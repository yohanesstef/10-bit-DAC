magic
tech sky130A
magscale 1 2
timestamp 1751042016
<< pwell >>
rect -151 -134 689 1279
<< mvpsubdiff >>
rect -115 1185 653 1243
rect -115 -40 -57 1185
rect 595 -40 653 1185
rect -115 -98 653 -40
<< locali >>
rect -103 1197 641 1231
rect -103 -52 -69 1197
rect 607 -52 641 1197
rect -103 -86 641 -52
<< metal1 >>
rect 279 961 289 1013
rect 341 961 351 1013
rect 23 856 75 866
rect 23 794 75 804
rect 23 616 75 626
rect 23 554 75 564
rect 23 376 75 386
rect 23 314 75 324
rect 205 146 233 866
rect 279 721 289 773
rect 341 721 351 773
rect 279 481 289 533
rect 341 481 351 533
rect 481 297 509 1017
rect 279 241 289 293
rect 341 241 351 293
rect 23 136 75 146
rect 23 74 75 84
<< via1 >>
rect 289 961 341 1013
rect 23 804 75 856
rect 23 564 75 616
rect 23 324 75 376
rect 289 721 341 773
rect 289 481 341 533
rect 289 241 341 293
rect 23 84 75 136
<< metal2 >>
rect 279 989 289 1013
rect 23 961 289 989
rect 341 961 351 1013
rect 23 862 51 961
rect 23 856 75 862
rect 23 794 75 804
rect 279 749 289 773
rect 23 721 289 749
rect 341 721 351 773
rect 23 622 51 721
rect 23 616 75 622
rect 23 554 75 564
rect 279 509 289 533
rect 23 481 289 509
rect 341 481 351 533
rect 23 382 51 481
rect 23 376 75 382
rect 23 314 75 324
rect 279 269 289 293
rect 23 241 289 269
rect 341 241 351 293
rect 23 142 51 241
rect 23 136 75 142
rect 23 74 75 84
use sky130_fd_pr__nfet_g5v0d10v5_MU5DNH  sky130_fd_pr__nfet_g5v0d10v5_MU5DNH_0
timestamp 1750848845
transform 1 0 131 0 1 495
box -108 -459 108 459
use sky130_fd_pr__nfet_g5v0d10v5_MU5DNH  sky130_fd_pr__nfet_g5v0d10v5_MU5DNH_1
timestamp 1750848845
transform 1 0 407 0 1 646
box -108 -459 108 459
<< end >>
