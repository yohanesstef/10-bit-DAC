magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1073 307 1073
<< psubdiff >>
rect -271 1003 -175 1037
rect 175 1003 271 1037
rect -271 941 -237 1003
rect 237 941 271 1003
rect -271 -1003 -237 -941
rect 237 -1003 271 -941
rect -271 -1037 -175 -1003
rect 175 -1037 271 -1003
<< psubdiffcont >>
rect -175 1003 175 1037
rect -271 -941 -237 941
rect 237 -941 271 941
rect -175 -1037 175 -1003
<< xpolycontact >>
rect -141 475 141 907
rect -141 -907 141 -475
<< xpolyres >>
rect -141 -475 141 475
<< locali >>
rect -271 1003 -175 1037
rect 175 1003 271 1037
rect -271 941 -237 1003
rect 237 941 271 1003
rect -271 -1003 -237 -941
rect 237 -1003 271 -941
rect -271 -1037 -175 -1003
rect 175 -1037 271 -1003
<< viali >>
rect -125 492 125 889
rect -125 -889 125 -492
<< metal1 >>
rect -131 889 131 901
rect -131 492 -125 889
rect 125 492 131 889
rect -131 480 131 492
rect -131 -492 131 -480
rect -131 -889 -125 -492
rect 125 -889 131 -492
rect -131 -901 131 -889
<< properties >>
string FIXED_BBOX -254 -1020 254 1020
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 4.91 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 7.231k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
