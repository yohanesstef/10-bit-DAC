magic
tech sky130A
magscale 1 2
timestamp 1748944356
<< xpolycontact >>
rect -141 60 141 492
rect -141 -492 141 -60
<< xpolyres >>
rect -141 -60 141 60
<< viali >>
rect -125 77 125 474
rect -125 -474 125 -77
<< metal1 >>
rect -131 474 131 486
rect -131 77 -125 474
rect 125 77 131 474
rect -131 65 131 77
rect -131 -77 131 -65
rect -131 -474 -125 -77
rect 125 -474 131 -77
rect -131 -486 131 -474
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 0.759 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 1.343k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
