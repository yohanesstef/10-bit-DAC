magic
tech sky130A
magscale 1 2
timestamp 1751042016
<< mvnmos >>
rect -129 -73 -29 11
rect 29 -73 129 11
<< mvndiff >>
rect -187 -1 -129 11
rect -187 -61 -175 -1
rect -141 -61 -129 -1
rect -187 -73 -129 -61
rect -29 -1 29 11
rect -29 -61 -17 -1
rect 17 -61 29 -1
rect -29 -73 29 -61
rect 129 -1 187 11
rect 129 -61 141 -1
rect 175 -61 187 -1
rect 129 -73 187 -61
<< mvndiffc >>
rect -175 -61 -141 -1
rect -17 -61 17 -1
rect 141 -61 175 -1
<< poly >>
rect -129 83 -29 99
rect -129 49 -113 83
rect -45 49 -29 83
rect -129 11 -29 49
rect 29 83 129 99
rect 29 49 45 83
rect 113 49 129 83
rect 29 11 129 49
rect -129 -99 -29 -73
rect 29 -99 129 -73
<< polycont >>
rect -113 49 -45 83
rect 45 49 113 83
<< locali >>
rect -129 49 -113 83
rect -45 49 -29 83
rect 29 49 45 83
rect 113 49 129 83
rect -175 -1 -141 15
rect -175 -77 -141 -61
rect -17 -1 17 15
rect -17 -77 17 -61
rect 141 -1 175 15
rect 141 -77 175 -61
<< viali >>
rect -105 49 -53 83
rect 53 49 105 83
rect -175 -61 -141 -1
rect -17 -61 17 -1
rect 141 -61 175 -1
<< metal1 >>
rect -117 83 -41 89
rect -117 49 -105 83
rect -53 49 -41 83
rect -117 43 -41 49
rect 41 83 117 89
rect 41 49 53 83
rect 105 49 117 83
rect 41 43 117 49
rect -181 -1 -135 11
rect -181 -61 -175 -1
rect -141 -61 -135 -1
rect -181 -73 -135 -61
rect -23 -1 23 11
rect -23 -61 -17 -1
rect 17 -61 23 -1
rect -23 -73 23 -61
rect 135 -1 181 11
rect 135 -61 141 -1
rect 175 -61 181 -1
rect 135 -73 181 -61
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.420 l 0.50 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
