magic
tech sky130A
magscale 1 2
timestamp 1749638674
<< error_p >>
rect -224 -182 -194 114
rect -158 -116 -128 48
rect 128 -116 158 48
rect -158 -120 158 -116
rect 194 -182 224 114
rect -224 -186 224 -182
<< nwell >>
rect -194 -182 194 148
<< mvpmos >>
rect -100 -120 100 48
<< mvpdiff >>
rect -158 -120 -100 48
rect 100 -120 158 48
<< poly >>
rect -100 129 100 145
rect -100 95 -84 129
rect 84 95 100 129
rect -100 48 100 95
rect -100 -146 100 -120
<< polycont >>
rect -84 95 84 129
<< locali >>
rect -100 95 -84 129
rect 84 95 100 129
<< viali >>
rect -42 95 42 129
<< metal1 >>
rect -54 129 54 135
rect -54 95 -42 129
rect 42 95 54 129
rect -54 89 54 95
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.84 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 50 viadrn 50 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
