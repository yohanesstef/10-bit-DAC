.subckt rseg_3_v3 v0 v1 v2 v3 v4 v5 v6 v7 v8 v9 v10 v11 v12 v13 v14 v15 v16 gnd
XR1 v0 v1 gnd sky130_fd_pr__res_xhigh_po_1p41 L=3.1677 mult=1 m=1
XR2 v1 v2 gnd sky130_fd_pr__res_xhigh_po_1p41 L=3.2702 mult=1 m=1
XR3 v2 v3 gnd sky130_fd_pr__res_xhigh_po_1p41 L=3.3214 mult=1 m=1
XR4 v3 v4 gnd sky130_fd_pr__res_xhigh_po_1p41 L=3.3727 mult=1 m=1
XR5 v4 v5 gnd sky130_fd_pr__res_xhigh_po_1p41 L=3.5265 mult=1 m=1
XR6 v5 v6 gnd sky130_fd_pr__res_xhigh_po_1p41 L=3.5777 mult=1 m=1
XR7 v6 v7 gnd sky130_fd_pr__res_xhigh_po_1p41 L=3.6802 mult=1 m=1
XR8 v7 v8 gnd sky130_fd_pr__res_xhigh_po_1p41 L=3.8340 mult=1 m=1
XR9 v8 v9 gnd sky130_fd_pr__res_xhigh_po_1p41 L=3.9364 mult=1 m=1
XR10 v9 v10 gnd sky130_fd_pr__res_xhigh_po_1p41 L=4.0902 mult=1 m=1
XR11 v10 v11 gnd sky130_fd_pr__res_xhigh_po_1p41 L=4.1928 mult=1 m=1
XR12 v11 v12 gnd sky130_fd_pr__res_xhigh_po_1p41 L=4.4490 mult=1 m=1
XR13 v12 v13 gnd sky130_fd_pr__res_xhigh_po_1p41 L=4.6028 mult=1 m=1
XR14 v13 v14 gnd sky130_fd_pr__res_xhigh_po_1p41 L=4.8590 mult=1 m=1
XR15 v14 v15 gnd sky130_fd_pr__res_xhigh_po_1p41 L=5.1153 mult=1 m=1
XR16 v15 v16 gnd sky130_fd_pr__res_xhigh_po_1p41 L=5.4229 mult=1 m=1
.ends