magic
tech sky130A
magscale 1 2
timestamp 1748963013
use sky130_fd_pr__res_xhigh_po_1p41_RP2U3Z  sky130_fd_pr__res_xhigh_po_1p41_RP2U3Z_0
timestamp 1748962452
transform 0 1 2700 1 0 -22895
box -141 -902 141 902
use sky130_fd_pr__res_xhigh_po_1p41_2NUKZQ  XR2 ~/10-bit-DAC/mag
timestamp 1748936551
transform 0 -1 2638 -1 0 -23219
box -141 -840 141 840
use sky130_fd_pr__res_xhigh_po_1p41_95YJ9M  XR3 ~/10-bit-DAC/mag
timestamp 1748936551
transform 0 -1 2587 -1 0 -23543
box -141 -789 141 789
use sky130_fd_pr__res_xhigh_po_1p41_GVNVJY  XR4 ~/10-bit-DAC/mag
timestamp 1748936551
transform 0 -1 2551 -1 0 -23867
box -141 -753 141 753
use sky130_fd_pr__res_xhigh_po_1p41_EEL3HT  XR5 ~/10-bit-DAC/mag
timestamp 1748936551
transform 0 -1 2526 -1 0 -24191
box -141 -728 141 728
use sky130_fd_pr__res_xhigh_po_1p41_S3DKJW  XR6 ~/10-bit-DAC/mag
timestamp 1748936551
transform 0 -1 2500 -1 0 -24515
box -141 -702 141 702
use sky130_fd_pr__res_xhigh_po_1p41_FZ95UC  XR7 ~/10-bit-DAC/mag
timestamp 1748936551
transform 0 -1 2480 -1 0 -24839
box -141 -682 141 682
use sky130_fd_pr__res_xhigh_po_1p41_GXMA4A  XR8 ~/10-bit-DAC/mag
timestamp 1748936551
transform 0 -1 2464 -1 0 -25163
box -141 -666 141 666
<< end >>
