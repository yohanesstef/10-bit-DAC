magic
tech sky130A
magscale 1 2
timestamp 1749478639
<< metal1 >>
rect 1979 -14566 2007 -14365
rect 2251 -14565 2279 -14364
rect 2525 -14567 2553 -14366
rect 2803 -14563 2831 -14362
rect 3082 -14576 3110 -14375
rect 3356 -14583 3384 -14382
rect 3629 -14587 3657 -14386
rect 3900 -14586 3928 -14385
rect 4180 -14581 4208 -14380
rect 4455 -14581 4483 -14380
use hnmos_16  hnmos_16_0
timestamp 1749478417
transform 1 0 1950 0 1 -14653
box -7 -5 4409 193
<< end >>
