magic
tech sky130A
magscale 1 2
timestamp 1748944356
<< xpolycontact >>
rect -141 101 141 533
rect -141 -533 141 -101
<< xpolyres >>
rect -141 -101 141 101
<< viali >>
rect -125 118 125 515
rect -125 -515 125 -118
<< metal1 >>
rect -131 515 131 527
rect -131 118 -125 515
rect 125 118 131 515
rect -131 106 131 118
rect -131 -118 131 -106
rect -131 -515 -125 -118
rect 125 -515 131 -118
rect -131 -527 131 -515
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.169 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 1.925k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
