magic
tech sky130A
magscale 1 2
timestamp 1750848845
<< pwell >>
rect -278 -629 278 629
<< mvnmos >>
rect -50 287 50 371
rect -50 47 50 131
rect -50 -193 50 -109
rect -50 -433 50 -349
<< mvndiff >>
rect -108 359 -50 371
rect -108 299 -96 359
rect -62 299 -50 359
rect -108 287 -50 299
rect 50 359 108 371
rect 50 299 62 359
rect 96 299 108 359
rect 50 287 108 299
rect -108 119 -50 131
rect -108 59 -96 119
rect -62 59 -50 119
rect -108 47 -50 59
rect 50 119 108 131
rect 50 59 62 119
rect 96 59 108 119
rect 50 47 108 59
rect -108 -121 -50 -109
rect -108 -181 -96 -121
rect -62 -181 -50 -121
rect -108 -193 -50 -181
rect 50 -121 108 -109
rect 50 -181 62 -121
rect 96 -181 108 -121
rect 50 -193 108 -181
rect -108 -361 -50 -349
rect -108 -421 -96 -361
rect -62 -421 -50 -361
rect -108 -433 -50 -421
rect 50 -361 108 -349
rect 50 -421 62 -361
rect 96 -421 108 -361
rect 50 -433 108 -421
<< mvndiffc >>
rect -96 299 -62 359
rect 62 299 96 359
rect -96 59 -62 119
rect 62 59 96 119
rect -96 -181 -62 -121
rect 62 -181 96 -121
rect -96 -421 -62 -361
rect 62 -421 96 -361
<< mvpsubdiff >>
rect -242 581 242 593
rect -242 547 -134 581
rect 134 547 242 581
rect -242 535 242 547
rect -242 485 -184 535
rect -242 -485 -230 485
rect -196 -485 -184 485
rect 184 485 242 535
rect -242 -535 -184 -485
rect 184 -485 196 485
rect 230 -485 242 485
rect 184 -535 242 -485
rect -242 -547 242 -535
rect -242 -581 -134 -547
rect 134 -581 242 -547
rect -242 -593 242 -581
<< mvpsubdiffcont >>
rect -134 547 134 581
rect -230 -485 -196 485
rect 196 -485 230 485
rect -134 -581 134 -547
<< poly >>
rect -50 443 50 459
rect -50 409 -34 443
rect 34 409 50 443
rect -50 371 50 409
rect -50 261 50 287
rect -50 203 50 219
rect -50 169 -34 203
rect 34 169 50 203
rect -50 131 50 169
rect -50 21 50 47
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -219 50 -193
rect -50 -277 50 -261
rect -50 -311 -34 -277
rect 34 -311 50 -277
rect -50 -349 50 -311
rect -50 -459 50 -433
<< polycont >>
rect -34 409 34 443
rect -34 169 34 203
rect -34 -71 34 -37
rect -34 -311 34 -277
<< locali >>
rect -230 547 -134 581
rect 134 547 230 581
rect -230 485 -196 547
rect 196 485 230 547
rect -50 409 -34 443
rect 34 409 50 443
rect -96 359 -62 375
rect -96 283 -62 299
rect 62 359 96 375
rect 62 283 96 299
rect -50 169 -34 203
rect 34 169 50 203
rect -96 119 -62 135
rect -96 43 -62 59
rect 62 119 96 135
rect 62 43 96 59
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -197 -62 -181
rect 62 -121 96 -105
rect 62 -197 96 -181
rect -50 -311 -34 -277
rect 34 -311 50 -277
rect -96 -361 -62 -345
rect -96 -437 -62 -421
rect 62 -361 96 -345
rect 62 -437 96 -421
rect -230 -547 -196 -485
rect 196 -547 230 -485
rect -230 -581 -134 -547
rect 134 -581 230 -547
<< viali >>
rect -26 409 26 443
rect -96 299 -62 359
rect 62 299 96 359
rect -26 169 26 203
rect -96 59 -62 119
rect 62 59 96 119
rect -26 -71 26 -37
rect -96 -181 -62 -121
rect 62 -181 96 -121
rect -26 -311 26 -277
rect -96 -421 -62 -361
rect 62 -421 96 -361
<< metal1 >>
rect -38 443 38 449
rect -38 409 -26 443
rect 26 409 38 443
rect -38 403 38 409
rect -102 359 -56 371
rect -102 299 -96 359
rect -62 299 -56 359
rect -102 287 -56 299
rect 56 359 102 371
rect 56 299 62 359
rect 96 299 102 359
rect 56 287 102 299
rect -38 203 38 209
rect -38 169 -26 203
rect 26 169 38 203
rect -38 163 38 169
rect -102 119 -56 131
rect -102 59 -96 119
rect -62 59 -56 119
rect -102 47 -56 59
rect 56 119 102 131
rect 56 59 62 119
rect 96 59 102 119
rect 56 47 102 59
rect -38 -37 38 -31
rect -38 -71 -26 -37
rect 26 -71 38 -37
rect -38 -77 38 -71
rect -102 -121 -56 -109
rect -102 -181 -96 -121
rect -62 -181 -56 -121
rect -102 -193 -56 -181
rect 56 -121 102 -109
rect 56 -181 62 -121
rect 96 -181 102 -121
rect 56 -193 102 -181
rect -38 -277 38 -271
rect -38 -311 -26 -277
rect 26 -311 38 -277
rect -38 -317 38 -311
rect -102 -361 -56 -349
rect -102 -421 -96 -361
rect -62 -421 -56 -361
rect -102 -433 -56 -421
rect 56 -361 102 -349
rect 56 -421 62 -361
rect 96 -421 102 -361
rect 56 -433 102 -421
<< properties >>
string FIXED_BBOX -213 -564 213 564
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.420 l 0.50 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
