magic
tech sky130A
timestamp 1748954881
<< end >>
