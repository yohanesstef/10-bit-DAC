magic
tech sky130A
magscale 1 2
timestamp 1750079478
<< pwell >>
rect -35 -39 7037 5101
<< mvpsubdiffcont >>
rect 74 5018 6928 5052
rect 14 3536 48 4992
rect 6954 3536 6988 4992
rect 14 3502 6988 3536
rect 14 2020 48 3502
rect 6954 2020 6988 3502
rect 14 1986 6988 2020
rect 14 1032 48 1986
rect 6954 1032 6988 1986
rect 14 998 6988 1032
rect 14 70 48 998
rect 6954 70 6988 998
rect 74 10 6928 44
<< viali >>
rect 14 5018 74 5052
rect 74 5018 6928 5052
rect 6928 5018 6988 5052
rect 14 4992 48 5018
rect 14 3536 48 4992
rect 6954 4992 6988 5018
rect 6954 3536 6988 4992
rect 14 3502 6988 3536
rect 14 2020 48 3502
rect 6954 2020 6988 3502
rect 14 1986 6988 2020
rect 14 1032 48 1986
rect 6954 1032 6988 1986
rect 14 998 6988 1032
rect 14 70 48 998
rect 14 44 48 70
rect 6954 70 6988 998
rect 6954 44 6988 70
rect 14 10 74 44
rect 74 10 6928 44
rect 6928 10 6988 44
<< metal2 >>
rect 3022 4909 3032 4965
rect 3088 4909 3098 4965
rect 3148 4733 3158 4789
rect 3214 4733 3224 4789
rect 3904 4645 3914 4701
rect 3970 4645 3980 4701
rect 2931 4525 3728 4527
rect 2931 4469 3662 4525
rect 3718 4469 3728 4525
rect 2931 4467 3728 4469
rect 3778 4117 3788 4173
rect 3844 4117 3854 4173
rect 3274 4029 3284 4085
rect 3340 4029 3350 4085
rect 3400 3733 3478 3735
rect 3400 3677 3410 3733
rect 3466 3677 3478 3733
rect 3400 3675 3478 3677
rect 3524 3645 3602 3647
rect 3524 3589 3536 3645
rect 3592 3589 3602 3645
rect 3524 3587 3602 3589
rect 3406 3449 3602 3451
rect 3406 3393 3536 3449
rect 3592 3393 3602 3449
rect 3406 3391 3602 3393
rect 3400 3361 3596 3363
rect 3400 3305 3410 3361
rect 3466 3305 3596 3361
rect 3400 3303 3596 3305
rect 3274 2953 3284 3009
rect 3340 2953 3350 3009
rect 3778 2865 3788 2921
rect 3844 2865 3854 2921
rect 3652 2569 4198 2571
rect 3652 2513 3662 2569
rect 3718 2513 4198 2569
rect 3652 2511 4198 2513
rect 3904 2337 3914 2393
rect 3970 2337 3980 2393
rect 3148 2249 3158 2305
rect 3214 2249 3224 2305
rect 3022 2073 3032 2129
rect 3088 2073 3098 2129
<< via2 >>
rect 3032 4909 3088 4965
rect 3158 4733 3214 4789
rect 3914 4645 3970 4701
rect 3662 4469 3718 4525
rect 3788 4117 3844 4173
rect 3284 4029 3340 4085
rect 3410 3677 3466 3733
rect 3536 3589 3592 3645
rect 3536 3393 3592 3449
rect 3410 3305 3466 3361
rect 3284 2953 3340 3009
rect 3788 2865 3844 2921
rect 3662 2513 3718 2569
rect 3914 2337 3970 2393
rect 3158 2249 3214 2305
rect 3032 2073 3088 2129
<< metal3 >>
rect 3027 4965 3093 4975
rect 3027 4909 3032 4965
rect 3088 4909 3093 4965
rect 3027 2129 3093 4909
rect 3027 2073 3032 2129
rect 3088 2073 3093 2129
rect 3027 1757 3093 2073
rect 3153 4789 3219 4794
rect 3153 4733 3158 4789
rect 3214 4733 3219 4789
rect 3153 2305 3219 4733
rect 3909 4701 3975 4711
rect 3909 4645 3914 4701
rect 3970 4645 3975 4701
rect 3657 4525 3723 4535
rect 3657 4469 3662 4525
rect 3718 4469 3723 4525
rect 3153 2249 3158 2305
rect 3214 2249 3219 2305
rect 3153 2043 3219 2249
rect 3279 4085 3345 4090
rect 3279 4029 3284 4085
rect 3340 4029 3345 4085
rect 3279 3009 3345 4029
rect 3279 2953 3284 3009
rect 3340 2953 3345 3009
rect 3279 2043 3345 2953
rect 3405 3733 3471 3738
rect 3405 3677 3410 3733
rect 3466 3677 3471 3733
rect 3405 3361 3471 3677
rect 3405 3305 3410 3361
rect 3466 3305 3471 3361
rect 3405 2043 3471 3305
rect 3531 3645 3597 3650
rect 3531 3589 3536 3645
rect 3592 3589 3597 3645
rect 3531 3449 3597 3589
rect 3531 3393 3536 3449
rect 3592 3393 3597 3449
rect 3531 2043 3597 3393
rect 3657 2569 3723 4469
rect 3657 2513 3662 2569
rect 3718 2513 3723 2569
rect 3657 2043 3723 2513
rect 3783 4173 3849 4178
rect 3783 4117 3788 4173
rect 3844 4117 3849 4173
rect 3783 2921 3849 4117
rect 3783 2865 3788 2921
rect 3844 2865 3849 2921
rect 3783 2043 3849 2865
rect 3909 2393 3975 4645
rect 3909 2337 3914 2393
rect 3970 2337 3975 2393
rect 3909 2043 3975 2337
use cm_ncell1  cm_ncell1_0
timestamp 1750060524
transform 1 0 29 0 1 972
box -38 -985 6982 1071
use cm_ncell2  cm_ncell2_0
timestamp 1750079478
transform 1 0 -15 0 1 3492
box 6 -1529 7026 1583
<< end >>
