magic
tech sky130A
magscale 1 2
timestamp 1749621435
<< error_p >>
rect -29 341 29 347
rect -29 307 -17 341
rect -29 301 29 307
<< nmos >>
rect -15 -331 15 269
<< ndiff >>
rect -73 257 -15 269
rect -73 -319 -61 257
rect -27 -319 -15 257
rect -73 -331 -15 -319
rect 15 257 73 269
rect 15 -319 27 257
rect 61 -319 73 257
rect 15 -331 73 -319
<< ndiffc >>
rect -61 -319 -27 257
rect 27 -319 61 257
<< poly >>
rect -33 341 33 357
rect -33 307 -17 341
rect 17 307 33 341
rect -33 291 33 307
rect -15 269 15 291
rect -15 -357 15 -331
<< polycont >>
rect -17 307 17 341
<< locali >>
rect -33 307 -17 341
rect 17 307 33 341
rect -61 257 -27 273
rect -61 -335 -27 -319
rect 27 257 61 273
rect 27 -335 61 -319
<< viali >>
rect -17 307 17 341
rect -61 -319 -27 257
rect 27 -319 61 257
<< metal1 >>
rect -29 341 29 347
rect -29 307 -17 341
rect 17 307 29 341
rect -29 301 29 307
rect -67 257 -21 269
rect -67 -319 -61 257
rect -27 -319 -21 257
rect -67 -331 -21 -319
rect 21 257 67 269
rect 21 -319 27 257
rect 61 -319 67 257
rect 21 -331 67 -319
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
