magic
tech sky130A
magscale 1 2
timestamp 1751042016
<< metal1 >>
rect 40745 21212 40805 21218
rect 40481 20870 40541 20876
rect 39087 19788 39147 19794
rect 38735 19578 38795 19584
rect 38735 14697 38795 19518
rect 38735 14631 38795 14637
rect 38823 19358 38883 19364
rect 38823 14609 38883 19298
rect 38823 14543 38883 14549
rect 38911 19192 38971 19198
rect 38911 14521 38971 19132
rect 38911 14455 38971 14461
rect 38999 18850 39059 18856
rect 38999 14433 39059 18790
rect 38999 14367 39059 14373
rect 39087 14345 39147 19728
rect 39087 14279 39147 14285
rect 39175 19446 39235 19452
rect 39175 14257 39235 19386
rect 40481 19358 40541 20810
rect 40481 19292 40541 19298
rect 40569 20528 40629 20534
rect 40569 19192 40629 20468
rect 40569 19126 40629 19132
rect 40657 20186 40717 20192
rect 39175 14191 39235 14197
rect 39263 19104 39323 19110
rect 39263 14169 39323 19044
rect 40657 18850 40717 20126
rect 40745 19578 40805 21152
rect 40745 19512 40805 19518
rect 40657 18784 40717 18790
rect 39263 14103 39323 14109
rect 39351 18762 39411 18768
rect 39351 14081 39411 18702
rect 39351 14015 39411 14021
rect 39439 18364 39499 18370
rect 39439 13993 39499 18304
rect 39791 18276 39851 18282
rect 39439 13927 39499 13933
rect 39527 18023 39587 18029
rect 39527 13905 39587 17963
rect 39527 13839 39587 13845
rect 39615 17680 39675 17686
rect 39615 13817 39675 17620
rect 39615 13751 39675 13757
rect 39703 17338 39763 17344
rect 39703 13729 39763 17278
rect 39703 13663 39763 13669
rect 39791 13641 39851 18216
rect 39791 13575 39851 13581
rect 39879 17934 39939 17940
rect 39879 13553 39939 17874
rect 40495 17592 40555 17598
rect 39879 13487 39939 13493
rect 39967 16532 40027 16538
rect 39967 13465 40027 16472
rect 40495 16532 40555 17532
rect 40495 16466 40555 16472
rect 40583 17250 40643 17256
rect 39967 13399 40027 13405
rect 40055 16444 40115 16450
rect 40055 13377 40115 16384
rect 40583 16444 40643 17190
rect 40583 16378 40643 16384
rect 40055 13311 40115 13317
rect 40143 16356 40203 16362
rect 40143 13289 40203 16296
rect 40143 13223 40203 13229
rect 40231 16268 40291 16274
rect 40231 13201 40291 16208
rect 40231 13135 40291 13141
rect 40319 15366 40379 15372
rect 40319 13113 40379 15306
rect 40319 13047 40379 13053
rect 40407 15278 40467 15284
rect 40407 13025 40467 15218
rect 40987 14376 41047 14382
rect 40407 12959 40467 12965
rect 40495 13386 40555 13392
rect 40495 12761 40555 13326
rect 40495 12695 40555 12701
rect 40583 13298 40643 13304
rect 40583 12673 40643 13238
rect 40987 12937 41047 14316
rect 40987 12871 41047 12877
rect 41075 14288 41135 14294
rect 41075 12849 41135 14228
rect 41075 12783 41135 12789
rect 40577 12613 40583 12673
rect 40643 12613 40649 12673
rect 40577 12525 40583 12585
rect 40643 12525 40649 12585
rect 40495 12497 40555 12503
rect 40407 12409 40467 12415
rect 40319 12321 40379 12327
rect 40231 12233 40291 12239
rect 40143 12145 40203 12151
rect 40055 12057 40115 12063
rect 39967 11969 40027 11975
rect 39879 11881 39939 11887
rect 39791 11793 39851 11799
rect 39791 8117 39851 11733
rect 39879 8205 39939 11821
rect 39967 8293 40027 11909
rect 40055 9283 40115 11997
rect 40143 10328 40203 12085
rect 40231 10416 40291 12173
rect 40319 11318 40379 12261
rect 40407 11406 40467 12349
rect 40495 12308 40555 12437
rect 40583 12396 40643 12525
rect 40583 12330 40643 12336
rect 40495 12242 40555 12248
rect 40407 11340 40467 11346
rect 40319 11252 40379 11258
rect 40231 10350 40291 10356
rect 40143 10262 40203 10268
rect 40055 9217 40115 9223
rect 39967 8227 40027 8233
rect 39879 8139 39939 8145
rect 41075 8205 41135 8211
rect 39791 8051 39851 8057
rect 40987 8117 41047 8123
rect 40987 6313 41047 8057
rect 41075 7303 41135 8145
rect 41075 7237 41135 7243
rect 40987 6247 41047 6253
<< via1 >>
rect 40745 21152 40805 21212
rect 40481 20810 40541 20870
rect 39087 19728 39147 19788
rect 38735 19518 38795 19578
rect 38735 14637 38795 14697
rect 38823 19298 38883 19358
rect 38823 14549 38883 14609
rect 38911 19132 38971 19192
rect 38911 14461 38971 14521
rect 38999 18790 39059 18850
rect 38999 14373 39059 14433
rect 39087 14285 39147 14345
rect 39175 19386 39235 19446
rect 40481 19298 40541 19358
rect 40569 20468 40629 20528
rect 40569 19132 40629 19192
rect 40657 20126 40717 20186
rect 39175 14197 39235 14257
rect 39263 19044 39323 19104
rect 40745 19518 40805 19578
rect 40657 18790 40717 18850
rect 39263 14109 39323 14169
rect 39351 18702 39411 18762
rect 39351 14021 39411 14081
rect 39439 18304 39499 18364
rect 39791 18216 39851 18276
rect 39439 13933 39499 13993
rect 39527 17963 39587 18023
rect 39527 13845 39587 13905
rect 39615 17620 39675 17680
rect 39615 13757 39675 13817
rect 39703 17278 39763 17338
rect 39703 13669 39763 13729
rect 39791 13581 39851 13641
rect 39879 17874 39939 17934
rect 40495 17532 40555 17592
rect 39879 13493 39939 13553
rect 39967 16472 40027 16532
rect 40495 16472 40555 16532
rect 40583 17190 40643 17250
rect 39967 13405 40027 13465
rect 40055 16384 40115 16444
rect 40583 16384 40643 16444
rect 40055 13317 40115 13377
rect 40143 16296 40203 16356
rect 40143 13229 40203 13289
rect 40231 16208 40291 16268
rect 40231 13141 40291 13201
rect 40319 15306 40379 15366
rect 40319 13053 40379 13113
rect 40407 15218 40467 15278
rect 40987 14316 41047 14376
rect 40407 12965 40467 13025
rect 40495 13326 40555 13386
rect 40495 12701 40555 12761
rect 40583 13238 40643 13298
rect 40987 12877 41047 12937
rect 41075 14228 41135 14288
rect 41075 12789 41135 12849
rect 40583 12613 40643 12673
rect 40583 12525 40643 12585
rect 40495 12437 40555 12497
rect 40407 12349 40467 12409
rect 40319 12261 40379 12321
rect 40231 12173 40291 12233
rect 40143 12085 40203 12145
rect 40055 11997 40115 12057
rect 39967 11909 40027 11969
rect 39879 11821 39939 11881
rect 39791 11733 39851 11793
rect 40583 12336 40643 12396
rect 40495 12248 40555 12308
rect 40407 11346 40467 11406
rect 40319 11258 40379 11318
rect 40231 10356 40291 10416
rect 40143 10268 40203 10328
rect 40055 9223 40115 9283
rect 39967 8233 40027 8293
rect 39879 8145 39939 8205
rect 41075 8145 41135 8205
rect 39791 8057 39851 8117
rect 40987 8057 41047 8117
rect 41075 7243 41135 7303
rect 40987 6253 41047 6313
<< metal2 >>
rect 40739 21152 40745 21212
rect 40805 21152 40833 21212
rect 40475 20810 40481 20870
rect 40541 20810 40833 20870
rect 40563 20468 40569 20528
rect 40629 20468 40833 20528
rect 40651 20126 40657 20186
rect 40717 20126 40835 20186
rect 39081 19728 39087 19788
rect 39147 19728 40833 19788
rect 38729 19518 38735 19578
rect 38795 19518 40745 19578
rect 40805 19518 40811 19578
rect 39169 19386 39175 19446
rect 39235 19386 40833 19446
rect 38817 19298 38823 19358
rect 38883 19298 40481 19358
rect 40541 19298 40547 19358
rect 38905 19132 38911 19192
rect 38971 19132 40569 19192
rect 40629 19132 40635 19192
rect 39257 19044 39263 19104
rect 39323 19044 40833 19104
rect 38993 18790 38999 18850
rect 39059 18790 40657 18850
rect 40717 18790 40723 18850
rect 39345 18702 39351 18762
rect 39411 18702 40833 18762
rect 39433 18304 39439 18364
rect 39499 18304 40027 18364
rect 39785 18216 39791 18276
rect 39851 18216 40133 18276
rect 39521 17963 39527 18023
rect 39587 18022 39593 18023
rect 39587 17963 39992 18022
rect 39873 17874 39879 17934
rect 39939 17874 39991 17934
rect 39609 17620 39615 17680
rect 39675 17620 39991 17680
rect 40399 17532 40495 17592
rect 40555 17532 40561 17592
rect 39697 17278 39703 17338
rect 39763 17278 40045 17338
rect 40399 17190 40583 17250
rect 40643 17190 40649 17250
rect 39961 16472 39967 16532
rect 40027 16472 40495 16532
rect 40555 16472 40561 16532
rect 40049 16384 40055 16444
rect 40115 16384 40583 16444
rect 40643 16384 40649 16444
rect 40137 16296 40143 16356
rect 40203 16296 41182 16356
rect 40225 16208 40231 16268
rect 40291 16208 41182 16268
rect 40313 15306 40319 15366
rect 40379 15306 41182 15366
rect 40401 15218 40407 15278
rect 40467 15218 41182 15278
rect 15856 14637 38735 14697
rect 38795 14637 38801 14697
rect 15856 14549 38823 14609
rect 38883 14549 38889 14609
rect 15856 14461 38911 14521
rect 38971 14461 38977 14521
rect 15856 14373 38999 14433
rect 39059 14373 39065 14433
rect 15856 14285 39087 14345
rect 39147 14285 39153 14345
rect 40981 14316 40987 14376
rect 41047 14316 41182 14376
rect 15856 14197 39175 14257
rect 39235 14197 39241 14257
rect 41069 14228 41075 14288
rect 41135 14228 41182 14288
rect 15856 14109 39263 14169
rect 39323 14109 39329 14169
rect 15856 14021 39351 14081
rect 39411 14021 39417 14081
rect 15856 13933 39439 13993
rect 39499 13933 39505 13993
rect 15856 13845 39527 13905
rect 39587 13845 39593 13905
rect 15856 13757 39615 13817
rect 39675 13757 39681 13817
rect 15856 13669 39703 13729
rect 39763 13669 39769 13729
rect 15856 13581 39791 13641
rect 39851 13581 39857 13641
rect 15856 13493 39879 13553
rect 39939 13493 39945 13553
rect 15856 13405 39967 13465
rect 40027 13405 40033 13465
rect 15856 13317 40055 13377
rect 40115 13317 40121 13377
rect 40489 13326 40495 13386
rect 40555 13326 41182 13386
rect 15856 13229 40143 13289
rect 40203 13229 40209 13289
rect 40577 13238 40583 13298
rect 40643 13238 41425 13298
rect 15856 13141 40231 13201
rect 40291 13141 40297 13201
rect 15856 13053 40319 13113
rect 40379 13053 40385 13113
rect 15856 12965 40407 13025
rect 40467 12965 40473 13025
rect 15856 12877 40987 12937
rect 41047 12877 41053 12937
rect 15856 12789 41075 12849
rect 41135 12789 41141 12849
rect 15856 12701 40495 12761
rect 40555 12701 40561 12761
rect 15856 12613 40583 12673
rect 40643 12613 40649 12673
rect 15856 12525 40583 12585
rect 40643 12525 40649 12585
rect 15856 12437 40495 12497
rect 40555 12437 40561 12497
rect 15856 12349 40407 12409
rect 40467 12349 40473 12409
rect 40577 12336 40583 12396
rect 40643 12336 41182 12396
rect 15856 12261 40319 12321
rect 40379 12261 40385 12321
rect 40489 12248 40495 12308
rect 40555 12248 41182 12308
rect 15856 12173 40231 12233
rect 40291 12173 40297 12233
rect 15856 12085 40143 12145
rect 40203 12085 40209 12145
rect 15856 11997 40055 12057
rect 40115 11997 40121 12057
rect 15856 11909 39967 11969
rect 40027 11909 40033 11969
rect 15856 11821 39879 11881
rect 39939 11821 39945 11881
rect 15856 11733 39791 11793
rect 39851 11733 39857 11793
rect 40401 11346 40407 11406
rect 40467 11346 41182 11406
rect 40313 11258 40319 11318
rect 40379 11258 41182 11318
rect 40225 10356 40231 10416
rect 40291 10356 41182 10416
rect 40137 10268 40143 10328
rect 40203 10268 41182 10328
rect 40049 9223 40055 9283
rect 40115 9223 41182 9283
rect 39961 8233 39967 8293
rect 40027 8233 41187 8293
rect 39873 8145 39879 8205
rect 39939 8145 41075 8205
rect 41135 8145 41141 8205
rect 39785 8057 39791 8117
rect 39851 8057 40987 8117
rect 41047 8057 41053 8117
rect 41069 7243 41075 7303
rect 41135 7243 41184 7303
rect 40981 6253 40987 6313
rect 41047 6253 41190 6313
use top_dcell_bias  top_dcell_bias_0
timestamp 1751030423
transform 1 0 36407 0 1 18556
box -1184 -17354 10416 4891
<< labels >>
flabel space 41553 10066 41553 10066 0 FreeSans 4800 0 0 0 b[0]
flabel space 41488 11133 41488 11133 0 FreeSans 4800 0 0 0 b[1]
flabel space 41837 12124 41837 12124 0 FreeSans 4800 0 0 0 b[2]
flabel space 41681 13093 41681 13093 0 FreeSans 4800 0 0 0 b[3]
flabel space 41640 14029 41640 14029 0 FreeSans 4800 0 0 0 b[4]
flabel space 41547 14965 41547 14965 0 FreeSans 4800 0 0 0 b[5]
flabel space 41560 16047 41560 16047 0 FreeSans 4800 0 0 0 b[6]
flabel space 42322 17678 42322 17678 0 FreeSans 4800 0 0 0 DEC2
flabel space 41520 18935 41520 18935 0 FreeSans 4800 0 0 0 DEC1
flabel space 41600 20366 41600 20366 0 FreeSans 4800 0 0 0 DEC0
flabel space 41535 6045 41535 6045 0 FreeSans 4800 0 0 0 S1
flabel space 41715 6995 41715 6995 0 FreeSans 4800 0 0 0 S2
flabel space 41686 7954 41686 7954 0 FreeSans 4800 0 0 0 S3
flabel space 41705 8950 41705 8950 0 FreeSans 4800 0 0 0 S4
<< end >>
