magic
tech sky130A
magscale 1 2
timestamp 1743275510
<< pwell >>
rect -201 -659 201 659
<< psubdiff >>
rect -165 589 -69 623
rect 69 589 165 623
rect -165 527 -131 589
rect 131 527 165 589
rect -165 -589 -131 -527
rect 131 -589 165 -527
rect -165 -623 -69 -589
rect 69 -623 165 -589
<< psubdiffcont >>
rect -69 589 69 623
rect -165 -527 -131 527
rect 131 -527 165 527
rect -69 -623 69 -589
<< xpolycontact >>
rect -35 61 35 493
rect -35 -493 35 -61
<< xpolyres >>
rect -35 -61 35 61
<< locali >>
rect -165 589 -69 623
rect 69 589 165 623
rect -165 527 -131 589
rect 131 527 165 589
rect -165 -589 -131 -527
rect 131 -589 165 -527
rect -165 -623 -69 -589
rect 69 -623 165 -589
<< viali >>
rect -19 78 19 475
rect -19 -475 19 -78
<< metal1 >>
rect -25 475 25 487
rect -25 78 -19 475
rect 19 78 25 475
rect -25 66 25 78
rect -25 -78 25 -66
rect -25 -475 -19 -78
rect 19 -475 25 -78
rect -25 -487 25 -475
<< properties >>
string FIXED_BBOX -148 -606 148 606
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.769 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 5.469k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
