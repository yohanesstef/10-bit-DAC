magic
tech sky130A
magscale 1 2
timestamp 1751060805
<< metal1 >>
rect 14088 25946 14148 25952
rect 1273 25246 1673 25252
rect 1273 24177 1673 24646
rect 3802 25246 4202 25252
rect 3802 24320 4202 24646
rect 8227 25246 8627 25252
rect 8227 24318 8627 24646
rect 13078 25246 13478 25252
rect 13078 24333 13478 24646
rect 13066 21778 13478 24333
rect 13078 16009 13478 21778
rect 14088 14507 14148 25346
rect 14199 25246 14259 25252
rect 14199 14700 14259 24646
rect 15962 16593 16022 16599
rect 15612 16505 15672 16511
rect 14199 14634 14259 14640
rect 14806 16241 14866 16247
rect 14806 14620 14866 16181
rect 15156 16153 15216 16159
rect 15156 14620 15216 16093
rect 15612 14620 15672 16445
rect 15962 14620 16022 16533
rect 19953 16593 20013 18516
rect 19953 16527 20013 16533
rect 20230 16505 20290 18428
rect 20230 16439 20290 16445
rect 21944 16241 22004 17876
rect 21944 16175 22004 16181
rect 22220 16153 22280 18015
rect 22220 16087 22280 16093
rect 16150 14700 16210 14706
rect 16150 14554 16210 14640
rect 13068 6319 13494 12285
rect 14206 12281 14266 13123
rect 14302 12809 14362 13123
rect 14460 12897 14520 13123
rect 16300 12985 16360 13101
rect 16458 13073 16518 13101
rect 16458 13007 16518 13013
rect 16300 12919 16360 12925
rect 14460 12831 14520 12837
rect 14302 12743 14362 12749
rect 14206 12215 14266 12221
rect 16554 12193 16614 13101
rect 34310 12281 34370 12287
rect 16554 12127 16614 12133
rect 19209 12193 19269 12199
rect 19209 10387 19269 12133
rect 34310 10382 34370 12221
rect 13094 1303 13494 6319
rect 13094 697 13494 703
<< via1 >>
rect 14088 25346 14148 25946
rect 1273 24646 1673 25246
rect 3802 24646 4202 25246
rect 8227 24646 8627 25246
rect 13078 24646 13478 25246
rect 14199 24646 14259 25246
rect 15962 16533 16022 16593
rect 15612 16445 15672 16505
rect 14199 14640 14259 14700
rect 14806 16181 14866 16241
rect 15156 16093 15216 16153
rect 19953 16533 20013 16593
rect 20230 16445 20290 16505
rect 21944 16181 22004 16241
rect 22220 16093 22280 16153
rect 16150 14640 16210 14700
rect 1273 14078 1393 14278
rect 16458 13013 16518 13073
rect 16300 12925 16360 12985
rect 14460 12837 14520 12897
rect 14302 12749 14362 12809
rect 14206 12221 14266 12281
rect 34310 12221 34370 12281
rect 16554 12133 16614 12193
rect 19209 12133 19269 12193
rect 13094 703 13494 1303
<< metal2 >>
rect 12718 27146 13118 27246
rect 12718 26946 12818 27146
rect 13018 26946 13118 27146
rect 12718 26846 13118 26946
rect 15956 16533 15962 16593
rect 16022 16533 19953 16593
rect 20013 16533 20019 16593
rect 15606 16445 15612 16505
rect 15672 16445 20230 16505
rect 20290 16445 20296 16505
rect 14800 16181 14806 16241
rect 14866 16181 21944 16241
rect 22004 16181 22010 16241
rect 15150 16093 15156 16153
rect 15216 16093 22220 16153
rect 22280 16093 22286 16153
rect 14193 14640 14199 14700
rect 14259 14640 16150 14700
rect 16210 14640 16216 14700
rect 241 14278 641 14378
rect 13806 14302 14056 14358
rect 14112 14302 14122 14358
rect 241 14078 1273 14278
rect 1393 14137 1399 14278
rect 1393 14078 4340 14137
rect 241 13978 641 14078
rect 1219 14077 4340 14078
rect 13806 13945 13866 14302
rect 16800 14222 17206 14252
rect 16800 14164 17148 14194
rect 12976 13885 13866 13945
rect 13926 14052 14056 14108
rect 14112 14052 14122 14108
rect 13926 13857 13986 14052
rect 16788 13973 17090 14003
rect 16800 13915 17032 13945
rect 12976 13797 13986 13857
rect 14046 13803 14056 13859
rect 14112 13803 14122 13859
rect 14046 13769 14122 13803
rect 12976 13709 14122 13769
rect 16800 13724 16974 13754
rect 12976 13621 14122 13681
rect 16800 13666 16916 13696
rect 14046 13610 14122 13621
rect 12976 13533 13986 13593
rect 14046 13554 14056 13610
rect 14112 13554 14122 13610
rect 13926 13361 13986 13533
rect 16798 13475 16858 13505
rect 13926 13305 14056 13361
rect 14112 13305 14122 13361
rect 16770 13161 16800 13417
rect 16828 13249 16858 13475
rect 16886 13337 16916 13666
rect 16944 13425 16974 13724
rect 17002 13513 17032 13915
rect 17060 13601 17090 13973
rect 17118 13689 17148 14164
rect 17176 13777 17206 14222
rect 17176 13747 17234 13777
rect 17118 13659 17234 13689
rect 17060 13571 17234 13601
rect 17002 13483 17234 13513
rect 16944 13395 17234 13425
rect 16886 13307 17234 13337
rect 16828 13219 17234 13249
rect 16770 13131 17234 13161
rect 16452 13013 16458 13073
rect 16518 13013 17234 13073
rect 16294 12925 16300 12985
rect 16360 12925 17234 12985
rect 14454 12837 14460 12897
rect 14520 12837 17234 12897
rect 14296 12749 14302 12809
rect 14362 12749 17377 12809
rect 14200 12221 14206 12281
rect 14266 12221 34310 12281
rect 34370 12221 34376 12281
rect 16548 12133 16554 12193
rect 16614 12133 19209 12193
rect 19269 12133 19275 12193
<< via2 >>
rect 12818 26946 13018 27146
rect 14056 14302 14112 14358
rect 14056 14052 14112 14108
rect 14056 13803 14112 13859
rect 14056 13554 14112 13610
rect 14056 13305 14112 13361
<< metal3 >>
rect 12813 27146 13023 27151
rect 12813 26946 12818 27146
rect 13018 26946 13023 27146
rect 12813 26941 13023 26946
rect 12852 24233 12984 26941
rect 14046 14358 14122 14363
rect 14046 14302 14056 14358
rect 14112 14302 14122 14358
rect 14046 14297 14122 14302
rect 14046 14108 14122 14113
rect 14046 14052 14056 14108
rect 14112 14052 14122 14108
rect 14046 14047 14122 14052
rect 14046 13859 14122 13864
rect 14046 13803 14056 13859
rect 14112 13803 14122 13859
rect 14046 13798 14122 13803
rect 14046 13610 14122 13615
rect 14046 13554 14056 13610
rect 14112 13554 14122 13610
rect 14046 13549 14122 13554
rect 14046 13361 14122 13366
rect 14046 13305 14056 13361
rect 14112 13305 14122 13361
rect 14046 13300 14122 13305
use top_buffer_opamp  top_buffer_opamp_0
timestamp 1751058216
transform -1 0 672 0 1 11001
box -12462 -8798 520 13398
use top_final_switch  top_final_switch_0
timestamp 1751053439
transform 1 0 -361 0 1 12
box 14407 13089 17161 14608
use top_rseg_n_dcell  top_rseg_n_dcell_0
timestamp 1751058216
transform 1 0 1378 0 1 1016
box -1226 -1019 49823 26230
<< end >>
