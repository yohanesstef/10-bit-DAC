magic
tech sky130A
magscale 1 2
timestamp 1750845353
<< error_p >>
rect -174 716 -144 748
rect 144 716 174 748
rect -174 532 174 716
rect -144 498 144 532
rect -174 396 -144 428
rect 144 396 174 428
rect -174 212 174 396
rect -144 178 144 212
rect -174 76 -144 108
rect 144 76 174 108
rect -174 -108 174 76
rect -144 -142 144 -108
rect -174 -244 -144 -212
rect 144 -244 174 -212
rect -174 -428 174 -244
rect -144 -462 144 -428
rect -174 -748 -144 -532
rect -108 -682 -78 -598
rect 78 -682 108 -598
rect 144 -748 174 -532
<< nwell >>
rect -144 498 144 782
rect -144 178 144 462
rect -144 -142 144 142
rect -144 -462 144 -178
rect -144 -782 144 -498
<< mvpmos >>
rect -50 598 50 682
rect -50 278 50 362
rect -50 -42 50 42
rect -50 -362 50 -278
rect -50 -682 50 -598
<< mvpdiff >>
rect -108 670 -50 682
rect -108 610 -96 670
rect -62 610 -50 670
rect -108 598 -50 610
rect 50 670 108 682
rect 50 610 62 670
rect 96 610 108 670
rect 50 598 108 610
rect -108 350 -50 362
rect -108 290 -96 350
rect -62 290 -50 350
rect -108 278 -50 290
rect 50 350 108 362
rect 50 290 62 350
rect 96 290 108 350
rect 50 278 108 290
rect -108 30 -50 42
rect -108 -30 -96 30
rect -62 -30 -50 30
rect -108 -42 -50 -30
rect 50 30 108 42
rect 50 -30 62 30
rect 96 -30 108 30
rect 50 -42 108 -30
rect -108 -290 -50 -278
rect -108 -350 -96 -290
rect -62 -350 -50 -290
rect -108 -362 -50 -350
rect 50 -290 108 -278
rect 50 -350 62 -290
rect 96 -350 108 -290
rect 50 -362 108 -350
rect -108 -610 -50 -598
rect -108 -670 -96 -610
rect -62 -670 -50 -610
rect -108 -682 -50 -670
rect 50 -610 108 -598
rect 50 -670 62 -610
rect 96 -670 108 -610
rect 50 -682 108 -670
<< mvpdiffc >>
rect -96 610 -62 670
rect 62 610 96 670
rect -96 290 -62 350
rect 62 290 96 350
rect -96 -30 -62 30
rect 62 -30 96 30
rect -96 -350 -62 -290
rect 62 -350 96 -290
rect -96 -670 -62 -610
rect 62 -670 96 -610
<< poly >>
rect -50 763 50 779
rect -50 729 -34 763
rect 34 729 50 763
rect -50 682 50 729
rect -50 551 50 598
rect -50 517 -34 551
rect 34 517 50 551
rect -50 501 50 517
rect -50 443 50 459
rect -50 409 -34 443
rect 34 409 50 443
rect -50 362 50 409
rect -50 231 50 278
rect -50 197 -34 231
rect 34 197 50 231
rect -50 181 50 197
rect -50 123 50 139
rect -50 89 -34 123
rect 34 89 50 123
rect -50 42 50 89
rect -50 -89 50 -42
rect -50 -123 -34 -89
rect 34 -123 50 -89
rect -50 -139 50 -123
rect -50 -197 50 -181
rect -50 -231 -34 -197
rect 34 -231 50 -197
rect -50 -278 50 -231
rect -50 -409 50 -362
rect -50 -443 -34 -409
rect 34 -443 50 -409
rect -50 -459 50 -443
rect -50 -517 50 -501
rect -50 -551 -34 -517
rect 34 -551 50 -517
rect -50 -598 50 -551
rect -50 -729 50 -682
rect -50 -763 -34 -729
rect 34 -763 50 -729
rect -50 -779 50 -763
<< polycont >>
rect -34 729 34 763
rect -34 517 34 551
rect -34 409 34 443
rect -34 197 34 231
rect -34 89 34 123
rect -34 -123 34 -89
rect -34 -231 34 -197
rect -34 -443 34 -409
rect -34 -551 34 -517
rect -34 -763 34 -729
<< locali >>
rect -50 729 -34 763
rect 34 729 50 763
rect -96 670 -62 686
rect -96 594 -62 610
rect 62 670 96 686
rect 62 594 96 610
rect -50 517 -34 551
rect 34 517 50 551
rect -50 409 -34 443
rect 34 409 50 443
rect -96 350 -62 366
rect -96 274 -62 290
rect 62 350 96 366
rect 62 274 96 290
rect -50 197 -34 231
rect 34 197 50 231
rect -50 89 -34 123
rect 34 89 50 123
rect -96 30 -62 46
rect -96 -46 -62 -30
rect 62 30 96 46
rect 62 -46 96 -30
rect -50 -123 -34 -89
rect 34 -123 50 -89
rect -50 -231 -34 -197
rect 34 -231 50 -197
rect -96 -290 -62 -274
rect -96 -366 -62 -350
rect 62 -290 96 -274
rect 62 -366 96 -350
rect -50 -443 -34 -409
rect 34 -443 50 -409
rect -50 -551 -34 -517
rect 34 -551 50 -517
rect -96 -610 -62 -594
rect -96 -686 -62 -670
rect 62 -610 96 -594
rect 62 -686 96 -670
rect -50 -763 -34 -729
rect 34 -763 50 -729
<< viali >>
rect -26 729 26 763
rect -96 610 -62 670
rect 62 610 96 670
rect -26 517 26 551
rect -26 409 26 443
rect -96 290 -62 350
rect 62 290 96 350
rect -26 197 26 231
rect -26 89 26 123
rect -96 -30 -62 30
rect 62 -30 96 30
rect -26 -123 26 -89
rect -26 -231 26 -197
rect -96 -350 -62 -290
rect 62 -350 96 -290
rect -26 -443 26 -409
rect -26 -551 26 -517
rect -96 -670 -62 -610
rect 62 -670 96 -610
rect -26 -763 26 -729
<< metal1 >>
rect -38 763 38 769
rect -38 729 -26 763
rect 26 729 38 763
rect -38 723 38 729
rect -102 670 -56 682
rect -102 610 -96 670
rect -62 610 -56 670
rect -102 598 -56 610
rect 56 670 102 682
rect 56 610 62 670
rect 96 610 102 670
rect 56 598 102 610
rect -38 551 38 557
rect -38 517 -26 551
rect 26 517 38 551
rect -38 511 38 517
rect -38 443 38 449
rect -38 409 -26 443
rect 26 409 38 443
rect -38 403 38 409
rect -102 350 -56 362
rect -102 290 -96 350
rect -62 290 -56 350
rect -102 278 -56 290
rect 56 350 102 362
rect 56 290 62 350
rect 96 290 102 350
rect 56 278 102 290
rect -38 231 38 237
rect -38 197 -26 231
rect 26 197 38 231
rect -38 191 38 197
rect -38 123 38 129
rect -38 89 -26 123
rect 26 89 38 123
rect -38 83 38 89
rect -102 30 -56 42
rect -102 -30 -96 30
rect -62 -30 -56 30
rect -102 -42 -56 -30
rect 56 30 102 42
rect 56 -30 62 30
rect 96 -30 102 30
rect 56 -42 102 -30
rect -38 -89 38 -83
rect -38 -123 -26 -89
rect 26 -123 38 -89
rect -38 -129 38 -123
rect -38 -197 38 -191
rect -38 -231 -26 -197
rect 26 -231 38 -197
rect -38 -237 38 -231
rect -102 -290 -56 -278
rect -102 -350 -96 -290
rect -62 -350 -56 -290
rect -102 -362 -56 -350
rect 56 -290 102 -278
rect 56 -350 62 -290
rect 96 -350 102 -290
rect 56 -362 102 -350
rect -38 -409 38 -403
rect -38 -443 -26 -409
rect 26 -443 38 -409
rect -38 -449 38 -443
rect -38 -517 38 -511
rect -38 -551 -26 -517
rect 26 -551 38 -517
rect -38 -557 38 -551
rect -102 -610 -56 -598
rect -102 -670 -96 -610
rect -62 -670 -56 -610
rect -102 -682 -56 -670
rect 56 -610 102 -598
rect 56 -670 62 -610
rect 96 -670 102 -610
rect 56 -682 102 -670
rect -38 -729 38 -723
rect -38 -763 -26 -729
rect 26 -763 38 -729
rect -38 -769 38 -763
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 0.50 m 5 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
