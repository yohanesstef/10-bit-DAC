magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -694 307 694
<< psubdiff >>
rect -271 624 -175 658
rect 175 624 271 658
rect -271 562 -237 624
rect 237 562 271 624
rect -271 -624 -237 -562
rect 237 -624 271 -562
rect -271 -658 -175 -624
rect 175 -658 271 -624
<< psubdiffcont >>
rect -175 624 175 658
rect -271 -562 -237 562
rect 237 -562 271 562
rect -175 -658 175 -624
<< xpolycontact >>
rect -141 96 141 528
rect -141 -528 141 -96
<< xpolyres >>
rect -141 -96 141 96
<< locali >>
rect -271 624 -175 658
rect 175 624 271 658
rect -271 562 -237 624
rect 237 562 271 624
rect -271 -624 -237 -562
rect 237 -624 271 -562
rect -271 -658 -175 -624
rect 175 -658 271 -624
<< viali >>
rect -125 113 125 510
rect -125 -510 125 -113
<< metal1 >>
rect -131 510 131 522
rect -131 113 -125 510
rect 125 113 131 510
rect -131 101 131 113
rect -131 -113 131 -101
rect -131 -510 -125 -113
rect 125 -510 131 -113
rect -131 -522 131 -510
<< properties >>
string FIXED_BBOX -254 -641 254 641
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.118 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 1.852k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
