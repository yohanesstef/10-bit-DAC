* PEX produced on Wed Jun 11 01:32:36 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from top_segment_2.ext - technology: sky130A

.subckt top_segment_2_posim V0 V48 DEC0[0] DEC0[1] DEC0[2] DEC1[0] DEC1[1] DEC1[2] DEC1[3]
+ DEC2[0] DEC2[1] DEC2[2] DEC2[3] VH VL GND
X0 rseg_2_v3_0.v47.t2 V48.t0 GND.t78 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X1 a_4370_4223.t1 DEC0[1].t0 rseg_2_v3_0.v31.t1 GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X2 a_6452_6264.t0 DEC1[3].t0 a_5474_4223.t0 GND.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X3 rseg_2_v3_0.v15.t0 rseg_2_v3_0.v14.t0 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=5.32
X4 a_2438_4223.t1 DEC0[0].t0 rseg_2_v3_0.v2.t1 GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X5 GND.t72 GND.t73 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X6 a_3818_4223.t1 DEC0[2].t0 rseg_2_v3_0.v43.t0 GND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X7 a_3266_4223.t3 DEC0[0].t1 rseg_2_v3_0.v8.t0 GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X8 a_4646_4223.t1 DEC0[2].t1 V48.t1 GND.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 a_6176_6264.t2 DEC1[3].t1 a_3542_4223.t0 GND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X10 rseg_2_v3_0.v17.t0 rseg_2_v3_0.v18.t0 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=5.06
X11 GND.t85 GND.t86 GND.t42 sky130_fd_pr__res_xhigh_po_1p41 l=5.22
X12 a_2990_4223.t1 DEC0[0].t2 rseg_2_v3_0.v6.t1 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X13 GND.t43 GND.t44 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X14 rseg_2_v3_0.v45.t1 rseg_2_v3_0.v46.t2 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=5.88
X15 a_6176_6264.t1 DEC1[0].t0 a_4094_4223.t0 GND.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X16 a_3266_4223.t4 DEC0[1].t1 rseg_2_v3_0.v24.t0 GND.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X17 rseg_2_v3_0.v33.t2 rseg_2_v3_0.v34.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X18 a_2162_4223.t2 DEC0[1].t2 rseg_2_v3_0.v16.t2 GND.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X19 a_3542_4223.t1 DEC0[2].t2 rseg_2_v3_0.v41.t1 GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X20 a_2990_4223.t2 DEC0[1].t3 rseg_2_v3_0.v22.t1 GND.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X21 a_3818_4223.t3 DEC0[1].t4 rseg_2_v3_0.v27.t1 GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X22 a_1886_4223.t2 DEC0[0].t3 rseg_2_v3_0.v1.t1 GND.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X23 a_3266_4223.t2 DEC0[2].t3 rseg_2_v3_0.v40.t1 GND.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X24 a_7004_6264.t3 DEC1[1].t0 a_2714_4223.t0 GND.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X25 GND.t65 GND.t66 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X26 a_5900_6264.t1 DEC1[0].t1 a_5198_4223.t1 GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X27 rseg_2_v3_0.v43.t2 rseg_2_v3_0.v44.t2 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=5.58
X28 rseg_2_v3_0.v17.t2 rseg_2_v3_0.v16.t3 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X29 rseg_2_v3_0.v13.t0 rseg_2_v3_0.v12.t0 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=5.58
X30 a_1886_4223.t3 DEC0[1].t5 rseg_2_v3_0.v17.t1 GND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X31 VH.t0 DEC2[3].t0 a_7004_6264.t4 GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X32 GND.t32 GND.t33 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=11.57
X33 a_2714_4223.t3 DEC0[1].t6 rseg_2_v3_0.v20.t1 GND.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X34 a_1334_4223.t0 DEC0[2].t4 rseg_2_v3_0.v37.t1 GND.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X35 a_3542_4223.t3 DEC0[1].t7 rseg_2_v3_0.v25.t0 GND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X36 rseg_2_v3_0.v25.t2 rseg_2_v3_0.v26.t2 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X37 a_2162_4223.t0 DEC0[2].t5 rseg_2_v3_0.v32.t2 GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X38 rseg_2_v3_0.v3.t0 rseg_2_v3_0.v2.t0 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=9.22
X39 a_2990_4223.t0 DEC0[2].t6 rseg_2_v3_0.v38.t2 GND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X40 a_6728_6264.t4 DEC1[1].t1 a_1610_4223.t0 GND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X41 a_1610_4223.t2 DEC0[0].t4 rseg_2_v3_0.v3.t2 GND.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X42 rseg_2_v3_0.v39.t2 rseg_2_v3_0.v40.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X43 rseg_2_v3_0.v15.t1 rseg_2_v3_0.v16.t0 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X44 rseg_2_v3_0.v9.t0 rseg_2_v3_0.v10.t0 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=6.14
X45 rseg_2_v3_0.v7.t0 rseg_2_v3_0.v6.t0 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=7.01
X46 VL.t0 DEC2[3].t1 a_6728_6264.t0 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X47 rseg_2_v3_0.v1.t0 V0.t0 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=11.57
X48 VH.t3 DEC2[1].t0 a_6452_6264.t3 GND.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X49 rseg_2_v3_0.v37.t0 rseg_2_v3_0.v38.t1 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=5.01
X50 a_2714_4223.t1 DEC0[2].t7 rseg_2_v3_0.v36.t0 GND.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X51 a_1334_4223.t1 DEC0[0].t5 rseg_2_v3_0.v5.t1 GND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X52 a_2162_4223.t1 DEC0[0].t6 V0.t1 GND.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X53 rseg_2_v3_0.v25.t1 rseg_2_v3_0.v24.t2 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X54 a_4922_4223.t2 DEC0[0].t7 rseg_2_v3_0.v14.t2 GND.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X55 a_5474_4223.t2 DEC0[1].t8 rseg_2_v3_0.v26.t0 GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X56 GND.t87 GND.t88 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X57 VL.t3 DEC2[1].t1 a_6176_6264.t4 GND.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X58 GND.t61 GND.t62 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X59 a_1058_4223.t3 DEC0[1].t9 rseg_2_v3_0.v23.t1 GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X60 a_2438_4223.t0 DEC0[2].t8 rseg_2_v3_0.v34.t1 GND.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X61 a_1058_4223.t2 DEC0[0].t8 rseg_2_v3_0.v7.t1 GND.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X62 rseg_2_v3_0.v13.t1 rseg_2_v3_0.v14.t1 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=5.47
X63 a_5900_6264.t2 DEC1[1].t2 a_2162_4223.t3 GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X64 rseg_2_v3_0.v3.t1 rseg_2_v3_0.v4.t1 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=8.5
X65 rseg_2_v3_0.v21.t1 rseg_2_v3_0.v22.t2 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=4.81
X66 a_3818_4223.t2 DEC0[0].t9 rseg_2_v3_0.v11.t0 GND.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X67 a_4646_4223.t2 DEC0[0].t10 rseg_2_v3_0.v16.t1 GND.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X68 rseg_2_v3_0.v5.t2 rseg_2_v3_0.v6.t2 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=7.42
X69 rseg_2_v3_0.v35.t0 rseg_2_v3_0.v34.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=4.81
X70 rseg_2_v3_0.v1.t2 rseg_2_v3_0.v2.t2 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=10.24
X71 a_5474_4223.t1 DEC0[0].t11 rseg_2_v3_0.v10.t1 GND.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X72 a_1610_4223.t3 DEC0[1].t10 rseg_2_v3_0.v19.t1 GND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X73 rseg_2_v3_0.v23.t0 rseg_2_v3_0.v22.t0 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X74 a_2438_4223.t2 DEC0[1].t11 rseg_2_v3_0.v18.t1 GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X75 rseg_2_v3_0.v31.t0 rseg_2_v3_0.v32.t1 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X76 a_1058_4223.t0 DEC0[2].t9 rseg_2_v3_0.v39.t1 GND.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X77 VL.t1 DEC2[2].t0 a_6452_6264.t1 GND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X78 GND.t59 GND.t60 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X79 a_1886_4223.t1 DEC0[2].t10 rseg_2_v3_0.v33.t1 GND.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X80 a_6452_6264.t4 DEC1[1].t3 a_2438_4223.t3 GND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X81 rseg_2_v3_0.v45.t2 rseg_2_v3_0.v44.t1 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=5.73
X82 rseg_2_v3_0.v21.t2 rseg_2_v3_0.v20.t2 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X83 rseg_2_v3_0.v29.t1 rseg_2_v3_0.v30.t0 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X84 a_7004_6264.t0 DEC1[2].t0 a_3266_4223.t0 GND.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X85 a_4922_4223.t1 DEC0[2].t11 rseg_2_v3_0.v46.t1 GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X86 a_5198_4223.t4 DEC0[1].t12 rseg_2_v3_0.v28.t2 GND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X87 rseg_2_v3_0.v23.t2 rseg_2_v3_0.v24.t1 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X88 a_5198_4223.t3 DEC0[0].t12 rseg_2_v3_0.v12.t1 GND.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X89 a_4094_4223.t2 DEC0[0].t13 rseg_2_v3_0.v13.t2 GND.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X90 a_1334_4223.t3 DEC0[1].t13 rseg_2_v3_0.v21.t0 GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X91 a_1610_4223.t1 DEC0[2].t12 rseg_2_v3_0.v35.t1 GND.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X92 rseg_2_v3_0.v35.t2 rseg_2_v3_0.v36.t1 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X93 rseg_2_v3_0.v31.t2 rseg_2_v3_0.v30.t2 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X94 a_6176_6264.t3 DEC1[1].t4 a_1886_4223.t0 GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X95 a_5900_6264.t4 DEC1[2].t1 a_2714_4223.t4 GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X96 rseg_2_v3_0.v47.t1 rseg_2_v3_0.v46.t0 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=6.09
X97 a_6728_6264.t5 DEC1[2].t2 a_1058_4223.t1 GND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X98 VH.t2 DEC2[2].t1 a_6728_6264.t1 GND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X99 rseg_2_v3_0.v19.t0 rseg_2_v3_0.v20.t0 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X100 rseg_2_v3_0.v29.t0 rseg_2_v3_0.v28.t1 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X101 a_4094_4223.t3 DEC0[1].t14 rseg_2_v3_0.v29.t2 GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X102 a_5474_4223.t3 DEC0[2].t13 rseg_2_v3_0.v42.t0 GND.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X103 a_4922_4223.t3 DEC0[1].t15 rseg_2_v3_0.v30.t1 GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X104 a_6452_6264.t5 DEC1[2].t3 a_2990_4223.t3 GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X105 a_7004_6264.t1 DEC1[3].t2 a_5198_4223.t0 GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X106 a_4370_4223.t0 DEC0[2].t14 rseg_2_v3_0.v47.t0 GND.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X107 a_5198_4223.t2 DEC0[2].t15 rseg_2_v3_0.v44.t0 GND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X108 rseg_2_v3_0.v7.t2 rseg_2_v3_0.v8.t2 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=6.65
X109 rseg_2_v3_0.v43.t1 rseg_2_v3_0.v42.t1 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=5.47
X110 rseg_2_v3_0.v9.t2 rseg_2_v3_0.v8.t1 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X111 rseg_2_v3_0.v27.t2 rseg_2_v3_0.v26.t1 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X112 a_7004_6264.t2 DEC1[0].t2 a_4646_4223.t0 GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X113 GND.t75 GND.t76 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X114 a_6728_6264.t3 DEC1[0].t3 a_4370_4223.t3 GND.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X115 rseg_2_v3_0.v5.t0 rseg_2_v3_0.v4.t0 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=7.88
X116 GND.t103 GND.t104 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X117 rseg_2_v3_0.v41.t0 rseg_2_v3_0.v40.t0 GND.t42 sky130_fd_pr__res_xhigh_po_1p41 l=5.22
X118 rseg_2_v3_0.v39.t0 rseg_2_v3_0.v38.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=5.01
X119 GND.t101 GND.t102 GND.t78 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X120 a_6176_6264.t5 DEC1[2].t4 a_1334_4223.t2 GND.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X121 VH.t1 DEC2[0].t0 a_6176_6264.t0 GND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X122 rseg_2_v3_0.v37.t2 rseg_2_v3_0.v36.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=4.91
X123 a_4646_4223.t3 DEC0[1].t16 rseg_2_v3_0.v32.t3 GND.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X124 a_5900_6264.t0 DEC1[3].t3 a_3266_4223.t1 GND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X125 a_6728_6264.t2 DEC1[3].t4 a_3818_4223.t0 GND.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X126 a_4094_4223.t1 DEC0[2].t16 rseg_2_v3_0.v45.t0 GND.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X127 a_2714_4223.t2 DEC0[0].t14 rseg_2_v3_0.v4.t2 GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X128 rseg_2_v3_0.v11.t2 rseg_2_v3_0.v12.t2 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=5.73
X129 a_3542_4223.t2 DEC0[0].t15 rseg_2_v3_0.v9.t1 GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X130 a_4370_4223.t2 DEC0[0].t16 rseg_2_v3_0.v15.t2 GND.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X131 rseg_2_v3_0.v27.t0 rseg_2_v3_0.v28.t0 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X132 rseg_2_v3_0.v19.t2 rseg_2_v3_0.v18.t2 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=4.96
X133 rseg_2_v3_0.v41.t2 rseg_2_v3_0.v42.t2 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=5.32
X134 rseg_2_v3_0.v11.t1 rseg_2_v3_0.v10.t2 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=5.94
X135 a_6452_6264.t2 DEC1[0].t4 a_4922_4223.t0 GND.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X136 VL.t2 DEC2[0].t1 a_5900_6264.t3 GND.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X137 rseg_2_v3_0.v33.t0 rseg_2_v3_0.v32.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X138 GND.t2 GND.t3 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=6.65
R0 rseg_2_v3_0.v47.t0 rseg_2_v3_0.v47.n0 237.56
R1 rseg_2_v3_0.v47.n0 rseg_2_v3_0.v47.t1 10.6178
R2 rseg_2_v3_0.v47.n0 rseg_2_v3_0.v47.t2 10.5739
R3 V48.n0 V48.t1 238.077
R4 V48.n0 V48.t0 10.612
R5 V48 V48.n0 1.29821
R6 GND.n81 GND.n33 32327.7
R7 GND.n33 GND.n32 32324.4
R8 GND.n83 GND.n32 32321.1
R9 GND.n83 GND.n81 32317.8
R10 GND.n78 GND.n53 10050.6
R11 GND.n78 GND.n54 10050.6
R12 GND.n60 GND.n53 9474.26
R13 GND.n69 GND.n54 9474.26
R14 GND.n102 GND.n3 8548.9
R15 GND.n101 GND.n3 8548.9
R16 GND.n90 GND.n19 8548.9
R17 GND.n89 GND.n19 8548.9
R18 GND.n102 GND.n4 7972.6
R19 GND.n94 GND.n4 7972.6
R20 GND.n94 GND.n14 7972.6
R21 GND.n90 GND.n14 7972.6
R22 GND.n101 GND.n5 7972.6
R23 GND.n95 GND.n5 7972.6
R24 GND.n95 GND.n13 7972.6
R25 GND.n89 GND.n13 7972.6
R26 GND.n73 GND.n59 4597.17
R27 GND.n65 GND.n59 4597.17
R28 GND.n73 GND.n60 4020.88
R29 GND.n69 GND.n65 4020.88
R30 GND.n77 GND.n76 1153.51
R31 GND.n76 GND.n75 1083.11
R32 GND.n61 GND.n16 1083.11
R33 GND.n91 GND.n18 981.836
R34 GND.n83 GND.n82 926.929
R35 GND.n93 GND.n15 911.436
R36 GND.n93 GND.n92 911.436
R37 GND.n92 GND.n91 911.436
R38 GND.n62 GND.n61 739.765
R39 GND.n104 GND.n1 675.013
R40 GND.n63 GND.n2 601.977
R41 GND.n92 GND.n16 601.977
R42 GND.n62 GND.n15 601.977
R43 GND.n70 GND.n60 576.293
R44 GND.n70 GND.n69 576.293
R45 GND.n52 GND.n14 576.293
R46 GND.n52 GND.n13 576.293
R47 GND.n67 GND.n4 576.293
R48 GND.n67 GND.n5 576.293
R49 GND.n103 GND.n2 568.095
R50 GND.n84 GND.n23 566.203
R51 GND.n6 GND.n1 542.871
R52 GND.n74 GND.n56 530.072
R53 GND.n96 GND.n12 514.26
R54 GND.n100 GND.n99 496.188
R55 GND.n88 GND.n87 494.683
R56 GND.n87 GND.n18 487.154
R57 GND.n39 GND.n38 483.003
R58 GND.n98 GND.n97 475.86
R59 GND.n21 GND.n20 472.471
R60 GND.n85 GND.n84 461.243
R61 GND.n38 GND.n37 461.243
R62 GND.n75 GND.n74 459.671
R63 GND.n64 GND.n63 459.671
R64 GND.n100 GND.n6 438.966
R65 GND.n88 GND.n21 438.966
R66 GND.n97 GND.n96 435.577
R67 GND.n64 GND.n0 415.248
R68 GND.n99 GND.n98 415.248
R69 GND.n20 GND.n12 397.176
R70 GND.n86 GND.n85 390.416
R71 GND.n63 GND.n62 343.341
R72 GND.n15 GND.n2 343.341
R73 GND.n46 GND.n23 312.353
R74 GND.n104 GND.n103 306.825
R75 GND GND.n0 303.06
R76 GND.n48 GND.n47 299.553
R77 GND GND.n104 298.918
R78 GND.n47 GND.n46 253.26
R79 GND.n40 GND.n39 251.339
R80 GND.n42 GND.n41 249.207
R81 GND.n44 GND.n43 229.579
R82 GND.n50 GND.n49 226.463
R83 GND.n57 GND.n33 212.213
R84 GND.n41 GND.n40 188.194
R85 GND.n99 GND.n7 184.471
R86 GND.n97 GND.n11 184.471
R87 GND.n30 GND.n12 184.471
R88 GND.n27 GND.n21 184.471
R89 GND.n87 GND.n86 184.471
R90 GND.n36 GND.n6 184.471
R91 GND.n45 GND.n44 179.019
R92 GND.n37 GND.n36 179.004
R93 GND.n26 GND.n22 173.474
R94 GND.t71 GND.t89 173.19
R95 GND.t92 GND.t71 173.19
R96 GND.t82 GND.t92 173.19
R97 GND.t53 GND.t11 173.19
R98 GND.t12 GND.t0 173.19
R99 GND.t0 GND.t41 173.19
R100 GND.t41 GND.t7 173.19
R101 GND.t47 GND.t48 173.19
R102 GND.t48 GND.t91 173.19
R103 GND.t91 GND.t98 173.19
R104 GND.t81 GND.t51 173.19
R105 GND.t51 GND.t16 173.19
R106 GND.t16 GND.t39 173.19
R107 GND.t55 GND.t39 173.19
R108 GND.t55 GND.t36 173.19
R109 GND.t8 GND.t36 173.19
R110 GND.t9 GND.t8 173.19
R111 GND.t99 GND.t9 173.19
R112 GND.t56 GND.t99 173.19
R113 GND.t31 GND.t56 173.19
R114 GND.t13 GND.t23 173.19
R115 GND.n35 GND.n34 170.487
R116 GND.n25 GND.n24 170.274
R117 GND.t1 GND.t31 165.66
R118 GND.t46 GND.t63 155.619
R119 GND.t54 GND.t83 155.619
R120 GND.t77 GND.t80 155.619
R121 GND.n10 GND.n9 152.139
R122 GND.n31 GND.n30 151.696
R123 GND.n29 GND.n28 151.5
R124 GND.n67 GND.n8 146.25
R125 GND.n68 GND.n67 146.25
R126 GND.n52 GND.n17 146.25
R127 GND.n79 GND.n52 146.25
R128 GND.n19 GND.n18 146.25
R129 GND.n82 GND.n19 146.25
R130 GND.n59 GND.n56 146.25
R131 GND.n59 GND.n58 146.25
R132 GND.n70 GND.n55 146.25
R133 GND.n71 GND.n70 146.25
R134 GND.n78 GND.n77 146.25
R135 GND.n79 GND.n78 146.25
R136 GND.n3 GND.n1 146.25
R137 GND.n57 GND.n3 146.25
R138 GND.n80 GND.t84 143.697
R139 GND.n43 GND.n42 143.393
R140 GND.n28 GND.n27 138.897
R141 GND.t35 GND.t70 138.049
R142 GND.t21 GND.t93 138.049
R143 GND.t22 GND.t17 138.049
R144 GND.t30 GND.t49 138.049
R145 GND.n49 GND.n48 135.073
R146 GND.t89 GND.n57 133.657
R147 GND.t7 GND.n79 133.657
R148 GND.n79 GND.t47 133.657
R149 GND.n82 GND.t13 133.657
R150 GND.n11 GND.n10 133.137
R151 GND.n86 GND.n22 131.857
R152 GND.t25 GND.t57 131.774
R153 GND.t94 GND.t96 131.774
R154 GND.n34 GND.n7 125.457
R155 GND.t10 GND.t78 124.873
R156 GND.n36 GND.n35 120.55
R157 GND.t19 GND.t27 120.48
R158 GND.t50 GND.t58 120.48
R159 GND.n56 GND.n0 114.825
R160 GND.t6 GND.t12 110.439
R161 GND.n27 GND.n26 110.311
R162 GND.n58 GND.t10 107.302
R163 GND.n9 GND.n7 106.257
R164 GND.t24 GND.t4 106.047
R165 GND.t95 GND.t40 105.419
R166 GND.t28 GND.t37 105.419
R167 GND.t100 GND.t74 102.909
R168 GND.n24 GND.n11 96.4436
R169 GND.n72 GND.t79 95.3798
R170 GND.n66 GND.t26 95.3798
R171 GND.n71 GND.t18 92.2424
R172 GND.t68 GND.n68 92.2424
R173 GND.t98 GND.t15 92.2424
R174 GND.n30 GND.n29 88.9769
R175 GND.t20 GND.t34 87.8499
R176 GND.t14 GND.t52 87.8499
R177 GND.t97 GND.t5 85.9674
R178 GND.t37 GND.t34 85.3399
R179 GND.t20 GND.t52 85.3399
R180 GND.t67 GND.n71 80.9474
R181 GND.n68 GND.t38 80.9474
R182 GND.t15 GND.t81 80.9474
R183 GND.n75 GND.n55 70.4005
R184 GND.n63 GND.n55 70.4005
R185 GND.n77 GND.n16 70.4005
R186 GND.n92 GND.n17 70.4005
R187 GND.n20 GND.n17 70.4005
R188 GND.n15 GND.n8 70.4005
R189 GND.n98 GND.n8 70.4005
R190 GND.t79 GND.t100 70.28
R191 GND.t74 GND.t19 70.28
R192 GND.t29 GND.t95 67.77
R193 GND.t40 GND.t28 67.77
R194 GND.n58 GND.t29 65.8875
R195 GND.t11 GND.t6 62.7501
R196 GND.t90 GND.n66 60.2401
R197 GND.t27 GND.t24 52.7101
R198 GND.t64 GND.t67 52.7101
R199 GND.t38 GND.t50 52.7101
R200 GND.t58 GND.t35 52.7101
R201 GND.t5 GND.t105 52.0826
R202 GND.t42 GND.t82 41.4152
R203 GND.t18 GND.t25 41.4152
R204 GND.t57 GND.t94 41.4152
R205 GND.t96 GND.t68 41.4152
R206 GND.n35 GND.t102 39.3159
R207 GND.n34 GND.t103 39.3159
R208 GND.n9 GND.t104 39.3159
R209 GND.n10 GND.t61 39.3159
R210 GND.n24 GND.t62 39.3159
R211 GND.n25 GND.t43 39.3159
R212 GND.n29 GND.t44 39.3159
R213 GND.n28 GND.t65 39.3159
R214 GND.n26 GND.t66 39.3159
R215 GND.n22 GND.t32 39.3159
R216 GND.n85 GND.t33 39.3159
R217 GND.n23 GND.t3 39.3159
R218 GND.n46 GND.t2 39.3159
R219 GND.n47 GND.t73 39.3159
R220 GND.n48 GND.t72 39.3159
R221 GND.n49 GND.t76 39.3159
R222 GND.n45 GND.t75 39.3159
R223 GND.n44 GND.t60 39.3159
R224 GND.n43 GND.t59 39.3159
R225 GND.n42 GND.t88 39.3159
R226 GND.n41 GND.t87 39.3159
R227 GND.n40 GND.t86 39.3159
R228 GND.n39 GND.t85 39.3159
R229 GND.n37 GND.t101 39.3159
R230 GND.t70 GND.t21 35.1403
R231 GND.t93 GND.t97 35.1403
R232 GND.t105 GND.t22 35.1403
R233 GND.t17 GND.t30 35.1403
R234 GND.t49 GND.t90 35.1403
R235 GND.t26 GND.t46 17.5704
R236 GND.t54 GND.t63 17.5704
R237 GND.t80 GND.t83 17.5704
R238 GND.t69 GND.t77 17.5704
R239 GND.t84 GND.t53 17.5704
R240 GND.n65 GND.n64 17.2064
R241 GND.n72 GND.n65 17.2064
R242 GND.n74 GND.n73 17.2064
R243 GND.n73 GND.n72 17.2064
R244 GND.t4 GND.t64 14.4329
R245 GND.n84 GND.n83 13.296
R246 GND.n38 GND.n33 13.296
R247 GND.n51 GND.t69 11.2954
R248 GND.n89 GND.n88 8.47876
R249 GND.t55 GND.n89 8.47876
R250 GND.n96 GND.n95 8.47876
R251 GND.n95 GND.t54 8.47876
R252 GND.n101 GND.n100 8.47876
R253 GND.t20 GND.n101 8.47876
R254 GND.n91 GND.n90 8.47876
R255 GND.n90 GND.t55 8.47876
R256 GND.n94 GND.n93 8.47876
R257 GND.t54 GND.n94 8.47876
R258 GND.n103 GND.n102 8.47876
R259 GND.n102 GND.t20 8.47876
R260 GND.n72 GND.t14 7.53045
R261 GND.t23 GND.t1 7.53045
R262 GND.n61 GND.n54 7.13465
R263 GND.n66 GND.n54 7.13465
R264 GND.n76 GND.n53 7.13465
R265 GND.n66 GND.n53 7.13465
R266 GND.n31 GND.n25 6.4005
R267 GND.t45 GND.t42 6.27546
R268 GND.n50 GND.n45 3.11845
R269 GND.n32 GND.n31 2.51123
R270 GND.n51 GND.n32 2.51123
R271 GND.n81 GND.n50 2.51123
R272 GND.n81 GND.n80 2.51123
R273 GND.t78 GND.t45 0.627996
R274 GND.n80 GND.n51 0.627996
R275 DEC0[1].n0 DEC0[1].t8 213.218
R276 DEC0[1].n15 DEC0[1].t9 212.554
R277 DEC0[1].n14 DEC0[1].t13 212.554
R278 DEC0[1].n13 DEC0[1].t10 212.554
R279 DEC0[1].n12 DEC0[1].t5 212.554
R280 DEC0[1].n11 DEC0[1].t2 212.554
R281 DEC0[1].n10 DEC0[1].t11 212.554
R282 DEC0[1].n9 DEC0[1].t6 212.554
R283 DEC0[1].n8 DEC0[1].t3 212.554
R284 DEC0[1].n7 DEC0[1].t1 212.554
R285 DEC0[1].n6 DEC0[1].t7 212.554
R286 DEC0[1].n5 DEC0[1].t4 212.554
R287 DEC0[1].n4 DEC0[1].t14 212.554
R288 DEC0[1].n3 DEC0[1].t0 212.554
R289 DEC0[1].n2 DEC0[1].t16 212.554
R290 DEC0[1].n1 DEC0[1].t15 212.554
R291 DEC0[1].n0 DEC0[1].t12 212.554
R292 DEC0[1].n1 DEC0[1].n0 0.663962
R293 DEC0[1].n2 DEC0[1].n1 0.663962
R294 DEC0[1].n3 DEC0[1].n2 0.663962
R295 DEC0[1].n4 DEC0[1].n3 0.663962
R296 DEC0[1].n5 DEC0[1].n4 0.663962
R297 DEC0[1].n6 DEC0[1].n5 0.663962
R298 DEC0[1].n7 DEC0[1].n6 0.663962
R299 DEC0[1].n8 DEC0[1].n7 0.663962
R300 DEC0[1].n9 DEC0[1].n8 0.663962
R301 DEC0[1].n10 DEC0[1].n9 0.663962
R302 DEC0[1].n11 DEC0[1].n10 0.663962
R303 DEC0[1].n12 DEC0[1].n11 0.663962
R304 DEC0[1].n13 DEC0[1].n12 0.663962
R305 DEC0[1].n14 DEC0[1].n13 0.663962
R306 DEC0[1].n15 DEC0[1].n14 0.663962
R307 DEC0[1] DEC0[1].n15 0.238481
R308 rseg_2_v3_0.v31.n0 rseg_2_v3_0.v31.t1 237.343
R309 rseg_2_v3_0.v31.n0 rseg_2_v3_0.v31.t2 10.6701
R310 rseg_2_v3_0.v31.t0 rseg_2_v3_0.v31.n0 10.5739
R311 a_4370_4223.n0 a_4370_4223.t2 251.719
R312 a_4370_4223.t0 a_4370_4223.n1 248.475
R313 a_4370_4223.n0 a_4370_4223.t1 241.631
R314 a_4370_4223.n1 a_4370_4223.t3 238.916
R315 a_4370_4223.n1 a_4370_4223.n0 3.24425
R316 DEC1[3].n2 DEC1[3].t3 213.218
R317 DEC1[3].n0 DEC1[3].t2 213.218
R318 DEC1[3].n2 DEC1[3].t1 212.554
R319 DEC1[3].n1 DEC1[3].t0 212.554
R320 DEC1[3].n0 DEC1[3].t4 212.554
R321 DEC1[3].n1 DEC1[3].n0 0.663962
R322 DEC1[3] DEC1[3].n1 0.457231
R323 DEC1[3] DEC1[3].n2 0.207231
R324 a_5474_4223.n0 a_5474_4223.t3 250.803
R325 a_5474_4223.n1 a_5474_4223.t1 248.238
R326 a_5474_4223.n0 a_5474_4223.t2 240.714
R327 a_5474_4223.t0 a_5474_4223.n1 239.833
R328 a_5474_4223.n1 a_5474_4223.n0 2.56508
R329 a_6452_6264.n2 a_6452_6264.t4 242.181
R330 a_6452_6264.n0 a_6452_6264.t1 240.082
R331 a_6452_6264.n0 a_6452_6264.t3 239.415
R332 a_6452_6264.n2 a_6452_6264.t5 239.248
R333 a_6452_6264.n1 a_6452_6264.t2 239.248
R334 a_6452_6264.t0 a_6452_6264.n3 239.248
R335 a_6452_6264.n1 a_6452_6264.n0 3.40883
R336 a_6452_6264.n3 a_6452_6264.n1 2.93383
R337 a_6452_6264.n3 a_6452_6264.n2 2.93383
R338 rseg_2_v3_0.v15.n0 rseg_2_v3_0.v15.t2 237.542
R339 rseg_2_v3_0.v15.n0 rseg_2_v3_0.v15.t1 10.5773
R340 rseg_2_v3_0.v15.t0 rseg_2_v3_0.v15.n0 10.577
R341 rseg_2_v3_0.v14 rseg_2_v3_0.v14.t2 237.291
R342 rseg_2_v3_0.v14.n0 rseg_2_v3_0.v14.t0 10.5327
R343 rseg_2_v3_0.v14.n0 rseg_2_v3_0.v14.t1 10.5285
R344 rseg_2_v3_0.v14 rseg_2_v3_0.v14.n0 0.941624
R345 DEC0[0].n0 DEC0[0].t11 213.218
R346 DEC0[0].n15 DEC0[0].t8 212.554
R347 DEC0[0].n14 DEC0[0].t5 212.554
R348 DEC0[0].n13 DEC0[0].t4 212.554
R349 DEC0[0].n12 DEC0[0].t3 212.554
R350 DEC0[0].n11 DEC0[0].t6 212.554
R351 DEC0[0].n10 DEC0[0].t0 212.554
R352 DEC0[0].n9 DEC0[0].t14 212.554
R353 DEC0[0].n8 DEC0[0].t2 212.554
R354 DEC0[0].n7 DEC0[0].t1 212.554
R355 DEC0[0].n6 DEC0[0].t15 212.554
R356 DEC0[0].n5 DEC0[0].t9 212.554
R357 DEC0[0].n4 DEC0[0].t13 212.554
R358 DEC0[0].n3 DEC0[0].t16 212.554
R359 DEC0[0].n2 DEC0[0].t10 212.554
R360 DEC0[0].n1 DEC0[0].t7 212.554
R361 DEC0[0].n0 DEC0[0].t12 212.554
R362 DEC0[0].n1 DEC0[0].n0 0.663962
R363 DEC0[0].n2 DEC0[0].n1 0.663962
R364 DEC0[0].n3 DEC0[0].n2 0.663962
R365 DEC0[0].n4 DEC0[0].n3 0.663962
R366 DEC0[0].n5 DEC0[0].n4 0.663962
R367 DEC0[0].n6 DEC0[0].n5 0.663962
R368 DEC0[0].n7 DEC0[0].n6 0.663962
R369 DEC0[0].n8 DEC0[0].n7 0.663962
R370 DEC0[0].n9 DEC0[0].n8 0.663962
R371 DEC0[0].n10 DEC0[0].n9 0.663962
R372 DEC0[0].n11 DEC0[0].n10 0.663962
R373 DEC0[0].n12 DEC0[0].n11 0.663962
R374 DEC0[0].n13 DEC0[0].n12 0.663962
R375 DEC0[0].n14 DEC0[0].n13 0.663962
R376 DEC0[0].n15 DEC0[0].n14 0.663962
R377 DEC0[0] DEC0[0].n15 0.209635
R378 rseg_2_v3_0.v2 rseg_2_v3_0.v2.t1 237.231
R379 rseg_2_v3_0.v2.n0 rseg_2_v3_0.v2.t0 10.6565
R380 rseg_2_v3_0.v2.n0 rseg_2_v3_0.v2.t2 10.5285
R381 rseg_2_v3_0.v2 rseg_2_v3_0.v2.n0 0.81529
R382 a_2438_4223.t0 a_2438_4223.n1 249.335
R383 a_2438_4223.n0 a_2438_4223.t1 247.23
R384 a_2438_4223.n0 a_2438_4223.t3 241.299
R385 a_2438_4223.n1 a_2438_4223.t2 239.248
R386 a_2438_4223.n1 a_2438_4223.n0 2.10675
R387 DEC0[2].n12 DEC0[2].t9 213.218
R388 DEC0[2].n0 DEC0[2].t13 213.218
R389 DEC0[2].n12 DEC0[2].t4 212.554
R390 DEC0[2].n13 DEC0[2].t12 212.554
R391 DEC0[2].n14 DEC0[2].t10 212.554
R392 DEC0[2].n11 DEC0[2].t5 212.554
R393 DEC0[2].n10 DEC0[2].t8 212.554
R394 DEC0[2].n9 DEC0[2].t7 212.554
R395 DEC0[2].n8 DEC0[2].t6 212.554
R396 DEC0[2].n7 DEC0[2].t3 212.554
R397 DEC0[2].n6 DEC0[2].t2 212.554
R398 DEC0[2].n5 DEC0[2].t0 212.554
R399 DEC0[2].n4 DEC0[2].t16 212.554
R400 DEC0[2].n3 DEC0[2].t14 212.554
R401 DEC0[2].n2 DEC0[2].t1 212.554
R402 DEC0[2].n1 DEC0[2].t11 212.554
R403 DEC0[2].n0 DEC0[2].t15 212.554
R404 DEC0[2].n1 DEC0[2].n0 0.663962
R405 DEC0[2].n2 DEC0[2].n1 0.663962
R406 DEC0[2].n3 DEC0[2].n2 0.663962
R407 DEC0[2].n4 DEC0[2].n3 0.663962
R408 DEC0[2].n5 DEC0[2].n4 0.663962
R409 DEC0[2].n6 DEC0[2].n5 0.663962
R410 DEC0[2].n7 DEC0[2].n6 0.663962
R411 DEC0[2].n8 DEC0[2].n7 0.663962
R412 DEC0[2].n9 DEC0[2].n8 0.663962
R413 DEC0[2].n10 DEC0[2].n9 0.663962
R414 DEC0[2].n11 DEC0[2].n10 0.663962
R415 DEC0[2].n14 DEC0[2].n13 0.663962
R416 DEC0[2].n13 DEC0[2].n12 0.663962
R417 DEC0[2] DEC0[2].n14 0.442808
R418 DEC0[2] DEC0[2].n11 0.221654
R419 rseg_2_v3_0.v43 rseg_2_v3_0.v43.t0 236.737
R420 rseg_2_v3_0.v43.n0 rseg_2_v3_0.v43.t1 10.7705
R421 rseg_2_v3_0.v43.n0 rseg_2_v3_0.v43.t2 10.7347
R422 rseg_2_v3_0.v43 rseg_2_v3_0.v43.n0 2.74678
R423 a_3818_4223.n0 a_3818_4223.t2 250.986
R424 a_3818_4223.n1 a_3818_4223.t1 249.524
R425 a_3818_4223.n0 a_3818_4223.t3 240.898
R426 a_3818_4223.t0 a_3818_4223.n1 239.649
R427 a_3818_4223.n1 a_3818_4223.n0 1.46092
R428 rseg_2_v3_0.v8 rseg_2_v3_0.v8.t0 236.044
R429 rseg_2_v3_0.v8.n0 rseg_2_v3_0.v8.t1 13.9493
R430 rseg_2_v3_0.v8.n0 rseg_2_v3_0.v8.t2 11.0147
R431 rseg_2_v3_0.v8 rseg_2_v3_0.v8.n0 4.72836
R432 a_3266_4223.n1 a_3266_4223.t3 250.435
R433 a_3266_4223.n0 a_3266_4223.t2 249.549
R434 a_3266_4223.n1 a_3266_4223.t4 240.347
R435 a_3266_4223.n0 a_3266_4223.t1 240.2
R436 a_3266_4223.t0 a_3266_4223.n2 240.2
R437 a_3266_4223.n2 a_3266_4223.n0 0.633833
R438 a_3266_4223.n2 a_3266_4223.n1 0.252583
R439 a_4646_4223.n0 a_4646_4223.t2 251.903
R440 a_4646_4223.n1 a_4646_4223.t1 248.659
R441 a_4646_4223.n0 a_4646_4223.t3 241.815
R442 a_4646_4223.t0 a_4646_4223.n1 238.732
R443 a_4646_4223.n1 a_4646_4223.n0 3.24425
R444 a_3542_4223.n0 a_3542_4223.t2 250.619
R445 a_3542_4223.n1 a_3542_4223.t1 249.733
R446 a_3542_4223.n0 a_3542_4223.t3 240.531
R447 a_3542_4223.t0 a_3542_4223.n1 240.016
R448 a_3542_4223.n1 a_3542_4223.n0 0.885917
R449 a_6176_6264.n0 a_6176_6264.t3 241.998
R450 a_6176_6264.n3 a_6176_6264.t4 239.899
R451 a_6176_6264.t0 a_6176_6264.n3 239.264
R452 a_6176_6264.n0 a_6176_6264.t5 239.065
R453 a_6176_6264.n1 a_6176_6264.t2 239.065
R454 a_6176_6264.n2 a_6176_6264.t1 239.065
R455 a_6176_6264.n2 a_6176_6264.n1 2.93383
R456 a_6176_6264.n1 a_6176_6264.n0 2.93383
R457 a_6176_6264.n3 a_6176_6264.n2 2.7755
R458 rseg_2_v3_0.v17.n0 rseg_2_v3_0.v17.t1 242.224
R459 rseg_2_v3_0.v17.t0 rseg_2_v3_0.v17.n0 10.7373
R460 rseg_2_v3_0.v17.n0 rseg_2_v3_0.v17.t2 10.5739
R461 rseg_2_v3_0.v18 rseg_2_v3_0.v18.t1 237.379
R462 rseg_2_v3_0.v18.n0 rseg_2_v3_0.v18.t2 10.5307
R463 rseg_2_v3_0.v18.n0 rseg_2_v3_0.v18.t0 10.5295
R464 rseg_2_v3_0.v18 rseg_2_v3_0.v18.n0 0.875827
R465 rseg_2_v3_0.v6 rseg_2_v3_0.v6.t1 236.447
R466 rseg_2_v3_0.v6.n0 rseg_2_v3_0.v6.t0 10.5383
R467 rseg_2_v3_0.v6.n0 rseg_2_v3_0.v6.t2 10.5285
R468 rseg_2_v3_0.v6 rseg_2_v3_0.v6.n0 3.74096
R469 a_2990_4223.t0 a_2990_4223.n1 250.069
R470 a_2990_4223.n0 a_2990_4223.t1 249.745
R471 a_2990_4223.n0 a_2990_4223.t3 240.565
R472 a_2990_4223.n1 a_2990_4223.t2 239.982
R473 a_2990_4223.n1 a_2990_4223.n0 0.323417
R474 rseg_2_v3_0.v45 rseg_2_v3_0.v45.t0 237.129
R475 rseg_2_v3_0.v45.n0 rseg_2_v3_0.v45.t2 10.7707
R476 rseg_2_v3_0.v45.n0 rseg_2_v3_0.v45.t1 10.7066
R477 rseg_2_v3_0.v45 rseg_2_v3_0.v45.n0 1.36863
R478 rseg_2_v3_0.v46 rseg_2_v3_0.v46.t1 237.683
R479 rseg_2_v3_0.v46.n0 rseg_2_v3_0.v46.t2 10.7345
R480 rseg_2_v3_0.v46.n0 rseg_2_v3_0.v46.t0 10.6569
R481 rseg_2_v3_0.v46 rseg_2_v3_0.v46.n0 0.688382
R482 DEC1[0].n2 DEC1[0].t1 213.218
R483 DEC1[0].n0 DEC1[0].t2 213.218
R484 DEC1[0].n2 DEC1[0].t0 212.554
R485 DEC1[0].n1 DEC1[0].t4 212.554
R486 DEC1[0].n0 DEC1[0].t3 212.554
R487 DEC1[0].n1 DEC1[0].n0 0.663962
R488 DEC1[0] DEC1[0].n2 0.363481
R489 DEC1[0] DEC1[0].n1 0.300981
R490 a_4094_4223.n0 a_4094_4223.t2 251.352
R491 a_4094_4223.n1 a_4094_4223.t1 248.684
R492 a_4094_4223.n0 a_4094_4223.t3 241.264
R493 a_4094_4223.t0 a_4094_4223.n1 239.282
R494 a_4094_4223.n1 a_4094_4223.n0 2.66925
R495 rseg_2_v3_0.v24 rseg_2_v3_0.v24.t0 236.203
R496 rseg_2_v3_0.v24.n0 rseg_2_v3_0.v24.t2 13.842
R497 rseg_2_v3_0.v24.n0 rseg_2_v3_0.v24.t1 10.7995
R498 rseg_2_v3_0.v24 rseg_2_v3_0.v24.n0 4.72836
R499 rseg_2_v3_0.v33.n0 rseg_2_v3_0.v33.t1 237.419
R500 rseg_2_v3_0.v33.n0 rseg_2_v3_0.v33.t2 10.6701
R501 rseg_2_v3_0.v33.t0 rseg_2_v3_0.v33.n0 10.5739
R502 rseg_2_v3_0.v34 rseg_2_v3_0.v34.t1 237.16
R503 rseg_2_v3_0.v34.n0 rseg_2_v3_0.v34.t0 10.7369
R504 rseg_2_v3_0.v34.n0 rseg_2_v3_0.v34.t2 10.6502
R505 rseg_2_v3_0.v34 rseg_2_v3_0.v34.n0 0.682179
R506 rseg_2_v3_0.v16.n0 rseg_2_v3_0.v16.t2 237.774
R507 rseg_2_v3_0.v16.n1 rseg_2_v3_0.v16.t1 237.685
R508 rseg_2_v3_0.v16.t0 rseg_2_v3_0.v16.n1 10.613
R509 rseg_2_v3_0.v16.n0 rseg_2_v3_0.v16.t3 10.612
R510 rseg_2_v3_0.v16.n1 rseg_2_v3_0.v16.n0 3.39554
R511 a_2162_4223.t0 a_2162_4223.n1 248.969
R512 a_2162_4223.n0 a_2162_4223.t1 246.287
R513 a_2162_4223.n0 a_2162_4223.t3 241.666
R514 a_2162_4223.n1 a_2162_4223.t2 238.881
R515 a_2162_4223.n1 a_2162_4223.n0 2.68175
R516 rseg_2_v3_0.v41 rseg_2_v3_0.v41.t1 236.345
R517 rseg_2_v3_0.v41.n0 rseg_2_v3_0.v41.t0 10.7937
R518 rseg_2_v3_0.v41.n0 rseg_2_v3_0.v41.t2 10.6741
R519 rseg_2_v3_0.v41 rseg_2_v3_0.v41.n0 4.095
R520 rseg_2_v3_0.v22 rseg_2_v3_0.v22.t1 236.595
R521 rseg_2_v3_0.v22.n0 rseg_2_v3_0.v22.t0 10.5306
R522 rseg_2_v3_0.v22.n0 rseg_2_v3_0.v22.t2 10.5285
R523 rseg_2_v3_0.v22 rseg_2_v3_0.v22.n0 3.54826
R524 rseg_2_v3_0.v27 rseg_2_v3_0.v27.t1 236.52
R525 rseg_2_v3_0.v27.n0 rseg_2_v3_0.v27.t2 10.763
R526 rseg_2_v3_0.v27.n0 rseg_2_v3_0.v27.t0 10.7161
R527 rseg_2_v3_0.v27 rseg_2_v3_0.v27.n0 2.72817
R528 rseg_2_v3_0.v1.n0 rseg_2_v3_0.v1.t1 240.27
R529 rseg_2_v3_0.v1.n0 rseg_2_v3_0.v1.t2 10.7145
R530 rseg_2_v3_0.v1.t0 rseg_2_v3_0.v1.n0 10.5739
R531 a_1886_4223.n0 a_1886_4223.t1 249.153
R532 a_1886_4223.n1 a_1886_4223.t2 247.62
R533 a_1886_4223.t0 a_1886_4223.n1 241.482
R534 a_1886_4223.n0 a_1886_4223.t3 239.065
R535 a_1886_4223.n1 a_1886_4223.n0 1.53175
R536 rseg_2_v3_0.v40.n0 rseg_2_v3_0.v40.t1 240.804
R537 rseg_2_v3_0.v40.t0 rseg_2_v3_0.v40.n0 13.9465
R538 rseg_2_v3_0.v40.n0 rseg_2_v3_0.v40.t2 10.7604
R539 DEC1[1].n0 DEC1[1].t0 213.218
R540 DEC1[1] DEC1[1].t2 212.989
R541 DEC1[1].n2 DEC1[1].t4 212.554
R542 DEC1[1].n1 DEC1[1].t3 212.554
R543 DEC1[1].n0 DEC1[1].t1 212.554
R544 DEC1[1].n1 DEC1[1].n0 0.663962
R545 DEC1[1].n2 DEC1[1].n1 0.663962
R546 DEC1[1] DEC1[1].n2 0.228865
R547 a_2714_4223.n0 a_2714_4223.t1 249.702
R548 a_2714_4223.n2 a_2714_4223.t2 248.171
R549 a_2714_4223.n1 a_2714_4223.t4 240.933
R550 a_2714_4223.t0 a_2714_4223.n2 240.933
R551 a_2714_4223.n0 a_2714_4223.t3 239.614
R552 a_2714_4223.n1 a_2714_4223.n0 0.898417
R553 a_2714_4223.n2 a_2714_4223.n1 0.633833
R554 a_7004_6264.n0 a_7004_6264.t4 244.489
R555 a_7004_6264.n2 a_7004_6264.t3 242.548
R556 a_7004_6264.n1 a_7004_6264.t1 239.614
R557 a_7004_6264.n0 a_7004_6264.t2 239.614
R558 a_7004_6264.t0 a_7004_6264.n2 239.614
R559 a_7004_6264.n1 a_7004_6264.n0 2.93383
R560 a_7004_6264.n2 a_7004_6264.n1 2.93383
R561 a_5198_4223.n0 a_5198_4223.t2 251.168
R562 a_5198_4223.n2 a_5198_4223.t3 250.329
R563 a_5198_4223.n0 a_5198_4223.t4 241.082
R564 a_5198_4223.n1 a_5198_4223.t1 239.465
R565 a_5198_4223.t0 a_5198_4223.n2 239.465
R566 a_5198_4223.n2 a_5198_4223.n1 0.633833
R567 a_5198_4223.n1 a_5198_4223.n0 0.20675
R568 a_5900_6264.n0 a_5900_6264.t3 241.857
R569 a_5900_6264.n1 a_5900_6264.t2 241.815
R570 a_5900_6264.n1 a_5900_6264.t4 238.881
R571 a_5900_6264.n0 a_5900_6264.t1 238.881
R572 a_5900_6264.t0 a_5900_6264.n2 238.881
R573 a_5900_6264.n2 a_5900_6264.n0 2.93383
R574 a_5900_6264.n2 a_5900_6264.n1 2.93383
R575 rseg_2_v3_0.v44 rseg_2_v3_0.v44.t0 237.291
R576 rseg_2_v3_0.v44.n0 rseg_2_v3_0.v44.t2 10.7254
R577 rseg_2_v3_0.v44.n0 rseg_2_v3_0.v44.t1 10.6855
R578 rseg_2_v3_0.v44 rseg_2_v3_0.v44.n0 2.06796
R579 rseg_2_v3_0.v13 rseg_2_v3_0.v13.t2 237.06
R580 rseg_2_v3_0.v13.n0 rseg_2_v3_0.v13.t1 10.5763
R581 rseg_2_v3_0.v13.n0 rseg_2_v3_0.v13.t0 10.5739
R582 rseg_2_v3_0.v13 rseg_2_v3_0.v13.n0 1.61086
R583 rseg_2_v3_0.v12 rseg_2_v3_0.v12.t1 236.899
R584 rseg_2_v3_0.v12.n0 rseg_2_v3_0.v12.t0 10.5327
R585 rseg_2_v3_0.v12.n0 rseg_2_v3_0.v12.t2 10.5285
R586 rseg_2_v3_0.v12 rseg_2_v3_0.v12.n0 2.18861
R587 DEC2[3] DEC2[3].t0 212.907
R588 DEC2[3] DEC2[3].t1 212.864
R589 VH.n0 VH.t1 244.607
R590 VH VH.t0 239.375
R591 VH.n1 VH.t2 239.264
R592 VH.n0 VH.t3 234.399
R593 VH.n1 VH.n0 6.0755
R594 VH VH.n1 1.09842
R595 rseg_2_v3_0.v20 rseg_2_v3_0.v20.t1 236.987
R596 rseg_2_v3_0.v20.n0 rseg_2_v3_0.v20.t2 10.6247
R597 rseg_2_v3_0.v20.n0 rseg_2_v3_0.v20.t0 10.5295
R598 rseg_2_v3_0.v20 rseg_2_v3_0.v20.n0 2.10756
R599 rseg_2_v3_0.v37 rseg_2_v3_0.v37.t1 236.597
R600 rseg_2_v3_0.v37.n0 rseg_2_v3_0.v37.t0 10.7609
R601 rseg_2_v3_0.v37.n0 rseg_2_v3_0.v37.t2 10.7147
R602 rseg_2_v3_0.v37 rseg_2_v3_0.v37.n0 2.72245
R603 a_1334_4223.n0 a_1334_4223.t1 249.886
R604 a_1334_4223.t0 a_1334_4223.n1 247.333
R605 a_1334_4223.n1 a_1334_4223.t2 240.75
R606 a_1334_4223.n0 a_1334_4223.t3 239.798
R607 a_1334_4223.n1 a_1334_4223.n0 2.55258
R608 rseg_2_v3_0.v25 rseg_2_v3_0.v25.t0 236.129
R609 rseg_2_v3_0.v25.n0 rseg_2_v3_0.v25.t1 10.8275
R610 rseg_2_v3_0.v25.n0 rseg_2_v3_0.v25.t2 10.6741
R611 rseg_2_v3_0.v25 rseg_2_v3_0.v25.n0 4.11253
R612 rseg_2_v3_0.v26 rseg_2_v3_0.v26.t0 236.433
R613 rseg_2_v3_0.v26.n0 rseg_2_v3_0.v26.t2 10.7826
R614 rseg_2_v3_0.v26.n0 rseg_2_v3_0.v26.t1 10.6321
R615 rseg_2_v3_0.v26 rseg_2_v3_0.v26.n0 3.43753
R616 rseg_2_v3_0.v32.n0 rseg_2_v3_0.v32.t3 237.611
R617 rseg_2_v3_0.v32.n1 rseg_2_v3_0.v32.t2 237.554
R618 rseg_2_v3_0.v32.t0 rseg_2_v3_0.v32.n1 10.613
R619 rseg_2_v3_0.v32.n0 rseg_2_v3_0.v32.t1 10.612
R620 rseg_2_v3_0.v32.n1 rseg_2_v3_0.v32.n0 3.36262
R621 rseg_2_v3_0.v3 rseg_2_v3_0.v3.t2 239.756
R622 rseg_2_v3_0.v3.n0 rseg_2_v3_0.v3.t1 10.5893
R623 rseg_2_v3_0.v3.n0 rseg_2_v3_0.v3.t0 10.5739
R624 rseg_2_v3_0.v3 rseg_2_v3_0.v3.n0 1.55408
R625 rseg_2_v3_0.v38 rseg_2_v3_0.v38.t2 236.376
R626 rseg_2_v3_0.v38.n0 rseg_2_v3_0.v38.t0 10.7194
R627 rseg_2_v3_0.v38.n0 rseg_2_v3_0.v38.t1 10.686
R628 rseg_2_v3_0.v38 rseg_2_v3_0.v38.n0 3.41844
R629 a_1610_4223.n0 a_1610_4223.t2 249.518
R630 a_1610_4223.n1 a_1610_4223.t1 249.325
R631 a_1610_4223.t0 a_1610_4223.n1 241.115
R632 a_1610_4223.n0 a_1610_4223.t3 239.431
R633 a_1610_4223.n1 a_1610_4223.n0 0.19425
R634 a_6728_6264.n0 a_6728_6264.t4 242.364
R635 a_6728_6264.t0 a_6728_6264.n3 240.264
R636 a_6728_6264.n3 a_6728_6264.t1 239.631
R637 a_6728_6264.n0 a_6728_6264.t5 239.431
R638 a_6728_6264.n1 a_6728_6264.t2 239.431
R639 a_6728_6264.n2 a_6728_6264.t3 239.431
R640 a_6728_6264.n3 a_6728_6264.n2 4.04217
R641 a_6728_6264.n2 a_6728_6264.n1 2.93383
R642 a_6728_6264.n1 a_6728_6264.n0 2.93383
R643 rseg_2_v3_0.v39 rseg_2_v3_0.v39.t1 236.206
R644 rseg_2_v3_0.v39.n0 rseg_2_v3_0.v39.t2 10.7562
R645 rseg_2_v3_0.v39.n0 rseg_2_v3_0.v39.t0 10.7314
R646 rseg_2_v3_0.v39 rseg_2_v3_0.v39.n0 4.09296
R647 rseg_2_v3_0.v9 rseg_2_v3_0.v9.t1 236.276
R648 rseg_2_v3_0.v9.n0 rseg_2_v3_0.v9.t0 10.5784
R649 rseg_2_v3_0.v9.n0 rseg_2_v3_0.v9.t2 10.5739
R650 rseg_2_v3_0.v9 rseg_2_v3_0.v9.n0 4.16334
R651 rseg_2_v3_0.v10 rseg_2_v3_0.v10.t1 236.507
R652 rseg_2_v3_0.v10.n0 rseg_2_v3_0.v10.t2 10.5328
R653 rseg_2_v3_0.v10.n0 rseg_2_v3_0.v10.t0 10.5295
R654 rseg_2_v3_0.v10 rseg_2_v3_0.v10.n0 3.49115
R655 rseg_2_v3_0.v7 rseg_2_v3_0.v7.t1 238.972
R656 rseg_2_v3_0.v7.n0 rseg_2_v3_0.v7.t2 10.5816
R657 rseg_2_v3_0.v7.n0 rseg_2_v3_0.v7.t0 10.5739
R658 rseg_2_v3_0.v7 rseg_2_v3_0.v7.n0 4.43733
R659 VL.n0 VL.t2 240.29
R660 VL VL.t0 239.346
R661 VL.n0 VL.t3 239.082
R662 VL.n1 VL.t1 239.082
R663 VL.n1 VL.n0 1.20883
R664 VL VL.n1 0.94425
R665 V0.n0 V0.t1 237.625
R666 V0.n0 V0.t0 10.612
R667 V0 V0.n0 2.7443
R668 DEC2[1] DEC2[1].t1 212.899
R669 DEC2[1] DEC2[1].t0 212.875
R670 rseg_2_v3_0.v36 rseg_2_v3_0.v36.t0 236.768
R671 rseg_2_v3_0.v36.n0 rseg_2_v3_0.v36.t2 10.7131
R672 rseg_2_v3_0.v36.n0 rseg_2_v3_0.v36.t1 10.6688
R673 rseg_2_v3_0.v36 rseg_2_v3_0.v36.n0 2.05079
R674 rseg_2_v3_0.v5 rseg_2_v3_0.v5.t1 239.363
R675 rseg_2_v3_0.v5.n0 rseg_2_v3_0.v5.t2 10.5837
R676 rseg_2_v3_0.v5.n0 rseg_2_v3_0.v5.t0 10.5739
R677 rseg_2_v3_0.v5 rseg_2_v3_0.v5.n0 3.00616
R678 a_4922_4223.n0 a_4922_4223.t2 251.536
R679 a_4922_4223.n1 a_4922_4223.t1 250.017
R680 a_4922_4223.n0 a_4922_4223.t3 241.447
R681 a_4922_4223.t0 a_4922_4223.n1 239.1
R682 a_4922_4223.n1 a_4922_4223.n0 1.51925
R683 rseg_2_v3_0.v23 rseg_2_v3_0.v23.t1 236.137
R684 rseg_2_v3_0.v23.n0 rseg_2_v3_0.v23.t2 10.6507
R685 rseg_2_v3_0.v23.n0 rseg_2_v3_0.v23.t0 10.6439
R686 rseg_2_v3_0.v23 rseg_2_v3_0.v23.n0 4.1755
R687 a_1058_4223.n0 a_1058_4223.t2 250.252
R688 a_1058_4223.t0 a_1058_4223.n1 245.975
R689 a_1058_4223.n1 a_1058_4223.t1 240.382
R690 a_1058_4223.n0 a_1058_4223.t3 240.165
R691 a_1058_4223.n1 a_1058_4223.n0 4.27758
R692 rseg_2_v3_0.v4 rseg_2_v3_0.v4.t2 236.839
R693 rseg_2_v3_0.v4.n0 rseg_2_v3_0.v4.t0 10.5428
R694 rseg_2_v3_0.v4.n0 rseg_2_v3_0.v4.t1 10.5285
R695 rseg_2_v3_0.v4 rseg_2_v3_0.v4.n0 2.30299
R696 rseg_2_v3_0.v21 rseg_2_v3_0.v21.t0 236.529
R697 rseg_2_v3_0.v21.n0 rseg_2_v3_0.v21.t1 10.8508
R698 rseg_2_v3_0.v21.n0 rseg_2_v3_0.v21.t2 10.6202
R699 rseg_2_v3_0.v21 rseg_2_v3_0.v21.n0 2.7508
R700 rseg_2_v3_0.v11 rseg_2_v3_0.v11.t0 236.668
R701 rseg_2_v3_0.v11.n0 rseg_2_v3_0.v11.t2 10.5784
R702 rseg_2_v3_0.v11.n0 rseg_2_v3_0.v11.t1 10.5739
R703 rseg_2_v3_0.v11 rseg_2_v3_0.v11.n0 2.86211
R704 rseg_2_v3_0.v35 rseg_2_v3_0.v35.t1 236.988
R705 rseg_2_v3_0.v35.n0 rseg_2_v3_0.v35.t2 10.7851
R706 rseg_2_v3_0.v35.n0 rseg_2_v3_0.v35.t0 10.6941
R707 rseg_2_v3_0.v35 rseg_2_v3_0.v35.n0 1.35575
R708 rseg_2_v3_0.v19 rseg_2_v3_0.v19.t1 236.921
R709 rseg_2_v3_0.v19 rseg_2_v3_0.v19.n0 11.7546
R710 rseg_2_v3_0.v19.n0 rseg_2_v3_0.v19.t0 10.7127
R711 rseg_2_v3_0.v19.n0 rseg_2_v3_0.v19.t2 10.5739
R712 DEC2[2] DEC2[2].t0 212.887
R713 DEC2[2] DEC2[2].t1 212.887
R714 rseg_2_v3_0.v29 rseg_2_v3_0.v29.t2 236.911
R715 rseg_2_v3_0.v29.n0 rseg_2_v3_0.v29.t0 10.779
R716 rseg_2_v3_0.v29.n0 rseg_2_v3_0.v29.t1 10.6965
R717 rseg_2_v3_0.v29 rseg_2_v3_0.v29.n0 1.35861
R718 rseg_2_v3_0.v30 rseg_2_v3_0.v30.t1 237.215
R719 rseg_2_v3_0.v30.n0 rseg_2_v3_0.v30.t0 10.7421
R720 rseg_2_v3_0.v30.n0 rseg_2_v3_0.v30.t2 10.6502
R721 rseg_2_v3_0.v30 rseg_2_v3_0.v30.n0 0.682179
R722 DEC1[2].n0 DEC1[2].t0 213.218
R723 DEC1[2] DEC1[2].t1 212.982
R724 DEC1[2].n2 DEC1[2].t4 212.554
R725 DEC1[2].n1 DEC1[2].t3 212.554
R726 DEC1[2].n0 DEC1[2].t2 212.554
R727 DEC1[2].n1 DEC1[2].n0 0.663962
R728 DEC1[2].n2 DEC1[2].n1 0.663962
R729 DEC1[2] DEC1[2].n2 0.236077
R730 rseg_2_v3_0.v28 rseg_2_v3_0.v28.t2 236.825
R731 rseg_2_v3_0.v28.n0 rseg_2_v3_0.v28.t0 10.7162
R732 rseg_2_v3_0.v28.n0 rseg_2_v3_0.v28.t1 10.6741
R733 rseg_2_v3_0.v28 rseg_2_v3_0.v28.n0 2.05317
R734 rseg_2_v3_0.v42 rseg_2_v3_0.v42.t0 236.899
R735 rseg_2_v3_0.v42.n0 rseg_2_v3_0.v42.t2 10.7518
R736 rseg_2_v3_0.v42.n0 rseg_2_v3_0.v42.t1 10.6292
R737 rseg_2_v3_0.v42 rseg_2_v3_0.v42.n0 3.42215
R738 DEC2[0] DEC2[0].t1 212.895
R739 DEC2[0] DEC2[0].t0 212.876
C0 DEC0[0] V0 0.12956f
C1 VL DEC2[0] 0.14256f
C2 rseg_2_v3_0.v2 rseg_2_v3_0.v4 1.57718f
C3 rseg_2_v3_0.v37 rseg_2_v3_0.v39 2.25141f
C4 rseg_2_v3_0.v10 rseg_2_v3_0.v21 0.02734f
C5 rseg_2_v3_0.v44 V48 0.12159f
C6 rseg_2_v3_0.v13 rseg_2_v3_0.v4 0.01528f
C7 DEC0[0] rseg_2_v3_0.v6 0.05852f
C8 rseg_2_v3_0.v25 rseg_2_v3_0.v27 2.23765f
C9 rseg_2_v3_0.v20 rseg_2_v3_0.v18 1.68518f
C10 VL DEC2[3] 0.14124f
C11 DEC0[1] DEC0[2] 0.01836f
C12 rseg_2_v3_0.v42 rseg_2_v3_0.v44 2.28703f
C13 rseg_2_v3_0.v14 rseg_2_v3_0.v13 0.01875f
C14 rseg_2_v3_0.v12 rseg_2_v3_0.v10 1.96915f
C15 rseg_2_v3_0.v39 rseg_2_v3_0.v38 0.01848f
C16 rseg_2_v3_0.v5 DEC0[0] 0.05702f
C17 rseg_2_v3_0.v22 rseg_2_v3_0.v21 0.01929f
C18 DEC1[0] DEC1[3] 0.04353f
C19 rseg_2_v3_0.v37 rseg_2_v3_0.v38 0.01848f
C20 DEC2[1] VH 0.24374f
C21 rseg_2_v3_0.v11 DEC0[0] 0.05997f
C22 rseg_2_v3_0.v27 rseg_2_v3_0.v24 0.01605f
C23 rseg_2_v3_0.v9 rseg_2_v3_0.v10 0.01515f
C24 rseg_2_v3_0.v25 rseg_2_v3_0.v22 0.02066f
C25 rseg_2_v3_0.v36 DEC0[2] 0.05483f
C26 rseg_2_v3_0.v14 rseg_2_v3_0.v12 1.71248f
C27 rseg_2_v3_0.v27 rseg_2_v3_0.v20 0.02097f
C28 rseg_2_v3_0.v6 rseg_2_v3_0.v8 2.21718f
C29 DEC2[2] DEC2[3] 0.043f
C30 rseg_2_v3_0.v21 rseg_2_v3_0.v19 1.80576f
C31 DEC0[1] rseg_2_v3_0.v26 0.06616f
C32 VL VH 1.06154f
C33 rseg_2_v3_0.v45 DEC0[2] 0.0556f
C34 rseg_2_v3_0.v28 rseg_2_v3_0.v37 0.02568f
C35 rseg_2_v3_0.v41 rseg_2_v3_0.v43 2.32271f
C36 rseg_2_v3_0.v38 rseg_2_v3_0.v43 0.01984f
C37 rseg_2_v3_0.v2 DEC0[0] 0.05143f
C38 DEC1[2] DEC1[3] 0.04353f
C39 rseg_2_v3_0.v35 rseg_2_v3_0.v34 0.01927f
C40 rseg_2_v3_0.v44 DEC0[2] 0.05869f
C41 DEC0[1] rseg_2_v3_0.v29 0.05523f
C42 rseg_2_v3_0.v22 rseg_2_v3_0.v24 2.25734f
C43 rseg_2_v3_0.v38 rseg_2_v3_0.v41 0.01944f
C44 DEC2[2] VH 0.08999f
C45 rseg_2_v3_0.v7 DEC0[0] 0.03198f
C46 rseg_2_v3_0.v13 DEC0[0] 0.05597f
C47 rseg_2_v3_0.v22 rseg_2_v3_0.v20 1.96543f
C48 rseg_2_v3_0.v11 rseg_2_v3_0.v8 0.01317f
C49 rseg_2_v3_0.v45 rseg_2_v3_0.v36 0.02014f
C50 rseg_2_v3_0.v12 rseg_2_v3_0.v19 0.02582f
C51 rseg_2_v3_0.v5 V0 0.12611f
C52 DEC1[0] DEC2[0] 0.01817f
C53 VL DEC2[1] 0.08984f
C54 rseg_2_v3_0.v20 rseg_2_v3_0.v19 0.0191f
C55 rseg_2_v3_0.v10 rseg_2_v3_0.v23 1.77186f
C56 rseg_2_v3_0.v12 DEC0[0] 0.06103f
C57 rseg_2_v3_0.v5 rseg_2_v3_0.v6 0.01252f
C58 rseg_2_v3_0.v45 rseg_2_v3_0.v44 0.01616f
C59 DEC0[1] rseg_2_v3_0.v21 0.05959f
C60 rseg_2_v3_0.v9 DEC0[0] 0.04881f
C61 rseg_2_v3_0.v11 rseg_2_v3_0.v6 0.0142f
C62 rseg_2_v3_0.v2 V0 1.49083f
C63 rseg_2_v3_0.v7 rseg_2_v3_0.v8 0.01396f
C64 rseg_2_v3_0.v37 rseg_2_v3_0.v35 1.92248f
C65 DEC2[2] DEC2[1] 0.043f
C66 rseg_2_v3_0.v25 DEC0[1] 0.03841f
C67 VL DEC2[2] 0.19606f
C68 rseg_2_v3_0.v7 V0 0.15536f
C69 rseg_2_v3_0.v28 rseg_2_v3_0.v30 1.81252f
C70 rseg_2_v3_0.v22 rseg_2_v3_0.v23 0.02114f
C71 rseg_2_v3_0.v3 DEC0[0] 0.05382f
C72 DEC0[2] rseg_2_v3_0.v34 0.05127f
C73 rseg_2_v3_0.v28 rseg_2_v3_0.v27 0.01966f
C74 rseg_2_v3_0.v25 rseg_2_v3_0.v26 0.01965f
C75 rseg_2_v3_0.v46 V48 1.72319f
C76 DEC0[1] rseg_2_v3_0.v24 0.06816f
C77 rseg_2_v3_0.v7 rseg_2_v3_0.v6 0.01326f
C78 rseg_2_v3_0.v9 rseg_2_v3_0.v8 2.60553f
C79 rseg_2_v3_0.v20 DEC0[1] 0.0549f
C80 rseg_2_v3_0.v42 rseg_2_v3_0.v43 0.01692f
C81 rseg_2_v3_0.v36 rseg_2_v3_0.v34 1.75263f
C82 rseg_2_v3_0.v24 rseg_2_v3_0.v26 0.55358f
C83 rseg_2_v3_0.v45 rseg_2_v3_0.v34 0.02043f
C84 rseg_2_v3_0.v42 rseg_2_v3_0.v41 0.0174f
C85 rseg_2_v3_0.v7 rseg_2_v3_0.v5 2.80645f
C86 rseg_2_v3_0.v28 rseg_2_v3_0.v35 0.02519f
C87 rseg_2_v3_0.v39 DEC0[2] 0.03198f
C88 rseg_2_v3_0.v13 rseg_2_v3_0.v11 1.82582f
C89 rseg_2_v3_0.v18 rseg_2_v3_0.v19 0.02053f
C90 rseg_2_v3_0.v37 DEC0[2] 0.05934f
C91 rseg_2_v3_0.v9 rseg_2_v3_0.v6 0.01391f
C92 rseg_2_v3_0.v3 V0 0.1393f
C93 rseg_2_v3_0.v35 rseg_2_v3_0.v30 0.02497f
C94 rseg_2_v3_0.v22 rseg_2_v3_0.v27 0.02063f
C95 rseg_2_v3_0.v20 rseg_2_v3_0.v29 0.02078f
C96 rseg_2_v3_0.v23 rseg_2_v3_0.v8 0.05599f
C97 rseg_2_v3_0.v12 rseg_2_v3_0.v11 0.01623f
C98 rseg_2_v3_0.v13 rseg_2_v3_0.v2 0.01634f
C99 rseg_2_v3_0.v39 rseg_2_v3_0.v26 1.82529f
C100 DEC1[1] DEC1[2] 0.04353f
C101 DEC0[2] rseg_2_v3_0.v43 0.06041f
C102 rseg_2_v3_0.v37 rseg_2_v3_0.v26 0.02587f
C103 rseg_2_v3_0.v46 DEC0[2] 0.05546f
C104 DEC0[1] rseg_2_v3_0.v23 0.03299f
C105 rseg_2_v3_0.v37 rseg_2_v3_0.v36 0.01886f
C106 DEC0[0] rseg_2_v3_0.v4 0.0547f
C107 rseg_2_v3_0.v9 rseg_2_v3_0.v11 2.09225f
C108 rseg_2_v3_0.v10 DEC0[0] 0.06502f
C109 DEC0[2] rseg_2_v3_0.v41 0.05928f
C110 rseg_2_v3_0.v14 rseg_2_v3_0.v19 0.02577f
C111 rseg_2_v3_0.v38 DEC0[2] 0.05789f
C112 rseg_2_v3_0.v12 rseg_2_v3_0.v21 0.02654f
C113 rseg_2_v3_0.v5 rseg_2_v3_0.v3 2.48553f
C114 rseg_2_v3_0.v36 rseg_2_v3_0.v43 0.01986f
C115 rseg_2_v3_0.v20 rseg_2_v3_0.v21 0.02084f
C116 rseg_2_v3_0.v14 DEC0[0] 0.05687f
C117 rseg_2_v3_0.v12 rseg_2_v3_0.v13 0.01833f
C118 rseg_2_v3_0.v25 rseg_2_v3_0.v24 2.91357f
C119 rseg_2_v3_0.v45 rseg_2_v3_0.v43 1.98281f
C120 DEC0[1] rseg_2_v3_0.v18 0.05194f
C121 rseg_2_v3_0.v45 rseg_2_v3_0.v46 0.01575f
C122 rseg_2_v3_0.v28 DEC0[1] 0.06133f
C123 rseg_2_v3_0.v36 rseg_2_v3_0.v38 2.07263f
C124 rseg_2_v3_0.v10 rseg_2_v3_0.v8 0.53808f
C125 rseg_2_v3_0.v42 V48 0.15466f
C126 rseg_2_v3_0.v44 rseg_2_v3_0.v43 0.01659f
C127 rseg_2_v3_0.v44 rseg_2_v3_0.v46 1.94305f
C128 DEC0[1] rseg_2_v3_0.v30 0.05675f
C129 rseg_2_v3_0.v28 rseg_2_v3_0.v26 2.13767f
C130 rseg_2_v3_0.v4 V0 0.01681f
C131 rseg_2_v3_0.v27 DEC0[1] 0.05989f
C132 rseg_2_v3_0.v29 rseg_2_v3_0.v18 0.02109f
C133 rseg_2_v3_0.v28 rseg_2_v3_0.v29 0.01992f
C134 rseg_2_v3_0.v6 rseg_2_v3_0.v4 1.90109f
C135 DEC2[0] VH 0.10669f
C136 rseg_2_v3_0.v21 rseg_2_v3_0.v23 2.08874f
C137 rseg_2_v3_0.v27 rseg_2_v3_0.v26 0.0199f
C138 rseg_2_v3_0.v35 DEC0[2] 0.05522f
C139 rseg_2_v3_0.v22 DEC0[1] 0.06054f
C140 rseg_2_v3_0.v39 rseg_2_v3_0.v24 0.07044f
C141 DEC0[2] V48 0.05661f
C142 rseg_2_v3_0.v29 rseg_2_v3_0.v30 0.01993f
C143 rseg_2_v3_0.v5 rseg_2_v3_0.v4 0.01178f
C144 rseg_2_v3_0.v27 rseg_2_v3_0.v29 1.90818f
C145 DEC0[1] rseg_2_v3_0.v19 0.05518f
C146 rseg_2_v3_0.v11 rseg_2_v3_0.v4 0.01456f
C147 DEC2[3] VH 0.13063f
C148 rseg_2_v3_0.v42 DEC0[2] 0.06502f
C149 rseg_2_v3_0.v10 rseg_2_v3_0.v11 0.01566f
C150 DEC0[0] rseg_2_v3_0.v8 0.05056f
C151 rseg_2_v3_0.v36 rseg_2_v3_0.v35 0.01906f
C152 rseg_2_v3_0.v24 rseg_2_v3_0.v23 0.01963f
C153 DEC2[1] DEC2[0] 0.043f
C154 DEC0[1] DEC0[0] 0.01836f
C155 V48 GND 1.56118f
C156 DEC0[2] GND 5.41185f
C157 DEC0[1] GND 5.13285f
C158 V0 GND 2.40947f
C159 DEC0[0] GND 5.27522f
C160 VH GND 0.68034f
C161 VL GND 0.46529f
C162 DEC2[3] GND 0.60863f
C163 DEC2[2] GND 0.57813f
C164 DEC2[1] GND 0.57115f
C165 DEC2[0] GND 0.59373f
C166 DEC1[0] GND 1.4667f
C167 DEC1[3] GND 1.45153f
C168 DEC1[2] GND 1.46452f
C169 DEC1[1] GND 1.52774f
C170 rseg_2_v3_0.v42 GND 2.1743f
C171 rseg_2_v3_0.v44 GND 1.32207f
C172 rseg_2_v3_0.v46 GND 0.91672f
C173 rseg_2_v3_0.v45 GND 0.89932f
C174 rseg_2_v3_0.v43 GND 1.26475f
C175 rseg_2_v3_0.v41 GND 2.16252f
C176 rseg_2_v3_0.v38 GND 1.52048f
C177 rseg_2_v3_0.v36 GND 1.1614f
C178 rseg_2_v3_0.v34 GND 0.82727f
C179 rseg_2_v3_0.v35 GND 0.82365f
C180 rseg_2_v3_0.v37 GND 1.18969f
C181 rseg_2_v3_0.v39 GND 1.76674f
C182 rseg_2_v3_0.v26 GND 1.23612f
C183 rseg_2_v3_0.v28 GND 1.15392f
C184 rseg_2_v3_0.v30 GND 0.80858f
C185 rseg_2_v3_0.v29 GND 0.83077f
C186 rseg_2_v3_0.v27 GND 1.17794f
C187 rseg_2_v3_0.v25 GND 2.04014f
C188 rseg_2_v3_0.v24 GND 2.98762f
C189 rseg_2_v3_0.v22 GND 1.32334f
C190 rseg_2_v3_0.v20 GND 0.9106f
C191 rseg_2_v3_0.v18 GND 0.84609f
C192 rseg_2_v3_0.v19 GND 0.8303f
C193 rseg_2_v3_0.v21 GND 1.17765f
C194 rseg_2_v3_0.v23 GND 1.75309f
C195 rseg_2_v3_0.v10 GND 0.81139f
C196 rseg_2_v3_0.v12 GND 0.89682f
C197 rseg_2_v3_0.v14 GND 0.82563f
C198 rseg_2_v3_0.v13 GND 0.85946f
C199 rseg_2_v3_0.v11 GND 1.25295f
C200 rseg_2_v3_0.v9 GND 2.09094f
C201 rseg_2_v3_0.v8 GND 3.30542f
C202 rseg_2_v3_0.v6 GND 1.56789f
C203 rseg_2_v3_0.v4 GND 1.20222f
C204 rseg_2_v3_0.v2 GND 1.12435f
C205 rseg_2_v3_0.v3 GND 2.25075f
C206 rseg_2_v3_0.v5 GND 2.40032f
C207 rseg_2_v3_0.v7 GND 3.45704f
C208 rseg_2_v3_0.v42.t0 GND 0.01054f
C209 rseg_2_v3_0.v42.t1 GND 0.09055f
C210 rseg_2_v3_0.v42.t2 GND 0.10014f
C211 rseg_2_v3_0.v42.n0 GND 1.78741f
C212 rseg_2_v3_0.v28.t2 GND 0.01099f
C213 rseg_2_v3_0.v28.t1 GND 0.09795f
C214 rseg_2_v3_0.v28.t0 GND 0.10095f
C215 rseg_2_v3_0.v28.n0 GND 1.61052f
C216 rseg_2_v3_0.v11.t0 GND 0.01146f
C217 rseg_2_v3_0.v11.t2 GND 0.09471f
C218 rseg_2_v3_0.v11.t1 GND 0.09441f
C219 rseg_2_v3_0.v11.n0 GND 1.58504f
C220 rseg_2_v3_0.v21.t0 GND 0.01097f
C221 rseg_2_v3_0.v21.t2 GND 0.09398f
C222 rseg_2_v3_0.v21.t1 GND 0.10876f
C223 rseg_2_v3_0.v21.n0 GND 1.59653f
C224 a_1058_4223.t2 GND 0.15594f
C225 a_1058_4223.t3 GND 0.06377f
C226 a_1058_4223.n0 GND 5.11593f
C227 a_1058_4223.t1 GND 0.06506f
C228 a_1058_4223.n1 GND 3.89706f
C229 a_1058_4223.t0 GND 0.10224f
C230 rseg_2_v3_0.v23.t1 GND 0.01006f
C231 rseg_2_v3_0.v23.t2 GND 0.09028f
C232 rseg_2_v3_0.v23.t0 GND 0.08989f
C233 rseg_2_v3_0.v23.n0 GND 1.61436f
C234 a_4922_4223.t1 GND 0.1673f
C235 a_4922_4223.t2 GND 0.19205f
C236 a_4922_4223.t3 GND 0.07964f
C237 a_4922_4223.n0 GND 5.71483f
C238 a_4922_4223.n1 GND 4.4887f
C239 a_4922_4223.t0 GND 0.0575f
C240 rseg_2_v3_0.v5.t1 GND 0.03136f
C241 rseg_2_v3_0.v5.t2 GND 0.2006f
C242 rseg_2_v3_0.v5.t0 GND 0.19927f
C243 rseg_2_v3_0.v5.n0 GND 3.79324f
C244 rseg_2_v3_0.v36.t0 GND 0.01105f
C245 rseg_2_v3_0.v36.t2 GND 0.10186f
C246 rseg_2_v3_0.v36.t1 GND 0.09865f
C247 rseg_2_v3_0.v36.n0 GND 1.60945f
C248 rseg_2_v3_0.v7.t1 GND 0.01483f
C249 rseg_2_v3_0.v7.t2 GND 0.09877f
C250 rseg_2_v3_0.v7.t0 GND 0.09824f
C251 rseg_2_v3_0.v7.n0 GND 2.0341f
C252 rseg_2_v3_0.v10.t2 GND -0.04361f
C253 rseg_2_v3_0.v10.t0 GND -0.04348f
C254 rseg_2_v3_0.v10.n0 GND -0.75761f
C255 rseg_2_v3_0.v9.t1 GND 0.02389f
C256 rseg_2_v3_0.v9.t0 GND 0.20319f
C257 rseg_2_v3_0.v9.t2 GND 0.20254f
C258 rseg_2_v3_0.v9.n0 GND 3.55912f
C259 rseg_2_v3_0.v39.t1 GND 0.01071f
C260 rseg_2_v3_0.v39.t2 GND 0.10286f
C261 rseg_2_v3_0.v39.t0 GND 0.10091f
C262 rseg_2_v3_0.v39.n0 GND 1.7744f
C263 a_6728_6264.t4 GND 0.07551f
C264 a_6728_6264.t5 GND 0.0628f
C265 a_6728_6264.n0 GND 2.55379f
C266 a_6728_6264.t2 GND 0.0628f
C267 a_6728_6264.n1 GND 1.51601f
C268 a_6728_6264.t3 GND 0.0628f
C269 a_6728_6264.n2 GND 1.70138f
C270 a_6728_6264.t1 GND 0.06237f
C271 a_6728_6264.n3 GND 1.93846f
C272 a_6728_6264.t0 GND 0.06407f
C273 a_1610_4223.t1 GND 0.16728f
C274 a_1610_4223.t2 GND 0.17057f
C275 a_1610_4223.t3 GND 0.06972f
C276 a_1610_4223.n0 GND 4.89637f
C277 a_1610_4223.n1 GND 5.40937f
C278 a_1610_4223.t0 GND 0.0867f
C279 rseg_2_v3_0.v38.t2 GND 0.0214f
C280 rseg_2_v3_0.v38.t1 GND 0.19912f
C281 rseg_2_v3_0.v38.t0 GND 0.2041f
C282 rseg_2_v3_0.v38.n0 GND 3.48146f
C283 rseg_2_v3_0.v3.t2 GND 0.03192f
C284 rseg_2_v3_0.v3.t1 GND 0.19632f
C285 rseg_2_v3_0.v3.t0 GND 0.19438f
C286 rseg_2_v3_0.v3.n0 GND 3.27725f
C287 rseg_2_v3_0.v26.t1 GND 0.08808f
C288 rseg_2_v3_0.v26.t2 GND 0.09887f
C289 rseg_2_v3_0.v26.n0 GND 1.62687f
C290 rseg_2_v3_0.v25.t0 GND 0.02324f
C291 rseg_2_v3_0.v25.t2 GND 0.21195f
C292 rseg_2_v3_0.v25.t1 GND 0.23823f
C293 rseg_2_v3_0.v25.n0 GND 3.95638f
C294 a_1334_4223.t1 GND 0.16517f
C295 a_1334_4223.t3 GND 0.06747f
C296 a_1334_4223.n0 GND 5.15358f
C297 a_1334_4223.t2 GND 0.07601f
C298 a_1334_4223.n1 GND 4.60987f
C299 a_1334_4223.t0 GND 0.12791f
C300 rseg_2_v3_0.v37.t1 GND 0.01183f
C301 rseg_2_v3_0.v37.t2 GND 0.10716f
C302 rseg_2_v3_0.v37.t0 GND 0.11076f
C303 rseg_2_v3_0.v37.n0 GND 1.75654f
C304 rseg_2_v3_0.v44.t0 GND 0.0119f
C305 rseg_2_v3_0.v44.t2 GND 0.10582f
C306 rseg_2_v3_0.v44.t1 GND 0.10271f
C307 rseg_2_v3_0.v44.n0 GND 1.75822f
C308 a_5900_6264.t3 GND 0.03955f
C309 a_5900_6264.t1 GND 0.03423f
C310 a_5900_6264.n0 GND 1.24539f
C311 a_5900_6264.t2 GND 0.04042f
C312 a_5900_6264.t4 GND 0.03423f
C313 a_5900_6264.n1 GND 1.28824f
C314 a_5900_6264.n2 GND 0.78371f
C315 a_5900_6264.t0 GND 0.03423f
C316 a_5198_4223.t2 GND 0.16998f
C317 a_5198_4223.t4 GND 0.07011f
C318 a_5198_4223.n0 GND 4.88166f
C319 a_5198_4223.t1 GND 0.05584f
C320 a_5198_4223.n1 GND 0.59217f
C321 a_5198_4223.t3 GND 0.15734f
C322 a_5198_4223.n2 GND 4.21706f
C323 a_5198_4223.t0 GND 0.05584f
C324 a_7004_6264.t4 GND 0.04844f
C325 a_7004_6264.t2 GND 0.03452f
C326 a_7004_6264.n0 GND 1.72763f
C327 a_7004_6264.t1 GND 0.03452f
C328 a_7004_6264.n1 GND 0.84517f
C329 a_7004_6264.t3 GND 0.04172f
C330 a_7004_6264.n2 GND 1.43346f
C331 a_7004_6264.t0 GND 0.03452f
C332 a_2714_4223.t1 GND 0.1514f
C333 a_2714_4223.t3 GND 0.06185f
C334 a_2714_4223.n0 GND 4.46413f
C335 a_2714_4223.t4 GND 0.07321f
C336 a_2714_4223.n1 GND 1.20642f
C337 a_2714_4223.t2 GND 0.12979f
C338 a_2714_4223.n2 GND 4.33997f
C339 a_2714_4223.t0 GND 0.07321f
C340 rseg_2_v3_0.v40.t1 GND 0.02546f
C341 rseg_2_v3_0.v40.t2 GND 0.16114f
C342 rseg_2_v3_0.v40.n0 GND 4.57606f
C343 rseg_2_v3_0.v40.t0 GND 0.63734f
C344 a_1886_4223.t1 GND 0.17697f
C345 a_1886_4223.t3 GND 0.07252f
C346 a_1886_4223.n0 GND 5.33538f
C347 a_1886_4223.t2 GND 0.15093f
C348 a_1886_4223.n1 GND 5.6647f
C349 a_1886_4223.t0 GND 0.0995f
C350 rseg_2_v3_0.v1.t1 GND 0.01856f
C351 rseg_2_v3_0.v1.t2 GND 0.11517f
C352 rseg_2_v3_0.v1.n0 GND 1.95957f
C353 rseg_2_v3_0.v1.t0 GND 0.1067f
C354 rseg_2_v3_0.v27.t1 GND 0.01112f
C355 rseg_2_v3_0.v27.t2 GND 0.10492f
C356 rseg_2_v3_0.v27.t0 GND 0.10143f
C357 rseg_2_v3_0.v27.n0 GND 1.69051f
C358 rseg_2_v3_0.v22.t1 GND 0.01149f
C359 rseg_2_v3_0.v22.t0 GND 0.09509f
C360 rseg_2_v3_0.v22.t2 GND 0.09501f
C361 rseg_2_v3_0.v22.n0 GND 1.75955f
C362 rseg_2_v3_0.v41.t1 GND 0.02297f
C363 rseg_2_v3_0.v41.t2 GND 0.20624f
C364 rseg_2_v3_0.v41.t0 GND 0.22762f
C365 rseg_2_v3_0.v41.n0 GND 4.16348f
C366 a_2162_4223.t1 GND 0.06748f
C367 a_2162_4223.t3 GND 0.053f
C368 a_2162_4223.n0 GND 2.83277f
C369 a_2162_4223.t2 GND 0.03679f
C370 a_2162_4223.n1 GND 2.82036f
C371 a_2162_4223.t0 GND 0.08959f
C372 rseg_2_v3_0.v24.t0 GND 0.01594f
C373 rseg_2_v3_0.v24.t1 GND 0.16274f
C374 rseg_2_v3_0.v24.t2 GND 0.59169f
C375 rseg_2_v3_0.v24.n0 GND 3.93737f
C376 a_4094_4223.t1 GND 0.14562f
C377 a_4094_4223.t2 GND 0.18645f
C378 a_4094_4223.t3 GND 0.0771f
C379 a_4094_4223.n0 GND 5.74363f
C380 a_4094_4223.n1 GND 4.28874f
C381 a_4094_4223.t0 GND 0.05846f
C382 a_2990_4223.t1 GND 0.15567f
C383 a_2990_4223.t3 GND 0.07037f
C384 a_2990_4223.n0 GND 4.70467f
C385 a_2990_4223.t2 GND 0.06564f
C386 a_2990_4223.n1 GND 4.64301f
C387 a_2990_4223.t0 GND 0.16064f
C388 rseg_2_v3_0.v6.t1 GND 0.01011f
C389 rseg_2_v3_0.v6.t0 GND 0.08506f
C390 rseg_2_v3_0.v6.t2 GND 0.08454f
C391 rseg_2_v3_0.v6.n0 GND 1.70684f
C392 a_6176_6264.t4 GND 0.06307f
C393 a_6176_6264.t3 GND 0.07374f
C394 a_6176_6264.t5 GND 0.06204f
C395 a_6176_6264.n0 GND 2.40254f
C396 a_6176_6264.t2 GND 0.06204f
C397 a_6176_6264.n1 GND 1.44859f
C398 a_6176_6264.t1 GND 0.06204f
C399 a_6176_6264.n2 GND 1.42112f
C400 a_6176_6264.n3 GND 1.54318f
C401 a_6176_6264.t0 GND 0.06164f
C402 a_3542_4223.t1 GND 0.17175f
C403 a_3542_4223.t2 GND 0.1868f
C404 a_3542_4223.t3 GND 0.07658f
C405 a_3542_4223.n0 GND 5.49565f
C406 a_3542_4223.n1 GND 4.99847f
C407 a_3542_4223.t0 GND 0.07075f
C408 a_4646_4223.t1 GND 0.08612f
C409 a_4646_4223.t2 GND 0.11548f
C410 a_4646_4223.t3 GND 0.04818f
C411 a_4646_4223.n0 GND 3.58176f
C412 a_4646_4223.n1 GND 2.4369f
C413 a_4646_4223.t0 GND 0.03156f
C414 a_3266_4223.t2 GND 0.15559f
C415 a_3266_4223.t1 GND 0.06731f
C416 a_3266_4223.n0 GND 4.60037f
C417 a_3266_4223.t3 GND 0.16937f
C418 a_3266_4223.t4 GND 0.06934f
C419 a_3266_4223.n1 GND 4.88352f
C420 a_3266_4223.n2 GND 0.88718f
C421 a_3266_4223.t0 GND 0.06731f
C422 rseg_2_v3_0.v8.t0 GND 0.01313f
C423 rseg_2_v3_0.v8.t2 GND 0.15978f
C424 rseg_2_v3_0.v8.t1 GND 0.5213f
C425 rseg_2_v3_0.v8.n0 GND 3.70736f
C426 a_3818_4223.t1 GND 0.14851f
C427 a_3818_4223.t2 GND 0.17024f
C428 a_3818_4223.t3 GND 0.07006f
C429 a_3818_4223.n0 GND 5.08543f
C430 a_3818_4223.n1 GND 4.26715f
C431 a_3818_4223.t0 GND 0.05862f
C432 rseg_2_v3_0.v43.t0 GND 0.01122f
C433 rseg_2_v3_0.v43.t1 GND 0.10468f
C434 rseg_2_v3_0.v43.t2 GND 0.1019f
C435 rseg_2_v3_0.v43.n0 GND 1.77793f
C436 a_2438_4223.t1 GND 0.13926f
C437 a_2438_4223.t3 GND 0.0925f
C438 a_2438_4223.n0 GND 5.29359f
C439 a_2438_4223.t2 GND 0.07081f
C440 a_2438_4223.n1 GND 5.33076f
C441 a_2438_4223.t0 GND 0.17307f
C442 a_6452_6264.t1 GND 0.06308f
C443 a_6452_6264.t3 GND 0.0615f
C444 a_6452_6264.n0 GND 1.73123f
C445 a_6452_6264.t2 GND 0.06193f
C446 a_6452_6264.n1 GND 1.55195f
C447 a_6452_6264.t4 GND 0.07406f
C448 a_6452_6264.t5 GND 0.06193f
C449 a_6452_6264.n2 GND 2.46074f
C450 a_6452_6264.n3 GND 1.47166f
C451 a_6452_6264.t0 GND 0.06193f
C452 a_5474_4223.t3 GND 0.16318f
C453 a_5474_4223.t2 GND 0.06702f
C454 a_5474_4223.n0 GND 5.04796f
C455 a_5474_4223.t1 GND 0.12781f
C456 a_5474_4223.n1 GND 4.03512f
C457 a_5474_4223.t0 GND 0.05892f
C458 a_4370_4223.t2 GND 0.21223f
C459 a_4370_4223.t1 GND 0.08827f
C460 a_4370_4223.n0 GND 6.60332f
C461 a_4370_4223.t3 GND 0.0607f
C462 a_4370_4223.n1 GND 4.57762f
C463 a_4370_4223.t0 GND 0.15786f
.ends

