* PEX produced on Mon Jun  9 18:31:02 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from top_segment_4.ext - technology: sky130A

.subckt top_segment_4_posim V0 V63 DEC0 DEC1 DEC2 DEC3 b0 b1 b2 b3 bb0 bb1 bb2 bb3 VOUT
+ GND VPB
X0 rseg_4_routing_0/rseg_4_v3_0.v39.t2 rseg_4_routing_0/rseg_4_v3_0.v40.t2 GND.t7 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X1 rseg_4_routing_0/rseg_4_v3_0.v1.t0 V0.t1 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X2 a_31783_n8174.t4 b3.t0 a_36412_n5474.t2 VPB.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X3 a_33081_n6738.t3 DEC1.t0 rseg_4_routing_0/rseg_4_v3_0.v30.t1 VPB.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X4 rseg_4_routing_0/rseg_4_v3_0.v57.t2 DEC3.t0 a_31543_n6738.t3 VPB.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X5 rseg_4_routing_0/rseg_4_v3_0.v61.t1 rseg_4_routing_0/rseg_4_v3_0.v60.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=2.14
X6 GND.t21 GND.t22 GND.t7 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X7 a_32529_n6738.t1 DEC3.t1 rseg_4_routing_0/rseg_4_v3_0.v60.t1 VPB.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X8 rseg_4_routing_0/rseg_4_v3_0.v47.t1 rseg_4_routing_0/rseg_4_v3_0.v48.t1 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X9 a_36846_n4393.t2 b1.t0 a_35686_n4393.t1 VPB.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X10 a_32805_n6738.t4 DEC1.t1 rseg_4_routing_0/rseg_4_v3_0.v29.t1 VPB.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X11 a_33081_n6738.t0 DEC2.t0 rseg_4_routing_0/rseg_4_v3_0.v46.t1 VPB.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X12 rseg_4_routing_0/rseg_4_v3_0.v51.t0 rseg_4_routing_0/rseg_4_v3_0.v52.t1 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X13 rseg_4_routing_0/rseg_4_v3_0.v41.t2 DEC2.t1 a_31543_n6738.t1 VPB.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X14 a_35584_n5474.t2 bb3.t0 a_32529_n6738.t3 VPB.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X15 rseg_4_routing_0/rseg_4_v3_0.v55.t2 rseg_4_routing_0/rseg_4_v3_0.v56.t2 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.63
X16 rseg_4_routing_0/rseg_4_v3_0.v43.t0 rseg_4_routing_0/rseg_4_v3_0.v42.t1 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X17 GND.t18 GND.t19 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X18 rseg_4_routing_0/rseg_4_v3_0.v37.t1 rseg_4_routing_0/rseg_4_v3_0.v36.t1 GND.t7 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X19 a_36412_n5474.t0 bb3.t1 a_33357_n6738.t3 VPB.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X20 a_33081_n6738.t4 DEC3.t2 rseg_4_routing_0/rseg_4_v3_0.v62.t1 VPB.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X21 rseg_4_routing_0/rseg_4_v3_0.v33.t0 DEC2.t2 a_29969_n8174.t4 VPB.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X22 a_36266_n4393.t2 bb1.t0 a_35686_n4393.t0 VPB.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X23 rseg_4_routing_0/rseg_4_v3_0.v47.t2 rseg_4_routing_0/rseg_4_v3_0.v46.t2 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X24 rseg_4_routing_0/rseg_4_v3_0.v49.t1 rseg_4_routing_0/rseg_4_v3_0.v50.t1 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X25 a_30955_n8174.t4 DEC2.t3 rseg_4_routing_0/rseg_4_v3_0.v36.t2 VPB.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X26 rseg_4_routing_0/rseg_4_v3_0.v33.t1 rseg_4_routing_0/rseg_4_v3_0.v32.t2 GND.t7 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X27 GND.t5 GND.t6 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X28 a_35990_n4393.t0 bb2.t0 a_36412_n5474.t1 VPB.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X29 GND.t8 GND.t9 GND.t7 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X30 a_33357_n6738.t1 DEC3.t3 V63.t1 VPB.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X31 rseg_4_routing_0/rseg_4_v3_0.v3.t0 DEC0.t0 a_30521_n8174.t0 VPB.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X32 rseg_4_routing_0/rseg_4_v3_0.v17.t1 DEC1.t2 a_29969_n8174.t2 VPB.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X33 rseg_4_routing_0/rseg_4_v3_0.v27.t2 rseg_4_routing_0/rseg_4_v3_0.v26.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X34 rseg_4_routing_0/rseg_4_v3_0.v51.t2 rseg_4_routing_0/rseg_4_v3_0.v50.t2 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X35 GND.t25 GND.t26 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X36 rseg_4_routing_0/rseg_4_v3_0.v3.t1 rseg_4_routing_0/rseg_4_v3_0.v2.t1 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X37 a_31507_n8174.t4 DEC2.t4 rseg_4_routing_0/rseg_4_v3_0.v38.t2 VPB.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X38 rseg_4_routing_0/rseg_4_v3_0.v53.t1 rseg_4_routing_0/rseg_4_v3_0.v52.t0 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X39 rseg_4_routing_0/rseg_4_v3_0.v27.t0 rseg_4_routing_0/rseg_4_v3_0.v28.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X40 a_36846_n4393.t1 b2.t0 a_34638_n5474.t1 VPB.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X41 rseg_4_routing_0/rseg_4_v3_0.v51.t1 DEC3.t4 a_30521_n8174.t1 VPB.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X42 a_32529_n6738.t4 DEC0.t1 rseg_4_routing_0/rseg_4_v3_0.v12.t0 VPB.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X43 rseg_4_routing_0/rseg_4_v3_0.v18.t1 DEC1.t3 a_30245_n8174.t2 VPB.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X44 GND.t39 GND.t40 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.63
X45 rseg_4_routing_0/rseg_4_v3_0.v41.t1 rseg_4_routing_0/rseg_4_v3_0.v40.t1 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X46 rseg_4_routing_0/rseg_4_v3_0.v31.t1 rseg_4_routing_0/rseg_4_v3_0.v32.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X47 a_33357_n6738.t0 DEC0.t2 rseg_4_routing_0/rseg_4_v3_0.v15.t0 VPB.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X48 rseg_4_routing_0/rseg_4_v3_0.v10.t0 DEC0.t3 a_31819_n6738.t0 VPB.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X49 rseg_4_routing_0/rseg_4_v3_0.v55.t0 rseg_4_routing_0/rseg_4_v3_0.v54.t1 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X50 a_35686_n4393.t2 b0.t0 VOUT.t1 VPB.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X51 rseg_4_routing_0/rseg_4_v3_0.v39.t0 rseg_4_routing_0/rseg_4_v3_0.v38.t1 GND.t7 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X52 a_36266_n4393.t0 b2.t1 a_35190_n5474.t1 VPB.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X53 rseg_4_routing_0/rseg_4_v3_0.v45.t1 rseg_4_routing_0/rseg_4_v3_0.v46.t0 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X54 a_31231_n8174.t1 DEC3.t5 rseg_4_routing_0/rseg_4_v3_0.v53.t2 VPB.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X55 rseg_4_routing_0/rseg_4_v3_0.v49.t2 rseg_4_routing_0/rseg_4_v3_0.v48.t2 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X56 a_30955_n8174.t2 DEC1.t4 rseg_4_routing_0/rseg_4_v3_0.v20.t1 VPB.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X57 a_31783_n8174.t2 DEC1.t5 rseg_4_routing_0/rseg_4_v3_0.v23.t1 VPB.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X58 rseg_4_routing_0/rseg_4_v3_0.v42.t2 DEC2.t5 a_31819_n6738.t4 VPB.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X59 rseg_4_routing_0/rseg_4_v3_0.v25.t2 DEC1.t6 a_31543_n6738.t4 VPB.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X60 rseg_4_routing_0/rseg_4_v3_0.v53.t0 rseg_4_routing_0/rseg_4_v3_0.v54.t0 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X61 a_32529_n6738.t2 DEC1.t7 rseg_4_routing_0/rseg_4_v3_0.v28.t1 VPB.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X62 a_36570_n4393.t2 b1.t1 a_35382_n4393.t1 VPB.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X63 rseg_4_routing_0/rseg_4_v3_0.v29.t2 rseg_4_routing_0/rseg_4_v3_0.v28.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X64 a_32095_n6738.t3 bb3.t2 a_35466_n5474.t2 VPB.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X65 rseg_4_routing_0/rseg_4_v3_0.v58.t1 DEC3.t6 a_31819_n6738.t1 VPB.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X66 GND.t23 GND.t24 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X67 a_33357_n6738.t2 DEC1.t8 rseg_4_routing_0/rseg_4_v3_0.v31.t0 VPB.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X68 rseg_4_routing_0/rseg_4_v3_0.v15.t2 rseg_4_routing_0/rseg_4_v3_0.v14.t2 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X69 a_32529_n6738.t0 DEC2.t6 rseg_4_routing_0/rseg_4_v3_0.v44.t1 VPB.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X70 rseg_4_routing_0/rseg_4_v3_0.v57.t1 rseg_4_routing_0/rseg_4_v3_0.v58.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.78
X71 rseg_4_routing_0/rseg_4_v3_0.v49.t0 DEC3.t7 a_29969_n8174.t1 VPB.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X72 rseg_4_routing_0/rseg_4_v3_0.v26.t1 DEC1.t9 a_31819_n6738.t2 VPB.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X73 a_36570_n4393.t0 bb2.t1 a_35860_n5474.t0 VPB.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X74 a_32805_n6738.t3 DEC3.t8 rseg_4_routing_0/rseg_4_v3_0.v61.t0 VPB.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X75 rseg_4_routing_0/rseg_4_v3_0.v1.t1 DEC0.t4 a_29969_n8174.t0 VPB.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X76 rseg_4_routing_0/rseg_4_v3_0.v56.t1 DEC3.t9 a_31267_n6738.t1 VPB.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X77 rseg_4_routing_0/rseg_4_v3_0.v7.t1 rseg_4_routing_0/rseg_4_v3_0.v8.t1 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X78 a_33357_n6738.t4 DEC2.t7 rseg_4_routing_0/rseg_4_v3_0.v47.t0 VPB.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X79 V0.t0 DEC0.t5 a_29693_n8174.t0 VPB.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X80 rseg_4_routing_0/rseg_4_v3_0.v61.t2 rseg_4_routing_0/rseg_4_v3_0.v62.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=2.4
X81 a_35860_n5474.t2 bb3.t3 a_32805_n6738.t1 VPB.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X82 rseg_4_routing_0/rseg_4_v3_0.v37.t0 rseg_4_routing_0/rseg_4_v3_0.v38.t0 GND.t7 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X83 rseg_4_routing_0/rseg_4_v3_0.v33.t2 rseg_4_routing_0/rseg_4_v3_0.v34.t1 GND.t7 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X84 rseg_4_routing_0/rseg_4_v3_0.v35.t0 rseg_4_routing_0/rseg_4_v3_0.v36.t0 GND.t7 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X85 GND.t13 GND.t14 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X86 rseg_4_routing_0/rseg_4_v3_0.v23.t2 rseg_4_routing_0/rseg_4_v3_0.v24.t2 GND.t27 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X87 rseg_4_routing_0/rseg_4_v3_0.v50.t0 DEC3.t10 a_30245_n8174.t1 VPB.t87 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X88 rseg_4_routing_0/rseg_4_v3_0.v19.t1 rseg_4_routing_0/rseg_4_v3_0.v18.t0 GND.t32 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X89 rseg_4_routing_0/rseg_4_v3_0.v34.t0 DEC2.t8 a_30245_n8174.t4 VPB.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X90 rseg_4_routing_0/rseg_4_v3_0.v11.t2 rseg_4_routing_0/rseg_4_v3_0.v10.t2 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X91 rseg_4_routing_0/rseg_4_v3_0.v29.t0 rseg_4_routing_0/rseg_4_v3_0.v30.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X92 rseg_4_routing_0/rseg_4_v3_0.v13.t2 rseg_4_routing_0/rseg_4_v3_0.v12.t1 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X93 a_34638_n5474.t0 b3.t1 a_29693_n8174.t3 VPB.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X94 a_31507_n8174.t0 DEC0.t6 rseg_4_routing_0/rseg_4_v3_0.v6.t0 VPB.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X95 a_31231_n8174.t4 DEC2.t9 rseg_4_routing_0/rseg_4_v3_0.v37.t2 VPB.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X96 rseg_4_routing_0/rseg_4_v3_0.v32.t1 DEC2.t10 a_29693_n8174.t4 VPB.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X97 rseg_4_routing_0/rseg_4_v3_0.v8.t0 DEC0.t7 a_31267_n6738.t0 VPB.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X98 rseg_4_routing_0/rseg_4_v3_0.v9.t1 rseg_4_routing_0/rseg_4_v3_0.v10.t1 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X99 a_35466_n5474.t0 b3.t2 a_30521_n8174.t3 VPB.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X100 rseg_4_routing_0/rseg_4_v3_0.v25.t1 rseg_4_routing_0/rseg_4_v3_0.v24.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X101 a_35990_n4393.t2 bb1.t1 a_35382_n4393.t2 VPB.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X102 rseg_4_routing_0/rseg_4_v3_0.v11.t1 rseg_4_routing_0/rseg_4_v3_0.v12.t2 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X103 rseg_4_routing_0/rseg_4_v3_0.v11.t0 DEC0.t8 a_32095_n6738.t0 VPB.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X104 V63.t0 rseg_4_routing_0/rseg_4_v3_0.v62.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X105 a_30955_n8174.t0 DEC0.t9 rseg_4_routing_0/rseg_4_v3_0.v4.t0 VPB.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X106 a_31507_n8174.t3 b3.t3 a_36136_n5474.t1 VPB.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X107 rseg_4_routing_0/rseg_4_v3_0.v5.t2 rseg_4_routing_0/rseg_4_v3_0.v6.t1 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X108 rseg_4_routing_0/rseg_4_v3_0.v15.t1 rseg_4_routing_0/rseg_4_v3_0.v16.t0 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X109 a_31543_n6738.t0 bb3.t4 a_34914_n5474.t2 VPB.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X110 a_31231_n8174.t2 DEC1.t10 rseg_4_routing_0/rseg_4_v3_0.v21.t1 VPB.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X111 rseg_4_routing_0/rseg_4_v3_0.v3.t2 rseg_4_routing_0/rseg_4_v3_0.v4.t2 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X112 a_31783_n8174.t3 DEC2.t11 rseg_4_routing_0/rseg_4_v3_0.v39.t1 VPB.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X113 a_35990_n4393.t1 b2.t2 a_35466_n5474.t1 VPB.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X114 a_31783_n8174.t0 DEC0.t10 rseg_4_routing_0/rseg_4_v3_0.v7.t0 VPB.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X115 GND.t37 GND.t38 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X116 GND.t33 GND.t34 GND.t27 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X117 a_31507_n8174.t1 DEC3.t11 rseg_4_routing_0/rseg_4_v3_0.v54.t2 VPB.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X118 rseg_4_routing_0/rseg_4_v3_0.v16.t2 DEC1.t11 a_29693_n8174.t2 VPB.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X119 a_31231_n8174.t3 b3.t4 a_35860_n5474.t1 VPB.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X120 GND.t1 GND.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X121 a_32805_n6738.t2 DEC0.t11 rseg_4_routing_0/rseg_4_v3_0.v13.t0 VPB.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X122 rseg_4_routing_0/rseg_4_v3_0.v19.t2 DEC1.t12 a_30521_n8174.t2 VPB.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X123 GND.t35 GND.t36 GND.t27 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X124 rseg_4_routing_0/rseg_4_v3_0.v41.t0 rseg_4_routing_0/rseg_4_v3_0.v42.t0 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X125 a_31819_n6738.t3 bb3.t5 a_35190_n5474.t2 VPB.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X126 a_33081_n6738.t2 DEC0.t12 rseg_4_routing_0/rseg_4_v3_0.v14.t0 VPB.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X127 rseg_4_routing_0/rseg_4_v3_0.v21.t2 rseg_4_routing_0/rseg_4_v3_0.v20.t2 GND.t27 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X128 a_32805_n6738.t0 DEC2.t12 rseg_4_routing_0/rseg_4_v3_0.v45.t2 VPB.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X129 rseg_4_routing_0/rseg_4_v3_0.v59.t1 DEC3.t12 a_32095_n6738.t1 VPB.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X130 GND.t30 GND.t31 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X131 rseg_4_routing_0/rseg_4_v3_0.v17.t0 rseg_4_routing_0/rseg_4_v3_0.v16.t1 GND.t27 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X132 rseg_4_routing_0/rseg_4_v3_0.v40.t0 DEC2.t13 a_31267_n6738.t4 VPB.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X133 rseg_4_routing_0/rseg_4_v3_0.v59.t0 rseg_4_routing_0/rseg_4_v3_0.v60.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=2.04
X134 a_35382_n4393.t0 bb0.t0 VOUT.t0 VPB.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X135 GND.t10 GND.t11 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X136 rseg_4_routing_0/rseg_4_v3_0.v43.t1 DEC2.t14 a_32095_n6738.t4 VPB.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X137 rseg_4_routing_0/rseg_4_v3_0.v48.t0 DEC3.t13 a_29693_n8174.t1 VPB.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X138 a_36846_n4393.t0 bb2.t2 a_35584_n5474.t0 VPB.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X139 rseg_4_routing_0/rseg_4_v3_0.v43.t2 rseg_4_routing_0/rseg_4_v3_0.v44.t2 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X140 a_36136_n5474.t2 bb3.t6 a_33081_n6738.t1 VPB.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X141 rseg_4_routing_0/rseg_4_v3_0.v57.t0 rseg_4_routing_0/rseg_4_v3_0.v56.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X142 rseg_4_routing_0/rseg_4_v3_0.v17.t2 rseg_4_routing_0/rseg_4_v3_0.v18.t2 GND.t27 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X143 rseg_4_routing_0/rseg_4_v3_0.v59.t2 rseg_4_routing_0/rseg_4_v3_0.v58.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.94
X144 rseg_4_routing_0/rseg_4_v3_0.v1.t2 rseg_4_routing_0/rseg_4_v3_0.v2.t2 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X145 rseg_4_routing_0/rseg_4_v3_0.v31.t2 rseg_4_routing_0/rseg_4_v3_0.v30.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X146 rseg_4_routing_0/rseg_4_v3_0.v35.t2 rseg_4_routing_0/rseg_4_v3_0.v34.t2 GND.t7 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X147 a_36266_n4393.t1 bb2.t3 a_36136_n5474.t0 VPB.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X148 rseg_4_routing_0/rseg_4_v3_0.v2.t0 DEC0.t13 a_30245_n8174.t0 VPB.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X149 rseg_4_routing_0/rseg_4_v3_0.v7.t2 rseg_4_routing_0/rseg_4_v3_0.v6.t2 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X150 rseg_4_routing_0/rseg_4_v3_0.v13.t1 rseg_4_routing_0/rseg_4_v3_0.v14.t1 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X151 a_36570_n4393.t1 b2.t3 a_34914_n5474.t1 VPB.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X152 a_31231_n8174.t0 DEC0.t14 rseg_4_routing_0/rseg_4_v3_0.v5.t0 VPB.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X153 rseg_4_routing_0/rseg_4_v3_0.v21.t0 rseg_4_routing_0/rseg_4_v3_0.v22.t0 GND.t27 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X154 rseg_4_routing_0/rseg_4_v3_0.v5.t1 rseg_4_routing_0/rseg_4_v3_0.v4.t1 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X155 GND.t28 GND.t29 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X156 a_30955_n8174.t1 DEC3.t14 rseg_4_routing_0/rseg_4_v3_0.v52.t2 VPB.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X157 rseg_4_routing_0/rseg_4_v3_0.v19.t0 rseg_4_routing_0/rseg_4_v3_0.v20.t0 GND.t27 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X158 a_35190_n5474.t0 b3.t5 a_30245_n8174.t3 VPB.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X159 rseg_4_routing_0/rseg_4_v3_0.v9.t2 rseg_4_routing_0/rseg_4_v3_0.v8.t2 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X160 rseg_4_routing_0/rseg_4_v3_0.v23.t0 rseg_4_routing_0/rseg_4_v3_0.v22.t1 GND.t27 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X161 a_31783_n8174.t1 DEC3.t15 rseg_4_routing_0/rseg_4_v3_0.v55.t1 VPB.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X162 rseg_4_routing_0/rseg_4_v3_0.v35.t1 DEC2.t15 a_30521_n8174.t4 VPB.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X163 a_31507_n8174.t2 DEC1.t13 rseg_4_routing_0/rseg_4_v3_0.v22.t2 VPB.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X164 GND.t41 GND.t42 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X165 a_34914_n5474.t0 b3.t6 a_29969_n8174.t3 VPB.t71 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X166 a_31267_n6738.t3 bb3.t7 a_34638_n5474.t2 VPB.t86 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X167 rseg_4_routing_0/rseg_4_v3_0.v24.t1 DEC1.t14 a_31267_n6738.t2 VPB.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X168 rseg_4_routing_0/rseg_4_v3_0.v9.t0 DEC0.t15 a_31543_n6738.t2 VPB.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X169 GND.t16 GND.t17 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X170 rseg_4_routing_0/rseg_4_v3_0.v45.t0 rseg_4_routing_0/rseg_4_v3_0.v44.t0 GND.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X171 a_30955_n8174.t3 b3.t7 a_35584_n5474.t1 VPB.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X172 rseg_4_routing_0/rseg_4_v3_0.v27.t1 DEC1.t15 a_32095_n6738.t2 VPB.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X173 rseg_4_routing_0/rseg_4_v3_0.v25.t0 rseg_4_routing_0/rseg_4_v3_0.v26.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
R0 rseg_4_routing_0/rseg_4_v3_0.v39 rseg_4_routing_0/rseg_4_v3_0.v39.t1 674.658
R1 rseg_4_routing_0/rseg_4_v3_0.v39.n0 rseg_4_routing_0/rseg_4_v3_0.v39.t2 10.7653
R2 rseg_4_routing_0/rseg_4_v3_0.v39.n0 rseg_4_routing_0/rseg_4_v3_0.v39.t0 10.7376
R3 rseg_4_routing_0/rseg_4_v3_0.v39 rseg_4_routing_0/rseg_4_v3_0.v39.n0 4.0963
R4 rseg_4_routing_0/rseg_4_v3_0.v40 rseg_4_routing_0/rseg_4_v3_0.v40.t0 676.321
R5 rseg_4_routing_0/rseg_4_v3_0.v40.n0 rseg_4_routing_0/rseg_4_v3_0.v40.t1 13.4994
R6 rseg_4_routing_0/rseg_4_v3_0.v40.n0 rseg_4_routing_0/rseg_4_v3_0.v40.t2 10.7723
R7 rseg_4_routing_0/rseg_4_v3_0.v40 rseg_4_routing_0/rseg_4_v3_0.v40.n0 4.72836
R8 GND.n43 GND.n33 83508.7
R9 GND.n37 GND.n36 41345.1
R10 GND.n31 GND.n2 27409.3
R11 GND.n48 GND.n2 27409.3
R12 GND.n48 GND.n3 27406
R13 GND.n31 GND.n3 27406
R14 GND.n37 GND.n33 11233.5
R15 GND.n44 GND.n32 10335.8
R16 GND.n45 GND.n44 9944.8
R17 GND.n41 GND.n32 9286.94
R18 GND.n41 GND.n40 9174.63
R19 GND.n43 GND.n42 9053.82
R20 GND.n39 GND.n36 7714.56
R21 GND.n39 GND.n38 7518.99
R22 GND.n40 GND.n39 7478.84
R23 GND.n38 GND.n34 5608.79
R24 GND.n38 GND.n37 5016.48
R25 GND.n42 GND.n34 4715.04
R26 GND.n46 GND.n32 4451.25
R27 GND.n42 GND.n41 3889.56
R28 GND.n40 GND.n35 3752.03
R29 GND.n34 GND.n33 3562.79
R30 GND.n44 GND.n43 3153.67
R31 GND.t0 GND.t3 2122.95
R32 GND.t3 GND.t15 1868.79
R33 GND.n35 GND.t7 1788.29
R34 GND.n46 GND.t27 1746.89
R35 GND.t32 GND.t12 1737.69
R36 GND.n45 GND.t20 1727.34
R37 GND.n47 GND.t4 1239.73
R38 GND.t20 GND.n3 996.568
R39 GND.n36 GND.n2 966.668
R40 GND.n47 GND.t7 540.513
R41 GND.n14 GND.n13 475.536
R42 GND.n22 GND.n0 459.964
R43 GND.n13 GND.n12 458.043
R44 GND.n58 GND.n0 361.601
R45 GND.n36 GND.t0 242.656
R46 GND.n16 GND.n15 180.087
R47 GND.n52 GND.n51 171.339
R48 GND.n28 GND.n27 171.339
R49 GND.n20 GND.n19 171.126
R50 GND.n56 GND.n55 170.274
R51 GND.n7 GND.n6 170.274
R52 GND.n11 GND.n10 170.274
R53 GND.n24 GND.n23 170.06
R54 GND.n54 GND.n53 151.5
R55 GND.n9 GND.n8 151.5
R56 GND.n26 GND.n25 151.5
R57 GND.n18 GND.n17 148.087
R58 GND.n50 GND.n49 137.47
R59 GND.n12 GND.n11 137.419
R60 GND.n30 GND.n29 136.435
R61 GND.t15 GND.n35 134.554
R62 GND.t4 GND.n46 117.303
R63 GND.n15 GND.n14 102.433
R64 GND.n58 GND.n57 99.6436
R65 GND.n17 GND.n16 98.1667
R66 GND.t12 GND.n45 95.4527
R67 GND.n10 GND.n9 82.8067
R68 GND.n8 GND.n7 80.6733
R69 GND.n19 GND.n18 72.14
R70 GND.n21 GND.n20 72.14
R71 GND.n6 GND.n1 65.3133
R72 GND.n51 GND.n50 63.18
R73 GND.n29 GND.n28 61.0467
R74 GND.n27 GND.n26 61.0467
R75 GND.n53 GND.n52 58.9133
R76 GND.n55 GND.n54 56.78
R77 GND.n25 GND.n24 54.6467
R78 GND.n23 GND.n22 54.6467
R79 GND.n57 GND.n56 52.0867
R80 GND.n5 GND.t11 44.7381
R81 GND.n4 GND.t10 44.7381
R82 GND.n57 GND.t29 39.3159
R83 GND.n56 GND.t28 39.3159
R84 GND.n55 GND.t14 39.3159
R85 GND.n54 GND.t13 39.3159
R86 GND.n53 GND.t34 39.3159
R87 GND.n52 GND.t33 39.3159
R88 GND.n51 GND.t6 39.3159
R89 GND.n50 GND.t5 39.3159
R90 GND.n1 GND.t22 39.3159
R91 GND.n6 GND.t21 39.3159
R92 GND.n7 GND.t42 39.3159
R93 GND.n8 GND.t41 39.3159
R94 GND.n9 GND.t26 39.3159
R95 GND.n10 GND.t25 39.3159
R96 GND.n14 GND.t16 39.3159
R97 GND.n15 GND.t17 39.3159
R98 GND.n16 GND.t39 39.3159
R99 GND.n17 GND.t40 39.3159
R100 GND.n18 GND.t23 39.3159
R101 GND.n19 GND.t24 39.3159
R102 GND.n20 GND.t8 39.3159
R103 GND.n21 GND.t9 39.3159
R104 GND.n29 GND.t30 39.3159
R105 GND.n28 GND.t31 39.3159
R106 GND.n27 GND.t35 39.3159
R107 GND.n26 GND.t36 39.3159
R108 GND.n25 GND.t18 39.3159
R109 GND.n24 GND.t19 39.3159
R110 GND.n23 GND.t37 39.3159
R111 GND.n22 GND.t38 39.3159
R112 GND.n5 GND.t2 35.1381
R113 GND.n4 GND.t1 35.1381
R114 GND.n49 GND.n1 15.0979
R115 GND.n30 GND.n21 13.7851
R116 GND.n13 GND.n2 13.296
R117 GND.n3 GND.n0 13.296
R118 GND GND.n58 6.4005
R119 GND.n11 GND.n5 4.17828
R120 GND.n12 GND.n4 4.17828
R121 GND.n49 GND.n48 3.09574
R122 GND.n48 GND.n47 3.09574
R123 GND.n31 GND.n30 3.09574
R124 GND.n47 GND.n31 3.09574
R125 GND.t27 GND.t32 2.30055
R126 rseg_4_routing_0/rseg_4_v3_0.v1.n0 rseg_4_routing_0/rseg_4_v3_0.v1.t1 663.232
R127 rseg_4_routing_0/rseg_4_v3_0.v1.n0 rseg_4_routing_0/rseg_4_v3_0.v1.t2 10.6701
R128 rseg_4_routing_0/rseg_4_v3_0.v1.t0 rseg_4_routing_0/rseg_4_v3_0.v1.n0 10.5739
R129 V0.n0 V0.t0 668.13
R130 V0.n0 V0.t1 12.1073
R131 V0 V0.n0 0.274355
R132 b3.n0 b3.t1 217.555
R133 b3.n0 b3.t6 216.893
R134 b3.n1 b3.t5 216.893
R135 b3.n2 b3.t2 216.893
R136 b3.n3 b3.t7 216.893
R137 b3.n4 b3.t4 216.893
R138 b3.n5 b3.t3 216.893
R139 b3.n6 b3.t0 216.893
R140 b3.n6 b3.n5 0.663962
R141 b3.n5 b3.n4 0.663962
R142 b3.n4 b3.n3 0.663962
R143 b3.n3 b3.n2 0.663962
R144 b3.n2 b3.n1 0.663962
R145 b3.n1 b3.n0 0.663962
R146 b3 b3.n6 0.226462
R147 a_36412_n5474.n0 a_36412_n5474.t2 671.928
R148 a_36412_n5474.t0 a_36412_n5474.n0 671.475
R149 a_36412_n5474.n0 a_36412_n5474.t1 665.158
R150 a_31783_n8174.n0 a_31783_n8174.t1 673.378
R151 a_31783_n8174.t0 a_31783_n8174.n2 673.005
R152 a_31783_n8174.n1 a_31783_n8174.t4 669.523
R153 a_31783_n8174.n2 a_31783_n8174.t2 666.583
R154 a_31783_n8174.n0 a_31783_n8174.t3 666.583
R155 a_31783_n8174.n2 a_31783_n8174.n1 4.60675
R156 a_31783_n8174.n1 a_31783_n8174.n0 1.95467
R157 VPB.n93 VPB.n89 4436.17
R158 VPB.n93 VPB.n90 4436.17
R159 VPB.n95 VPB.n89 4436.17
R160 VPB.n95 VPB.n90 4436.17
R161 VPB.n101 VPB.n30 2671.14
R162 VPB.n101 VPB.n31 2671.14
R163 VPB.n103 VPB.n30 2671.14
R164 VPB.n103 VPB.n31 2671.14
R165 VPB.n82 VPB.n35 2671.14
R166 VPB.n84 VPB.n35 2671.14
R167 VPB.n84 VPB.n36 2671.14
R168 VPB.n82 VPB.n36 2671.14
R169 VPB.n125 VPB.n13 2671.14
R170 VPB.n125 VPB.n14 2671.14
R171 VPB.n127 VPB.n14 2671.14
R172 VPB.n127 VPB.n13 2671.14
R173 VPB.n117 VPB.n16 2671.14
R174 VPB.n119 VPB.n16 2671.14
R175 VPB.n119 VPB.n17 2671.14
R176 VPB.n117 VPB.n17 2671.14
R177 VPB.n109 VPB.n24 2671.14
R178 VPB.n109 VPB.n25 2671.14
R179 VPB.n111 VPB.n25 2671.14
R180 VPB.n111 VPB.n24 2671.14
R181 VPB.n71 VPB.n67 2671.14
R182 VPB.n73 VPB.n67 2671.14
R183 VPB.n73 VPB.n68 2671.14
R184 VPB.n71 VPB.n68 2671.14
R185 VPB.n63 VPB.n40 2671.14
R186 VPB.n63 VPB.n41 2671.14
R187 VPB.n61 VPB.n40 2671.14
R188 VPB.n61 VPB.n41 2671.14
R189 VPB.n54 VPB.n47 2671.14
R190 VPB.n54 VPB.n52 2671.14
R191 VPB.n56 VPB.n47 2671.14
R192 VPB.n56 VPB.n52 2671.14
R193 VPB.n133 VPB.n8 2671.14
R194 VPB.n133 VPB.n9 2671.14
R195 VPB.n135 VPB.n8 2671.14
R196 VPB.n135 VPB.n9 2671.14
R197 VPB.n142 VPB.n3 2671.14
R198 VPB.n142 VPB.n4 2671.14
R199 VPB.n140 VPB.n3 2671.14
R200 VPB.n140 VPB.n4 2671.14
R201 VPB.n86 VPB.n32 883.577
R202 VPB.n105 VPB.n28 883.577
R203 VPB.n92 VPB.n33 854.212
R204 VPB.n92 VPB.n91 854.212
R205 VPB.n96 VPB.n88 781.929
R206 VPB.n97 VPB.n96 781.929
R207 VPB.n81 VPB.n34 516.141
R208 VPB.n124 VPB.n123 516.141
R209 VPB.n70 VPB.n37 516.141
R210 VPB.n70 VPB.n69 516.141
R211 VPB.n143 VPB.n2 516.141
R212 VPB.n139 VPB.n2 516.141
R213 VPB.n60 VPB.n38 516.141
R214 VPB.t84 VPB.t23 475
R215 VPB.t54 VPB.t67 475
R216 VPB.t66 VPB.t8 475
R217 VPB.t28 VPB.t83 475
R218 VPB.t83 VPB.t24 475
R219 VPB.n100 VPB.n32 443.86
R220 VPB.n80 VPB.n79 443.86
R221 VPB.n79 VPB.n28 443.86
R222 VPB.n105 VPB.n104 443.86
R223 VPB.n104 VPB.n29 443.86
R224 VPB.n108 VPB.n107 443.86
R225 VPB.n19 VPB.n18 443.86
R226 VPB.n124 VPB.n122 443.86
R227 VPB.n69 VPB.n66 443.86
R228 VPB.n112 VPB.n23 443.86
R229 VPB.n113 VPB.n112 443.86
R230 VPB.n115 VPB.n114 443.86
R231 VPB.n114 VPB.n12 443.86
R232 VPB.n129 VPB.n128 443.86
R233 VPB.n128 VPB.n0 443.86
R234 VPB.n60 VPB.n59 443.86
R235 VPB.n58 VPB.n57 443.86
R236 VPB.n57 VPB.n46 443.86
R237 VPB.n136 VPB.n7 443.86
R238 VPB.n137 VPB.n136 443.86
R239 VPB.n139 VPB.n138 443.86
R240 VPB.t22 VPB.t53 431.25
R241 VPB.t82 VPB.t22 431.25
R242 VPB.t23 VPB.t82 431.25
R243 VPB.t10 VPB.t84 431.25
R244 VPB.t9 VPB.t10 431.25
R245 VPB.t67 VPB.t66 431.25
R246 VPB.t8 VPB.t28 431.25
R247 VPB.t74 VPB.t77 431.25
R248 VPB.t73 VPB.t74 431.25
R249 VPB.t70 VPB.t73 431.25
R250 VPB.t75 VPB.t72 431.25
R251 VPB.t72 VPB.t71 431.25
R252 VPB.t71 VPB.t76 431.25
R253 VPB.t33 VPB.t6 431.25
R254 VPB.t45 VPB.t33 431.25
R255 VPB.t79 VPB.t45 431.25
R256 VPB.t18 VPB.t60 431.25
R257 VPB.t1 VPB.t18 431.25
R258 VPB.t86 VPB.t1 431.25
R259 VPB.t52 VPB.t12 431.25
R260 VPB.t46 VPB.t52 431.25
R261 VPB.t81 VPB.t46 431.25
R262 VPB.t40 VPB.t48 431.25
R263 VPB.t48 VPB.t61 431.25
R264 VPB.t61 VPB.t11 431.25
R265 VPB.t85 VPB.t63 431.25
R266 VPB.t68 VPB.t85 431.25
R267 VPB.t29 VPB.t68 431.25
R268 VPB.t90 VPB.t41 431.25
R269 VPB.t56 VPB.t90 431.25
R270 VPB.t39 VPB.t56 431.25
R271 VPB.t0 VPB.t36 431.25
R272 VPB.t19 VPB.t0 431.25
R273 VPB.t50 VPB.t19 431.25
R274 VPB.t92 VPB.t37 431.25
R275 VPB.t37 VPB.t34 431.25
R276 VPB.t34 VPB.t16 431.25
R277 VPB.t88 VPB.t62 431.25
R278 VPB.t58 VPB.t88 431.25
R279 VPB.t44 VPB.t58 431.25
R280 VPB.t15 VPB.t64 431.25
R281 VPB.t59 VPB.t15 431.25
R282 VPB.t43 VPB.t59 431.25
R283 VPB.t31 VPB.t30 431.25
R284 VPB.t65 VPB.t31 431.25
R285 VPB.t57 VPB.t65 431.25
R286 VPB.t32 VPB.t87 431.25
R287 VPB.t87 VPB.t5 431.25
R288 VPB.t5 VPB.t14 431.25
R289 VPB.t93 VPB.t69 431.25
R290 VPB.t49 VPB.t93 431.25
R291 VPB.t17 VPB.t49 431.25
R292 VPB.t25 VPB.t26 431.25
R293 VPB.t26 VPB.t38 431.25
R294 VPB.t38 VPB.t20 431.25
R295 VPB.t89 VPB.t51 431.25
R296 VPB.t78 VPB.t89 431.25
R297 VPB.t42 VPB.t78 431.25
R298 VPB.t4 VPB.t13 431.25
R299 VPB.t13 VPB.t35 431.25
R300 VPB.t35 VPB.t2 431.25
R301 VPB.t91 VPB.t21 431.25
R302 VPB.t7 VPB.t91 431.25
R303 VPB.t47 VPB.t7 431.25
R304 VPB.t27 VPB.t80 431.25
R305 VPB.t80 VPB.t55 431.25
R306 VPB.t55 VPB.t3 431.25
R307 VPB.n18 VPB.n15 406.589
R308 VPB.t53 VPB.n89 379.062
R309 VPB.t24 VPB.n90 379.062
R310 VPB.t77 VPB.n30 379.062
R311 VPB.t76 VPB.n31 379.062
R312 VPB.t6 VPB.n82 379.062
R313 VPB.n84 VPB.t86 379.062
R314 VPB.t12 VPB.n13 379.062
R315 VPB.t11 VPB.n14 379.062
R316 VPB.t63 VPB.n117 379.062
R317 VPB.n119 VPB.t39 379.062
R318 VPB.t36 VPB.n24 379.062
R319 VPB.t16 VPB.n25 379.062
R320 VPB.t62 VPB.n71 379.062
R321 VPB.n73 VPB.t43 379.062
R322 VPB.t30 VPB.n40 379.062
R323 VPB.t14 VPB.n41 379.062
R324 VPB.t69 VPB.n47 379.062
R325 VPB.t20 VPB.n52 379.062
R326 VPB.t51 VPB.n8 379.062
R327 VPB.t2 VPB.n9 379.062
R328 VPB.t21 VPB.n3 379.062
R329 VPB.t3 VPB.n4 379.062
R330 VPB.n87 VPB.n34 371.2
R331 VPB.n77 VPB.n76 368.942
R332 VPB.n66 VPB.n23 368.942
R333 VPB.n99 VPB.n98 352.377
R334 VPB.n66 VPB.n65 343.341
R335 VPB.n39 VPB.n23 343.341
R336 VPB.n113 VPB.n21 343.341
R337 VPB.n115 VPB.n20 343.341
R338 VPB.n12 VPB.n10 343.341
R339 VPB.n131 VPB.n129 343.341
R340 VPB.n59 VPB.n58 339.954
R341 VPB.n44 VPB.n43 339.954
R342 VPB.n80 VPB.n78 332.8
R343 VPB.n28 VPB.n26 332.8
R344 VPB.n106 VPB.n105 332.8
R345 VPB.n29 VPB.n15 332.8
R346 VPB.n131 VPB.n130 320
R347 VPB.n65 VPB.n38 313.224
R348 VPB.n115 VPB.n113 310.966
R349 VPB.n50 VPB.n20 306.825
R350 VPB.n46 VPB.n7 297.788
R351 VPB.n50 VPB.n49 297.788
R352 VPB.n144 VPB.n1 295.154
R353 VPB.n122 VPB.n121 284.613
R354 VPB.n129 VPB.n12 284.613
R355 VPB.n49 VPB.n10 283.106
R356 VPB.n94 VPB.t9 281.25
R357 VPB.n76 VPB.n26 277.836
R358 VPB.n43 VPB.n39 277.836
R359 VPB.n107 VPB.n106 273.695
R360 VPB.n138 VPB.n137 272.565
R361 VPB.n130 VPB.n1 272.565
R362 VPB.n44 VPB.n21 269.93
R363 VPB.n78 VPB.n77 240.941
R364 VPB.n88 VPB.n87 236.8
R365 VPB.n99 VPB.n97 236.8
R366 VPB VPB.n144 225.882
R367 VPB.n102 VPB.t70 215.625
R368 VPB.n102 VPB.t75 215.625
R369 VPB.n83 VPB.t79 215.625
R370 VPB.t60 VPB.n83 215.625
R371 VPB.n126 VPB.t81 215.625
R372 VPB.n126 VPB.t40 215.625
R373 VPB.n118 VPB.t29 215.625
R374 VPB.t41 VPB.n118 215.625
R375 VPB.n110 VPB.t50 215.625
R376 VPB.n110 VPB.t92 215.625
R377 VPB.n72 VPB.t44 215.625
R378 VPB.t64 VPB.n72 215.625
R379 VPB.n62 VPB.t57 215.625
R380 VPB.n62 VPB.t32 215.625
R381 VPB.n55 VPB.t17 215.625
R382 VPB.n55 VPB.t25 215.625
R383 VPB.n134 VPB.t42 215.625
R384 VPB.n134 VPB.t4 215.625
R385 VPB.n141 VPB.t47 215.625
R386 VPB.n141 VPB.t27 215.625
R387 VPB.n78 VPB.n37 202.918
R388 VPB.n65 VPB.n64 202.918
R389 VPB.n53 VPB.n21 173.929
R390 VPB.n108 VPB.n26 166.024
R391 VPB.n64 VPB.n39 166.024
R392 VPB.n100 VPB.n99 163.766
R393 VPB.n132 VPB.n10 160.754
R394 VPB.n94 VPB.t54 150
R395 VPB.n144 VPB.n143 148.707
R396 VPB.n53 VPB.n20 137.036
R397 VPB.n132 VPB.n131 123.859
R398 VPB VPB.n0 117.46
R399 VPB.n87 VPB.n86 72.6593
R400 VPB.n97 VPB.n33 72.2828
R401 VPB.n91 VPB.n88 72.2828
R402 VPB.n98 VPB.n29 72.2828
R403 VPB.n86 VPB.n85 72.2828
R404 VPB.n85 VPB.n28 72.2828
R405 VPB.n81 VPB.n80 72.2828
R406 VPB.n32 VPB.n27 72.2828
R407 VPB.n105 VPB.n27 72.2828
R408 VPB.n123 VPB.n0 72.2828
R409 VPB.n122 VPB.n11 72.2828
R410 VPB.n129 VPB.n11 72.2828
R411 VPB.n116 VPB.n19 72.2828
R412 VPB.n116 VPB.n115 72.2828
R413 VPB.n107 VPB.n22 72.2828
R414 VPB.n113 VPB.n22 72.2828
R415 VPB.n76 VPB.n75 72.2828
R416 VPB.n75 VPB.n23 72.2828
R417 VPB.n77 VPB.n74 72.2828
R418 VPB.n74 VPB.n66 72.2828
R419 VPB.n121 VPB.n120 72.2828
R420 VPB.n120 VPB.n12 72.2828
R421 VPB.n43 VPB.n42 72.2828
R422 VPB.n59 VPB.n42 72.2828
R423 VPB.n45 VPB.n44 72.2828
R424 VPB.n58 VPB.n45 72.2828
R425 VPB.n51 VPB.n50 72.2828
R426 VPB.n51 VPB.n46 72.2828
R427 VPB.n49 VPB.n48 72.2828
R428 VPB.n48 VPB.n7 72.2828
R429 VPB.n130 VPB.n6 72.2828
R430 VPB.n137 VPB.n6 72.2828
R431 VPB.n5 VPB.n1 72.2828
R432 VPB.n138 VPB.n5 72.2828
R433 VPB.n90 VPB.n33 46.2505
R434 VPB.n91 VPB.n89 46.2505
R435 VPB.n98 VPB.n31 46.2505
R436 VPB.n85 VPB.n84 46.2505
R437 VPB.n82 VPB.n81 46.2505
R438 VPB.n30 VPB.n27 46.2505
R439 VPB.n123 VPB.n14 46.2505
R440 VPB.n13 VPB.n11 46.2505
R441 VPB.n117 VPB.n116 46.2505
R442 VPB.n25 VPB.n22 46.2505
R443 VPB.n75 VPB.n24 46.2505
R444 VPB.n74 VPB.n73 46.2505
R445 VPB.n71 VPB.n70 46.2505
R446 VPB.n120 VPB.n119 46.2505
R447 VPB.n42 VPB.n41 46.2505
R448 VPB.n47 VPB.n45 46.2505
R449 VPB.n52 VPB.n51 46.2505
R450 VPB.n48 VPB.n8 46.2505
R451 VPB.n9 VPB.n6 46.2505
R452 VPB.n5 VPB.n3 46.2505
R453 VPB.n4 VPB.n2 46.2505
R454 VPB.n40 VPB.n38 46.2505
R455 VPB.n106 VPB.n19 37.2711
R456 VPB.n121 VPB.n15 37.2711
R457 VPB.n35 VPB.n34 5.78175
R458 VPB.n83 VPB.n35 5.78175
R459 VPB.n101 VPB.n100 5.78175
R460 VPB.n102 VPB.n101 5.78175
R461 VPB.n79 VPB.n36 5.78175
R462 VPB.n83 VPB.n36 5.78175
R463 VPB.n104 VPB.n103 5.78175
R464 VPB.n103 VPB.n102 5.78175
R465 VPB.n67 VPB.n37 5.78175
R466 VPB.n72 VPB.n67 5.78175
R467 VPB.n109 VPB.n108 5.78175
R468 VPB.n110 VPB.n109 5.78175
R469 VPB.n18 VPB.n16 5.78175
R470 VPB.n118 VPB.n16 5.78175
R471 VPB.n125 VPB.n124 5.78175
R472 VPB.n126 VPB.n125 5.78175
R473 VPB.n69 VPB.n68 5.78175
R474 VPB.n72 VPB.n68 5.78175
R475 VPB.n112 VPB.n111 5.78175
R476 VPB.n111 VPB.n110 5.78175
R477 VPB.n114 VPB.n17 5.78175
R478 VPB.n118 VPB.n17 5.78175
R479 VPB.n128 VPB.n127 5.78175
R480 VPB.n127 VPB.n126 5.78175
R481 VPB.n61 VPB.n60 5.78175
R482 VPB.n62 VPB.n61 5.78175
R483 VPB.n57 VPB.n56 5.78175
R484 VPB.n56 VPB.n55 5.78175
R485 VPB.n136 VPB.n135 5.78175
R486 VPB.n135 VPB.n134 5.78175
R487 VPB.n140 VPB.n139 5.78175
R488 VPB.n141 VPB.n140 5.78175
R489 VPB.n64 VPB.n63 5.78175
R490 VPB.n63 VPB.n62 5.78175
R491 VPB.n54 VPB.n53 5.78175
R492 VPB.n55 VPB.n54 5.78175
R493 VPB.n133 VPB.n132 5.78175
R494 VPB.n134 VPB.n133 5.78175
R495 VPB.n143 VPB.n142 5.78175
R496 VPB.n142 VPB.n141 5.78175
R497 VPB.n93 VPB.n92 3.13609
R498 VPB.n94 VPB.n93 3.13609
R499 VPB.n96 VPB.n95 3.13609
R500 VPB.n95 VPB.n94 3.13609
R501 DEC1.n0 DEC1.t8 217.555
R502 DEC1.n7 DEC1.t11 217.555
R503 DEC1.n12 DEC1.t5 217.555
R504 DEC1.n5 DEC1.t6 216.893
R505 DEC1.n4 DEC1.t9 216.893
R506 DEC1.n3 DEC1.t15 216.893
R507 DEC1.n2 DEC1.t7 216.893
R508 DEC1.n1 DEC1.t1 216.893
R509 DEC1.n0 DEC1.t0 216.893
R510 DEC1.n7 DEC1.t2 216.893
R511 DEC1.n8 DEC1.t3 216.893
R512 DEC1.n9 DEC1.t12 216.893
R513 DEC1.n10 DEC1.t4 216.893
R514 DEC1.n11 DEC1.t10 216.893
R515 DEC1.n6 DEC1.t14 212.393
R516 DEC1.n13 DEC1.t13 212.393
R517 DEC1.n6 DEC1.n5 5.16396
R518 DEC1.n13 DEC1.n12 4.5005
R519 DEC1 DEC1.n13 1.88512
R520 DEC1 DEC1.n6 0.6755
R521 DEC1.n1 DEC1.n0 0.663962
R522 DEC1.n2 DEC1.n1 0.663962
R523 DEC1.n3 DEC1.n2 0.663962
R524 DEC1.n4 DEC1.n3 0.663962
R525 DEC1.n5 DEC1.n4 0.663962
R526 DEC1.n12 DEC1.n11 0.663962
R527 DEC1.n11 DEC1.n10 0.663962
R528 DEC1.n10 DEC1.n9 0.663962
R529 DEC1.n9 DEC1.n8 0.663962
R530 DEC1.n8 DEC1.n7 0.663962
R531 rseg_4_routing_0/rseg_4_v3_0.v30 rseg_4_routing_0/rseg_4_v3_0.v30.t1 675.843
R532 rseg_4_routing_0/rseg_4_v3_0.v30.n0 rseg_4_routing_0/rseg_4_v3_0.v30.t0 10.7393
R533 rseg_4_routing_0/rseg_4_v3_0.v30.n0 rseg_4_routing_0/rseg_4_v3_0.v30.t2 10.6478
R534 rseg_4_routing_0/rseg_4_v3_0.v30 rseg_4_routing_0/rseg_4_v3_0.v30.n0 0.682179
R535 a_33081_n6738.n1 a_33081_n6738.t2 672.764
R536 a_33081_n6738.n0 a_33081_n6738.t4 670.999
R537 a_33081_n6738.n0 a_33081_n6738.t1 666.655
R538 a_33081_n6738.n1 a_33081_n6738.t3 666.275
R539 a_33081_n6738.t0 a_33081_n6738.n2 666.275
R540 a_33081_n6738.n2 a_33081_n6738.n1 6.63383
R541 a_33081_n6738.n2 a_33081_n6738.n0 2.23175
R542 DEC3.n0 DEC3.t3 217.555
R543 DEC3.n10 DEC3.t13 217.555
R544 DEC3.n7 DEC3.t15 217.555
R545 DEC3.n6 DEC3.t9 216.893
R546 DEC3.n5 DEC3.t0 216.893
R547 DEC3.n4 DEC3.t6 216.893
R548 DEC3.n3 DEC3.t12 216.893
R549 DEC3.n2 DEC3.t1 216.893
R550 DEC3.n1 DEC3.t8 216.893
R551 DEC3.n0 DEC3.t2 216.893
R552 DEC3.n10 DEC3.t7 216.893
R553 DEC3.n11 DEC3.t10 216.893
R554 DEC3.n12 DEC3.t4 216.893
R555 DEC3.n9 DEC3.t14 216.893
R556 DEC3.n8 DEC3.t5 216.893
R557 DEC3.n7 DEC3.t11 216.893
R558 DEC3 DEC3.n6 6.64778
R559 DEC3 DEC3.n13 6.48592
R560 DEC3.n1 DEC3.n0 0.663962
R561 DEC3.n2 DEC3.n1 0.663962
R562 DEC3.n3 DEC3.n2 0.663962
R563 DEC3.n4 DEC3.n3 0.663962
R564 DEC3.n5 DEC3.n4 0.663962
R565 DEC3.n6 DEC3.n5 0.663962
R566 DEC3.n12 DEC3.n11 0.663962
R567 DEC3.n11 DEC3.n10 0.663962
R568 DEC3.n8 DEC3.n7 0.663962
R569 DEC3.n9 DEC3.n8 0.663962
R570 DEC3.n13 DEC3.n12 0.320692
R571 DEC3.n13 DEC3.n9 0.320692
R572 a_31543_n6738.n0 a_31543_n6738.t2 671.846
R573 a_31543_n6738.n2 a_31543_n6738.t3 667.794
R574 a_31543_n6738.t0 a_31543_n6738.n2 667.572
R575 a_31543_n6738.n0 a_31543_n6738.t4 665.36
R576 a_31543_n6738.n1 a_31543_n6738.t1 665.36
R577 a_31543_n6738.n1 a_31543_n6738.n0 6.63383
R578 a_31543_n6738.n2 a_31543_n6738.n1 4.51925
R579 rseg_4_routing_0/rseg_4_v3_0.v57 rseg_4_routing_0/rseg_4_v3_0.v57.t2 675.929
R580 rseg_4_routing_0/rseg_4_v3_0.v57.n0 rseg_4_routing_0/rseg_4_v3_0.v57.t0 10.7912
R581 rseg_4_routing_0/rseg_4_v3_0.v57.n0 rseg_4_routing_0/rseg_4_v3_0.v57.t1 10.6717
R582 rseg_4_routing_0/rseg_4_v3_0.v57 rseg_4_routing_0/rseg_4_v3_0.v57.n0 4.09783
R583 rseg_4_routing_0/rseg_4_v3_0.v61 rseg_4_routing_0/rseg_4_v3_0.v61.t0 675.904
R584 rseg_4_routing_0/rseg_4_v3_0.v61.n0 rseg_4_routing_0/rseg_4_v3_0.v61.t1 10.7652
R585 rseg_4_routing_0/rseg_4_v3_0.v61.n0 rseg_4_routing_0/rseg_4_v3_0.v61.t2 10.6927
R586 rseg_4_routing_0/rseg_4_v3_0.v61 rseg_4_routing_0/rseg_4_v3_0.v61.n0 1.36672
R587 rseg_4_routing_0/rseg_4_v3_0.v60 rseg_4_routing_0/rseg_4_v3_0.v60.t1 676.497
R588 rseg_4_routing_0/rseg_4_v3_0.v60.n0 rseg_4_routing_0/rseg_4_v3_0.v60.t0 10.7173
R589 rseg_4_routing_0/rseg_4_v3_0.v60.n0 rseg_4_routing_0/rseg_4_v3_0.v60.t2 10.675
R590 rseg_4_routing_0/rseg_4_v3_0.v60 rseg_4_routing_0/rseg_4_v3_0.v60.n0 2.06176
R591 a_32529_n6738.n1 a_32529_n6738.t4 672.396
R592 a_32529_n6738.n0 a_32529_n6738.t1 669.848
R593 a_32529_n6738.n0 a_32529_n6738.t3 666.222
R594 a_32529_n6738.n1 a_32529_n6738.t2 665.909
R595 a_32529_n6738.t0 a_32529_n6738.n2 665.909
R596 a_32529_n6738.n2 a_32529_n6738.n1 6.63383
R597 a_32529_n6738.n2 a_32529_n6738.n0 3.01508
R598 rseg_4_routing_0/rseg_4_v3_0.v47.t0 rseg_4_routing_0/rseg_4_v3_0.v47.n0 667.057
R599 rseg_4_routing_0/rseg_4_v3_0.v47.n0 rseg_4_routing_0/rseg_4_v3_0.v47.t2 10.6819
R600 rseg_4_routing_0/rseg_4_v3_0.v47.n0 rseg_4_routing_0/rseg_4_v3_0.v47.t1 10.5739
R601 rseg_4_routing_0/rseg_4_v3_0.v48.t0 rseg_4_routing_0/rseg_4_v3_0.v48.n0 668.13
R602 rseg_4_routing_0/rseg_4_v3_0.v48.n0 rseg_4_routing_0/rseg_4_v3_0.v48.t2 12.176
R603 rseg_4_routing_0/rseg_4_v3_0.v48.n0 rseg_4_routing_0/rseg_4_v3_0.v48.t1 12.0758
R604 b1.n0 b1.t0 217.555
R605 b1.n0 b1.t1 216.893
R606 b1 b1.n0 0.214442
R607 a_35686_n4393.n0 a_35686_n4393.t1 666.561
R608 a_35686_n4393.n0 a_35686_n4393.t2 666.096
R609 a_35686_n4393.t0 a_35686_n4393.n0 665.352
R610 a_36846_n4393.t0 a_36846_n4393.n0 667.659
R611 a_36846_n4393.n0 a_36846_n4393.t2 665.933
R612 a_36846_n4393.n0 a_36846_n4393.t1 665.299
R613 rseg_4_routing_0/rseg_4_v3_0.v29 rseg_4_routing_0/rseg_4_v3_0.v29.t1 675.904
R614 rseg_4_routing_0/rseg_4_v3_0.v29.n0 rseg_4_routing_0/rseg_4_v3_0.v29.t2 10.7799
R615 rseg_4_routing_0/rseg_4_v3_0.v29.n0 rseg_4_routing_0/rseg_4_v3_0.v29.t0 10.6965
R616 rseg_4_routing_0/rseg_4_v3_0.v29 rseg_4_routing_0/rseg_4_v3_0.v29.n0 1.35813
R617 a_32805_n6738.n1 a_32805_n6738.t2 672.581
R618 a_32805_n6738.n0 a_32805_n6738.t3 670.423
R619 a_32805_n6738.n0 a_32805_n6738.t1 666.391
R620 a_32805_n6738.n1 a_32805_n6738.t4 666.092
R621 a_32805_n6738.t0 a_32805_n6738.n2 666.092
R622 a_32805_n6738.n2 a_32805_n6738.n1 6.63383
R623 a_32805_n6738.n2 a_32805_n6738.n0 2.62342
R624 DEC2.n0 DEC2.t7 217.555
R625 DEC2.n7 DEC2.t10 217.555
R626 DEC2.n12 DEC2.t11 217.555
R627 DEC2.n5 DEC2.t1 216.893
R628 DEC2.n4 DEC2.t5 216.893
R629 DEC2.n3 DEC2.t14 216.893
R630 DEC2.n2 DEC2.t6 216.893
R631 DEC2.n1 DEC2.t12 216.893
R632 DEC2.n0 DEC2.t0 216.893
R633 DEC2.n7 DEC2.t2 216.893
R634 DEC2.n8 DEC2.t8 216.893
R635 DEC2.n9 DEC2.t15 216.893
R636 DEC2.n10 DEC2.t3 216.893
R637 DEC2.n11 DEC2.t9 216.893
R638 DEC2.n6 DEC2.t13 212.393
R639 DEC2.n13 DEC2.t4 212.393
R640 DEC2.n6 DEC2.n5 5.16396
R641 DEC2.n13 DEC2.n12 4.5005
R642 DEC2 DEC2.n13 1.89425
R643 DEC2.n1 DEC2.n0 0.663962
R644 DEC2.n2 DEC2.n1 0.663962
R645 DEC2.n3 DEC2.n2 0.663962
R646 DEC2.n4 DEC2.n3 0.663962
R647 DEC2.n5 DEC2.n4 0.663962
R648 DEC2.n12 DEC2.n11 0.663962
R649 DEC2.n11 DEC2.n10 0.663962
R650 DEC2.n10 DEC2.n9 0.663962
R651 DEC2.n9 DEC2.n8 0.663962
R652 DEC2.n8 DEC2.n7 0.663962
R653 DEC2 DEC2.n6 0.65675
R654 rseg_4_routing_0/rseg_4_v3_0.v46 rseg_4_routing_0/rseg_4_v3_0.v46.t1 676.005
R655 rseg_4_routing_0/rseg_4_v3_0.v46.n0 rseg_4_routing_0/rseg_4_v3_0.v46.t0 10.7355
R656 rseg_4_routing_0/rseg_4_v3_0.v46.n0 rseg_4_routing_0/rseg_4_v3_0.v46.t2 10.6512
R657 rseg_4_routing_0/rseg_4_v3_0.v46 rseg_4_routing_0/rseg_4_v3_0.v46.n0 0.683611
R658 rseg_4_routing_0/rseg_4_v3_0.v51 rseg_4_routing_0/rseg_4_v3_0.v51.t1 672.309
R659 rseg_4_routing_0/rseg_4_v3_0.v51.n0 rseg_4_routing_0/rseg_4_v3_0.v51.t0 10.8249
R660 rseg_4_routing_0/rseg_4_v3_0.v51.n0 rseg_4_routing_0/rseg_4_v3_0.v51.t2 10.5739
R661 rseg_4_routing_0/rseg_4_v3_0.v51 rseg_4_routing_0/rseg_4_v3_0.v51.n0 1.38332
R662 rseg_4_routing_0/rseg_4_v3_0.v52 rseg_4_routing_0/rseg_4_v3_0.v52.t2 672.956
R663 rseg_4_routing_0/rseg_4_v3_0.v52.n0 rseg_4_routing_0/rseg_4_v3_0.v52.t0 10.717
R664 rseg_4_routing_0/rseg_4_v3_0.v52.n0 rseg_4_routing_0/rseg_4_v3_0.v52.t1 10.6712
R665 rseg_4_routing_0/rseg_4_v3_0.v52 rseg_4_routing_0/rseg_4_v3_0.v52.n0 2.0484
R666 rseg_4_routing_0/rseg_4_v3_0.v41 rseg_4_routing_0/rseg_4_v3_0.v41.t2 675.929
R667 rseg_4_routing_0/rseg_4_v3_0.v41.n0 rseg_4_routing_0/rseg_4_v3_0.v41.t1 10.8167
R668 rseg_4_routing_0/rseg_4_v3_0.v41.n0 rseg_4_routing_0/rseg_4_v3_0.v41.t0 10.6741
R669 rseg_4_routing_0/rseg_4_v3_0.v41 rseg_4_routing_0/rseg_4_v3_0.v41.n0 4.10816
R670 bb3.n0 bb3.t1 217.555
R671 bb3.n6 bb3.t7 216.893
R672 bb3.n5 bb3.t4 216.893
R673 bb3.n4 bb3.t5 216.893
R674 bb3.n3 bb3.t2 216.893
R675 bb3.n2 bb3.t0 216.893
R676 bb3.n1 bb3.t3 216.893
R677 bb3.n0 bb3.t6 216.893
R678 bb3.n1 bb3.n0 0.663962
R679 bb3.n2 bb3.n1 0.663962
R680 bb3.n3 bb3.n2 0.663962
R681 bb3.n4 bb3.n3 0.663962
R682 bb3.n5 bb3.n4 0.663962
R683 bb3.n6 bb3.n5 0.663962
R684 bb3 bb3.n6 0.293769
R685 a_35584_n5474.n0 a_35584_n5474.t1 671.409
R686 a_35584_n5474.n0 a_35584_n5474.t2 670.924
R687 a_35584_n5474.t0 a_35584_n5474.n0 665.707
R688 rseg_4_routing_0/rseg_4_v3_0.v55 rseg_4_routing_0/rseg_4_v3_0.v55.t1 674.658
R689 rseg_4_routing_0/rseg_4_v3_0.v55.n0 rseg_4_routing_0/rseg_4_v3_0.v55.t2 10.7625
R690 rseg_4_routing_0/rseg_4_v3_0.v55.n0 rseg_4_routing_0/rseg_4_v3_0.v55.t0 10.7309
R691 rseg_4_routing_0/rseg_4_v3_0.v55 rseg_4_routing_0/rseg_4_v3_0.v55.n0 4.09058
R692 rseg_4_routing_0/rseg_4_v3_0.v56 rseg_4_routing_0/rseg_4_v3_0.v56.t1 676.321
R693 rseg_4_routing_0/rseg_4_v3_0.v56.n0 rseg_4_routing_0/rseg_4_v3_0.v56.t0 13.5978
R694 rseg_4_routing_0/rseg_4_v3_0.v56.n0 rseg_4_routing_0/rseg_4_v3_0.v56.t2 10.7628
R695 rseg_4_routing_0/rseg_4_v3_0.v56 rseg_4_routing_0/rseg_4_v3_0.v56.n0 4.72836
R696 rseg_4_routing_0/rseg_4_v3_0.v43 rseg_4_routing_0/rseg_4_v3_0.v43.t1 675.533
R697 rseg_4_routing_0/rseg_4_v3_0.v43.n0 rseg_4_routing_0/rseg_4_v3_0.v43.t0 10.7605
R698 rseg_4_routing_0/rseg_4_v3_0.v43.n0 rseg_4_routing_0/rseg_4_v3_0.v43.t2 10.7175
R699 rseg_4_routing_0/rseg_4_v3_0.v43 rseg_4_routing_0/rseg_4_v3_0.v43.n0 2.73151
R700 rseg_4_routing_0/rseg_4_v3_0.v42 rseg_4_routing_0/rseg_4_v3_0.v42.t2 676.712
R701 rseg_4_routing_0/rseg_4_v3_0.v42.n0 rseg_4_routing_0/rseg_4_v3_0.v42.t0 10.7728
R702 rseg_4_routing_0/rseg_4_v3_0.v42.n0 rseg_4_routing_0/rseg_4_v3_0.v42.t1 10.6268
R703 rseg_4_routing_0/rseg_4_v3_0.v42 rseg_4_routing_0/rseg_4_v3_0.v42.n0 3.43316
R704 rseg_4_routing_0/rseg_4_v3_0.v37 rseg_4_routing_0/rseg_4_v3_0.v37.t2 673.212
R705 rseg_4_routing_0/rseg_4_v3_0.v37.n0 rseg_4_routing_0/rseg_4_v3_0.v37.t0 10.7577
R706 rseg_4_routing_0/rseg_4_v3_0.v37.n0 rseg_4_routing_0/rseg_4_v3_0.v37.t1 10.7161
R707 rseg_4_routing_0/rseg_4_v3_0.v37 rseg_4_routing_0/rseg_4_v3_0.v37.n0 2.72817
R708 rseg_4_routing_0/rseg_4_v3_0.v36 rseg_4_routing_0/rseg_4_v3_0.v36.t2 672.795
R709 rseg_4_routing_0/rseg_4_v3_0.v36.n0 rseg_4_routing_0/rseg_4_v3_0.v36.t1 10.7151
R710 rseg_4_routing_0/rseg_4_v3_0.v36.n0 rseg_4_routing_0/rseg_4_v3_0.v36.t0 10.6684
R711 rseg_4_routing_0/rseg_4_v3_0.v36 rseg_4_routing_0/rseg_4_v3_0.v36.n0 2.05222
R712 a_33357_n6738.t0 a_33357_n6738.n2 672.947
R713 a_33357_n6738.n0 a_33357_n6738.t1 671.573
R714 a_33357_n6738.n0 a_33357_n6738.t3 666.919
R715 a_33357_n6738.n2 a_33357_n6738.t2 666.46
R716 a_33357_n6738.n1 a_33357_n6738.t4 666.46
R717 a_33357_n6738.n2 a_33357_n6738.n1 6.63383
R718 a_33357_n6738.n1 a_33357_n6738.n0 1.84008
R719 rseg_4_routing_0/rseg_4_v3_0.v62.n0 rseg_4_routing_0/rseg_4_v3_0.v62.t1 676.833
R720 rseg_4_routing_0/rseg_4_v3_0.v62.n0 rseg_4_routing_0/rseg_4_v3_0.v62.t2 10.7929
R721 rseg_4_routing_0/rseg_4_v3_0.v62.t0 rseg_4_routing_0/rseg_4_v3_0.v62.n0 10.5295
R722 a_29969_n8174.n0 a_29969_n8174.t1 672.278
R723 a_29969_n8174.t0 a_29969_n8174.n2 671.904
R724 a_29969_n8174.n1 a_29969_n8174.t3 671.547
R725 a_29969_n8174.n2 a_29969_n8174.t2 665.484
R726 a_29969_n8174.n0 a_29969_n8174.t4 665.484
R727 a_29969_n8174.n1 a_29969_n8174.n0 4.99842
R728 a_29969_n8174.n2 a_29969_n8174.n1 1.563
R729 rseg_4_routing_0/rseg_4_v3_0.v33.t0 rseg_4_routing_0/rseg_4_v3_0.v33.n0 663.232
R730 rseg_4_routing_0/rseg_4_v3_0.v33.n0 rseg_4_routing_0/rseg_4_v3_0.v33.t2 10.6713
R731 rseg_4_routing_0/rseg_4_v3_0.v33.n0 rseg_4_routing_0/rseg_4_v3_0.v33.t1 10.5739
R732 bb1.n0 bb1.t1 217.555
R733 bb1.n0 bb1.t0 216.893
R734 bb1 bb1.n0 0.166365
R735 a_36266_n4393.n0 a_36266_n4393.t2 668.659
R736 a_36266_n4393.n0 a_36266_n4393.t1 668.024
R737 a_36266_n4393.t0 a_36266_n4393.n0 665.667
R738 rseg_4_routing_0/rseg_4_v3_0.v49.t0 rseg_4_routing_0/rseg_4_v3_0.v49.n0 663.232
R739 rseg_4_routing_0/rseg_4_v3_0.v49.n0 rseg_4_routing_0/rseg_4_v3_0.v49.t1 10.6701
R740 rseg_4_routing_0/rseg_4_v3_0.v49.n0 rseg_4_routing_0/rseg_4_v3_0.v49.t2 10.5739
R741 rseg_4_routing_0/rseg_4_v3_0.v50 rseg_4_routing_0/rseg_4_v3_0.v50.t0 673.491
R742 rseg_4_routing_0/rseg_4_v3_0.v50.n0 rseg_4_routing_0/rseg_4_v3_0.v50.t2 10.7472
R743 rseg_4_routing_0/rseg_4_v3_0.v50.n0 rseg_4_routing_0/rseg_4_v3_0.v50.t1 10.6526
R744 rseg_4_routing_0/rseg_4_v3_0.v50 rseg_4_routing_0/rseg_4_v3_0.v50.n0 0.679794
R745 a_30955_n8174.n0 a_30955_n8174.t1 672.827
R746 a_30955_n8174.t0 a_30955_n8174.n2 672.455
R747 a_30955_n8174.n1 a_30955_n8174.t3 671.236
R748 a_30955_n8174.n2 a_30955_n8174.t2 666.034
R749 a_30955_n8174.n0 a_30955_n8174.t4 666.034
R750 a_30955_n8174.n2 a_30955_n8174.n1 5.78175
R751 a_30955_n8174.n1 a_30955_n8174.n0 0.779667
R752 rseg_4_routing_0/rseg_4_v3_0.v32.n0 rseg_4_routing_0/rseg_4_v3_0.v32.t1 668.13
R753 rseg_4_routing_0/rseg_4_v3_0.v32.n0 rseg_4_routing_0/rseg_4_v3_0.v32.t2 12.1392
R754 rseg_4_routing_0/rseg_4_v3_0.v32.t0 rseg_4_routing_0/rseg_4_v3_0.v32.n0 12.0768
R755 bb2.n0 bb2.t0 217.555
R756 bb2.n2 bb2.t2 216.893
R757 bb2.n1 bb2.t1 216.893
R758 bb2.n0 bb2.t3 216.893
R759 bb2.n1 bb2.n0 0.663962
R760 bb2.n2 bb2.n1 0.663962
R761 bb2 bb2.n2 0.28175
R762 a_35990_n4393.n0 a_35990_n4393.t2 670.064
R763 a_35990_n4393.t0 a_35990_n4393.n0 668.208
R764 a_35990_n4393.n0 a_35990_n4393.t1 665.85
R765 V63.n0 V63.t1 667.769
R766 V63.n0 V63.t0 10.5739
R767 V63 V63.n0 2.44409
R768 DEC0.n7 DEC0.t2 217.555
R769 DEC0.n3 DEC0.t5 217.555
R770 DEC0.n0 DEC0.t10 217.555
R771 DEC0.n13 DEC0.t7 216.893
R772 DEC0.n12 DEC0.t15 216.893
R773 DEC0.n11 DEC0.t3 216.893
R774 DEC0.n10 DEC0.t8 216.893
R775 DEC0.n9 DEC0.t1 216.893
R776 DEC0.n8 DEC0.t11 216.893
R777 DEC0.n7 DEC0.t12 216.893
R778 DEC0.n3 DEC0.t4 216.893
R779 DEC0.n4 DEC0.t13 216.893
R780 DEC0.n5 DEC0.t0 216.893
R781 DEC0.n2 DEC0.t9 216.893
R782 DEC0.n1 DEC0.t14 216.893
R783 DEC0.n0 DEC0.t6 216.893
R784 DEC0.n14 DEC0.n6 7.0505
R785 DEC0.n14 DEC0.n13 5.78319
R786 DEC0.n8 DEC0.n7 0.663962
R787 DEC0.n9 DEC0.n8 0.663962
R788 DEC0.n10 DEC0.n9 0.663962
R789 DEC0.n11 DEC0.n10 0.663962
R790 DEC0.n12 DEC0.n11 0.663962
R791 DEC0.n13 DEC0.n12 0.663962
R792 DEC0.n5 DEC0.n4 0.663962
R793 DEC0.n4 DEC0.n3 0.663962
R794 DEC0.n1 DEC0.n0 0.663962
R795 DEC0.n2 DEC0.n1 0.663962
R796 DEC0.n6 DEC0.n5 0.320692
R797 DEC0.n6 DEC0.n2 0.320692
R798 DEC0 DEC0.n14 0.0755
R799 a_30521_n8174.n0 a_30521_n8174.t1 672.644
R800 a_30521_n8174.t0 a_30521_n8174.n2 672.27
R801 a_30521_n8174.n1 a_30521_n8174.t3 671.963
R802 a_30521_n8174.n2 a_30521_n8174.t2 665.85
R803 a_30521_n8174.n0 a_30521_n8174.t4 665.85
R804 a_30521_n8174.n1 a_30521_n8174.n0 5.78175
R805 a_30521_n8174.n2 a_30521_n8174.n1 0.779667
R806 rseg_4_routing_0/rseg_4_v3_0.v3 rseg_4_routing_0/rseg_4_v3_0.v3.t0 672.309
R807 rseg_4_routing_0/rseg_4_v3_0.v3.n0 rseg_4_routing_0/rseg_4_v3_0.v3.t2 10.791
R808 rseg_4_routing_0/rseg_4_v3_0.v3.n0 rseg_4_routing_0/rseg_4_v3_0.v3.t1 10.6937
R809 rseg_4_routing_0/rseg_4_v3_0.v3 rseg_4_routing_0/rseg_4_v3_0.v3.n0 1.35575
R810 rseg_4_routing_0/rseg_4_v3_0.v17.n0 rseg_4_routing_0/rseg_4_v3_0.v17.t1 663.232
R811 rseg_4_routing_0/rseg_4_v3_0.v17.n0 rseg_4_routing_0/rseg_4_v3_0.v17.t2 10.6713
R812 rseg_4_routing_0/rseg_4_v3_0.v17.t0 rseg_4_routing_0/rseg_4_v3_0.v17.n0 10.5739
R813 rseg_4_routing_0/rseg_4_v3_0.v27 rseg_4_routing_0/rseg_4_v3_0.v27.t1 675.533
R814 rseg_4_routing_0/rseg_4_v3_0.v27.n0 rseg_4_routing_0/rseg_4_v3_0.v27.t2 10.7601
R815 rseg_4_routing_0/rseg_4_v3_0.v27.n0 rseg_4_routing_0/rseg_4_v3_0.v27.t0 10.7161
R816 rseg_4_routing_0/rseg_4_v3_0.v27 rseg_4_routing_0/rseg_4_v3_0.v27.n0 2.73056
R817 rseg_4_routing_0/rseg_4_v3_0.v26 rseg_4_routing_0/rseg_4_v3_0.v26.t1 676.553
R818 rseg_4_routing_0/rseg_4_v3_0.v26.n0 rseg_4_routing_0/rseg_4_v3_0.v26.t0 10.7808
R819 rseg_4_routing_0/rseg_4_v3_0.v26.n0 rseg_4_routing_0/rseg_4_v3_0.v26.t2 10.6292
R820 rseg_4_routing_0/rseg_4_v3_0.v26 rseg_4_routing_0/rseg_4_v3_0.v26.n0 3.43637
R821 rseg_4_routing_0/rseg_4_v3_0.v2 rseg_4_routing_0/rseg_4_v3_0.v2.t0 673.192
R822 rseg_4_routing_0/rseg_4_v3_0.v2.n0 rseg_4_routing_0/rseg_4_v3_0.v2.t1 10.7568
R823 rseg_4_routing_0/rseg_4_v3_0.v2.n0 rseg_4_routing_0/rseg_4_v3_0.v2.t2 10.6535
R824 rseg_4_routing_0/rseg_4_v3_0.v2 rseg_4_routing_0/rseg_4_v3_0.v2.n0 0.67884
R825 rseg_4_routing_0/rseg_4_v3_0.v38 rseg_4_routing_0/rseg_4_v3_0.v38.t2 673.412
R826 rseg_4_routing_0/rseg_4_v3_0.v38.n0 rseg_4_routing_0/rseg_4_v3_0.v38.t1 10.7203
R827 rseg_4_routing_0/rseg_4_v3_0.v38.n0 rseg_4_routing_0/rseg_4_v3_0.v38.t0 10.6908
R828 rseg_4_routing_0/rseg_4_v3_0.v38 rseg_4_routing_0/rseg_4_v3_0.v38.n0 3.42178
R829 a_31507_n8174.n0 a_31507_n8174.t1 673.193
R830 a_31507_n8174.t0 a_31507_n8174.n2 672.821
R831 a_31507_n8174.n1 a_31507_n8174.t3 670.087
R832 a_31507_n8174.n2 a_31507_n8174.t2 666.399
R833 a_31507_n8174.n0 a_31507_n8174.t4 666.399
R834 a_31507_n8174.n2 a_31507_n8174.n1 4.99842
R835 a_31507_n8174.n1 a_31507_n8174.n0 1.563
R836 rseg_4_routing_0/rseg_4_v3_0.v53 rseg_4_routing_0/rseg_4_v3_0.v53.t2 673.212
R837 rseg_4_routing_0/rseg_4_v3_0.v53.n0 rseg_4_routing_0/rseg_4_v3_0.v53.t0 10.7613
R838 rseg_4_routing_0/rseg_4_v3_0.v53.n0 rseg_4_routing_0/rseg_4_v3_0.v53.t1 10.7113
R839 rseg_4_routing_0/rseg_4_v3_0.v53 rseg_4_routing_0/rseg_4_v3_0.v53.n0 2.72292
R840 rseg_4_routing_0/rseg_4_v3_0.v28 rseg_4_routing_0/rseg_4_v3_0.v28.t1 675.814
R841 rseg_4_routing_0/rseg_4_v3_0.v28.n0 rseg_4_routing_0/rseg_4_v3_0.v28.t0 10.7162
R842 rseg_4_routing_0/rseg_4_v3_0.v28.n0 rseg_4_routing_0/rseg_4_v3_0.v28.t2 10.6712
R843 rseg_4_routing_0/rseg_4_v3_0.v28 rseg_4_routing_0/rseg_4_v3_0.v28.n0 2.05317
R844 b2.n0 b2.t0 217.555
R845 b2.n0 b2.t3 216.893
R846 b2.n1 b2.t1 216.893
R847 b2.n2 b2.t2 216.893
R848 b2.n2 b2.n1 0.663962
R849 b2.n1 b2.n0 0.663962
R850 b2 b2.n2 0.180788
R851 a_34638_n5474.t0 a_34638_n5474.n0 670.153
R852 a_34638_n5474.n0 a_34638_n5474.t2 669.817
R853 a_34638_n5474.n0 a_34638_n5474.t1 666.441
R854 rseg_4_routing_0/rseg_4_v3_0.v12 rseg_4_routing_0/rseg_4_v3_0.v12.t0 675.741
R855 rseg_4_routing_0/rseg_4_v3_0.v12.n0 rseg_4_routing_0/rseg_4_v3_0.v12.t2 10.7126
R856 rseg_4_routing_0/rseg_4_v3_0.v12.n0 rseg_4_routing_0/rseg_4_v3_0.v12.t1 10.6722
R857 rseg_4_routing_0/rseg_4_v3_0.v12 rseg_4_routing_0/rseg_4_v3_0.v12.n0 2.0546
R858 a_30245_n8174.n0 a_30245_n8174.t1 672.461
R859 a_30245_n8174.t0 a_30245_n8174.n2 672.087
R860 a_30245_n8174.n1 a_30245_n8174.t3 671.755
R861 a_30245_n8174.n2 a_30245_n8174.t2 665.667
R862 a_30245_n8174.n0 a_30245_n8174.t4 665.667
R863 a_30245_n8174.n1 a_30245_n8174.n0 5.39008
R864 a_30245_n8174.n2 a_30245_n8174.n1 1.17133
R865 rseg_4_routing_0/rseg_4_v3_0.v18 rseg_4_routing_0/rseg_4_v3_0.v18.t1 673.259
R866 rseg_4_routing_0/rseg_4_v3_0.v18.n0 rseg_4_routing_0/rseg_4_v3_0.v18.t0 10.7378
R867 rseg_4_routing_0/rseg_4_v3_0.v18.n0 rseg_4_routing_0/rseg_4_v3_0.v18.t2 10.6521
R868 rseg_4_routing_0/rseg_4_v3_0.v18 rseg_4_routing_0/rseg_4_v3_0.v18.n0 0.682657
R869 rseg_4_routing_0/rseg_4_v3_0.v31.t0 rseg_4_routing_0/rseg_4_v3_0.v31.n0 667.052
R870 rseg_4_routing_0/rseg_4_v3_0.v31.n0 rseg_4_routing_0/rseg_4_v3_0.v31.t2 10.6713
R871 rseg_4_routing_0/rseg_4_v3_0.v31.n0 rseg_4_routing_0/rseg_4_v3_0.v31.t1 10.5739
R872 rseg_4_routing_0/rseg_4_v3_0.v15.t0 rseg_4_routing_0/rseg_4_v3_0.v15.n0 667.052
R873 rseg_4_routing_0/rseg_4_v3_0.v15.n0 rseg_4_routing_0/rseg_4_v3_0.v15.t2 10.6701
R874 rseg_4_routing_0/rseg_4_v3_0.v15.n0 rseg_4_routing_0/rseg_4_v3_0.v15.t1 10.5739
R875 a_31819_n6738.t0 a_31819_n6738.n2 672.03
R876 a_31819_n6738.n0 a_31819_n6738.t1 668.37
R877 a_31819_n6738.n0 a_31819_n6738.t3 666.942
R878 a_31819_n6738.n2 a_31819_n6738.t2 665.543
R879 a_31819_n6738.n1 a_31819_n6738.t4 665.543
R880 a_31819_n6738.n2 a_31819_n6738.n1 6.63383
R881 a_31819_n6738.n1 a_31819_n6738.n0 4.12758
R882 rseg_4_routing_0/rseg_4_v3_0.v10 rseg_4_routing_0/rseg_4_v3_0.v10.t0 676.48
R883 rseg_4_routing_0/rseg_4_v3_0.v10.n0 rseg_4_routing_0/rseg_4_v3_0.v10.t1 10.7826
R884 rseg_4_routing_0/rseg_4_v3_0.v10.n0 rseg_4_routing_0/rseg_4_v3_0.v10.t2 10.6316
R885 rseg_4_routing_0/rseg_4_v3_0.v10 rseg_4_routing_0/rseg_4_v3_0.v10.n0 3.43753
R886 rseg_4_routing_0/rseg_4_v3_0.v54 rseg_4_routing_0/rseg_4_v3_0.v54.t2 673.572
R887 rseg_4_routing_0/rseg_4_v3_0.v54.n0 rseg_4_routing_0/rseg_4_v3_0.v54.t1 10.7178
R888 rseg_4_routing_0/rseg_4_v3_0.v54.n0 rseg_4_routing_0/rseg_4_v3_0.v54.t0 10.6903
R889 rseg_4_routing_0/rseg_4_v3_0.v54 rseg_4_routing_0/rseg_4_v3_0.v54.n0 3.41701
R890 b0 b0.t0 217.225
R891 VOUT.n0 VOUT.t1 665.933
R892 VOUT.n0 VOUT.t0 665.299
R893 VOUT VOUT.n0 0.0755
R894 a_35190_n5474.t0 a_35190_n5474.n0 670.519
R895 a_35190_n5474.n0 a_35190_n5474.t2 670.183
R896 a_35190_n5474.n0 a_35190_n5474.t1 666.073
R897 rseg_4_routing_0/rseg_4_v3_0.v45 rseg_4_routing_0/rseg_4_v3_0.v45.t2 675.904
R898 rseg_4_routing_0/rseg_4_v3_0.v45.n0 rseg_4_routing_0/rseg_4_v3_0.v45.t0 10.7766
R899 rseg_4_routing_0/rseg_4_v3_0.v45.n0 rseg_4_routing_0/rseg_4_v3_0.v45.t1 10.6951
R900 rseg_4_routing_0/rseg_4_v3_0.v45 rseg_4_routing_0/rseg_4_v3_0.v45.n0 1.35956
R901 a_31231_n8174.n0 a_31231_n8174.t1 673.01
R902 a_31231_n8174.t0 a_31231_n8174.n2 672.638
R903 a_31231_n8174.n1 a_31231_n8174.t3 670.662
R904 a_31231_n8174.n2 a_31231_n8174.t2 666.216
R905 a_31231_n8174.n0 a_31231_n8174.t4 666.216
R906 a_31231_n8174.n2 a_31231_n8174.n1 5.39008
R907 a_31231_n8174.n1 a_31231_n8174.n0 1.17133
R908 rseg_4_routing_0/rseg_4_v3_0.v20 rseg_4_routing_0/rseg_4_v3_0.v20.t1 672.722
R909 rseg_4_routing_0/rseg_4_v3_0.v20.n0 rseg_4_routing_0/rseg_4_v3_0.v20.t2 10.7152
R910 rseg_4_routing_0/rseg_4_v3_0.v20.n0 rseg_4_routing_0/rseg_4_v3_0.v20.t0 10.6722
R911 rseg_4_routing_0/rseg_4_v3_0.v20 rseg_4_routing_0/rseg_4_v3_0.v20.n0 2.05317
R912 rseg_4_routing_0/rseg_4_v3_0.v23 rseg_4_routing_0/rseg_4_v3_0.v23.t1 674.658
R913 rseg_4_routing_0/rseg_4_v3_0.v23.n0 rseg_4_routing_0/rseg_4_v3_0.v23.t2 10.7661
R914 rseg_4_routing_0/rseg_4_v3_0.v23.n0 rseg_4_routing_0/rseg_4_v3_0.v23.t0 10.7361
R915 rseg_4_routing_0/rseg_4_v3_0.v23 rseg_4_routing_0/rseg_4_v3_0.v23.n0 4.09773
R916 rseg_4_routing_0/rseg_4_v3_0.v25 rseg_4_routing_0/rseg_4_v3_0.v25.t2 675.929
R917 rseg_4_routing_0/rseg_4_v3_0.v25.n0 rseg_4_routing_0/rseg_4_v3_0.v25.t1 10.8219
R918 rseg_4_routing_0/rseg_4_v3_0.v25.n0 rseg_4_routing_0/rseg_4_v3_0.v25.t0 10.6741
R919 rseg_4_routing_0/rseg_4_v3_0.v25 rseg_4_routing_0/rseg_4_v3_0.v25.n0 4.11026
R920 a_35382_n4393.n0 a_35382_n4393.t1 666.692
R921 a_35382_n4393.t0 a_35382_n4393.n0 666.317
R922 a_35382_n4393.n0 a_35382_n4393.t2 665.484
R923 a_36570_n4393.t0 a_36570_n4393.n0 667.841
R924 a_36570_n4393.n0 a_36570_n4393.t2 667.34
R925 a_36570_n4393.n0 a_36570_n4393.t1 665.484
R926 a_35466_n5474.t0 a_35466_n5474.n0 670.775
R927 a_35466_n5474.n0 a_35466_n5474.t2 670.366
R928 a_35466_n5474.n0 a_35466_n5474.t1 665.89
R929 a_32095_n6738.t0 a_32095_n6738.n2 672.213
R930 a_32095_n6738.n0 a_32095_n6738.t1 668.944
R931 a_32095_n6738.n0 a_32095_n6738.t3 666.405
R932 a_32095_n6738.n2 a_32095_n6738.t2 665.726
R933 a_32095_n6738.n1 a_32095_n6738.t4 665.726
R934 a_32095_n6738.n2 a_32095_n6738.n1 6.63383
R935 a_32095_n6738.n1 a_32095_n6738.n0 3.73592
R936 rseg_4_routing_0/rseg_4_v3_0.v58 rseg_4_routing_0/rseg_4_v3_0.v58.t1 677.236
R937 rseg_4_routing_0/rseg_4_v3_0.v58.n0 rseg_4_routing_0/rseg_4_v3_0.v58.t0 10.7544
R938 rseg_4_routing_0/rseg_4_v3_0.v58.n0 rseg_4_routing_0/rseg_4_v3_0.v58.t2 10.6216
R939 rseg_4_routing_0/rseg_4_v3_0.v58 rseg_4_routing_0/rseg_4_v3_0.v58.n0 3.42573
R940 rseg_4_routing_0/rseg_4_v3_0.v14 rseg_4_routing_0/rseg_4_v3_0.v14.t0 675.77
R941 rseg_4_routing_0/rseg_4_v3_0.v14.n0 rseg_4_routing_0/rseg_4_v3_0.v14.t1 10.7383
R942 rseg_4_routing_0/rseg_4_v3_0.v14.n0 rseg_4_routing_0/rseg_4_v3_0.v14.t2 10.6502
R943 rseg_4_routing_0/rseg_4_v3_0.v14 rseg_4_routing_0/rseg_4_v3_0.v14.n0 0.682179
R944 rseg_4_routing_0/rseg_4_v3_0.v44 rseg_4_routing_0/rseg_4_v3_0.v44.t1 675.975
R945 rseg_4_routing_0/rseg_4_v3_0.v44.n0 rseg_4_routing_0/rseg_4_v3_0.v44.t2 10.7153
R946 rseg_4_routing_0/rseg_4_v3_0.v44.n0 rseg_4_routing_0/rseg_4_v3_0.v44.t0 10.6746
R947 rseg_4_routing_0/rseg_4_v3_0.v44 rseg_4_routing_0/rseg_4_v3_0.v44.n0 2.05556
R948 a_35860_n5474.n0 a_35860_n5474.t1 671.561
R949 a_35860_n5474.n0 a_35860_n5474.t2 671.109
R950 a_35860_n5474.t0 a_35860_n5474.n0 665.524
R951 a_31267_n6738.t0 a_31267_n6738.n2 671.663
R952 a_31267_n6738.n0 a_31267_n6738.t3 668.203
R953 a_31267_n6738.n0 a_31267_n6738.t1 667.22
R954 a_31267_n6738.n2 a_31267_n6738.t2 665.176
R955 a_31267_n6738.n1 a_31267_n6738.t4 665.176
R956 a_31267_n6738.n2 a_31267_n6738.n1 6.63383
R957 a_31267_n6738.n1 a_31267_n6738.n0 4.91092
R958 rseg_4_routing_0/rseg_4_v3_0.v7 rseg_4_routing_0/rseg_4_v3_0.v7.t0 674.658
R959 rseg_4_routing_0/rseg_4_v3_0.v7.n0 rseg_4_routing_0/rseg_4_v3_0.v7.t1 10.7657
R960 rseg_4_routing_0/rseg_4_v3_0.v7.n0 rseg_4_routing_0/rseg_4_v3_0.v7.t2 10.7357
R961 rseg_4_routing_0/rseg_4_v3_0.v7 rseg_4_routing_0/rseg_4_v3_0.v7.n0 4.09773
R962 rseg_4_routing_0/rseg_4_v3_0.v8 rseg_4_routing_0/rseg_4_v3_0.v8.t0 676.321
R963 rseg_4_routing_0/rseg_4_v3_0.v8.n0 rseg_4_routing_0/rseg_4_v3_0.v8.t2 13.4532
R964 rseg_4_routing_0/rseg_4_v3_0.v8.n0 rseg_4_routing_0/rseg_4_v3_0.v8.t1 10.7771
R965 rseg_4_routing_0/rseg_4_v3_0.v8 rseg_4_routing_0/rseg_4_v3_0.v8.n0 4.72836
R966 a_29693_n8174.n0 a_29693_n8174.t1 672.093
R967 a_29693_n8174.t0 a_29693_n8174.n2 671.721
R968 a_29693_n8174.n1 a_29693_n8174.t3 671.35
R969 a_29693_n8174.n2 a_29693_n8174.t2 665.299
R970 a_29693_n8174.n0 a_29693_n8174.t4 665.299
R971 a_29693_n8174.n1 a_29693_n8174.n0 4.60675
R972 a_29693_n8174.n2 a_29693_n8174.n1 1.95467
R973 rseg_4_routing_0/rseg_4_v3_0.v34 rseg_4_routing_0/rseg_4_v3_0.v34.t0 673.332
R974 rseg_4_routing_0/rseg_4_v3_0.v34.n0 rseg_4_routing_0/rseg_4_v3_0.v34.t2 10.7383
R975 rseg_4_routing_0/rseg_4_v3_0.v34.n0 rseg_4_routing_0/rseg_4_v3_0.v34.t1 10.6478
R976 rseg_4_routing_0/rseg_4_v3_0.v34 rseg_4_routing_0/rseg_4_v3_0.v34.n0 0.682179
R977 rseg_4_routing_0/rseg_4_v3_0.v35 rseg_4_routing_0/rseg_4_v3_0.v35.t1 672.309
R978 rseg_4_routing_0/rseg_4_v3_0.v35.n0 rseg_4_routing_0/rseg_4_v3_0.v35.t0 10.7751
R979 rseg_4_routing_0/rseg_4_v3_0.v35.n0 rseg_4_routing_0/rseg_4_v3_0.v35.t2 10.6965
R980 rseg_4_routing_0/rseg_4_v3_0.v35 rseg_4_routing_0/rseg_4_v3_0.v35.n0 1.35813
R981 rseg_4_routing_0/rseg_4_v3_0.v24 rseg_4_routing_0/rseg_4_v3_0.v24.t1 676.321
R982 rseg_4_routing_0/rseg_4_v3_0.v24.n0 rseg_4_routing_0/rseg_4_v3_0.v24.t0 13.4709
R983 rseg_4_routing_0/rseg_4_v3_0.v24.n0 rseg_4_routing_0/rseg_4_v3_0.v24.t2 10.7776
R984 rseg_4_routing_0/rseg_4_v3_0.v24 rseg_4_routing_0/rseg_4_v3_0.v24.n0 4.72836
R985 rseg_4_routing_0/rseg_4_v3_0.v19 rseg_4_routing_0/rseg_4_v3_0.v19.t2 672.309
R986 rseg_4_routing_0/rseg_4_v3_0.v19.n0 rseg_4_routing_0/rseg_4_v3_0.v19.t0 10.7857
R987 rseg_4_routing_0/rseg_4_v3_0.v19.n0 rseg_4_routing_0/rseg_4_v3_0.v19.t1 10.6946
R988 rseg_4_routing_0/rseg_4_v3_0.v19 rseg_4_routing_0/rseg_4_v3_0.v19.n0 1.3567
R989 rseg_4_routing_0/rseg_4_v3_0.v11 rseg_4_routing_0/rseg_4_v3_0.v11.t0 675.533
R990 rseg_4_routing_0/rseg_4_v3_0.v11.n0 rseg_4_routing_0/rseg_4_v3_0.v11.t2 10.7625
R991 rseg_4_routing_0/rseg_4_v3_0.v11.n0 rseg_4_routing_0/rseg_4_v3_0.v11.t1 10.7161
R992 rseg_4_routing_0/rseg_4_v3_0.v11 rseg_4_routing_0/rseg_4_v3_0.v11.n0 2.72817
R993 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v13.t0 675.904
R994 rseg_4_routing_0/rseg_4_v3_0.v13.n0 rseg_4_routing_0/rseg_4_v3_0.v13.t2 10.7856
R995 rseg_4_routing_0/rseg_4_v3_0.v13.n0 rseg_4_routing_0/rseg_4_v3_0.v13.t1 10.6951
R996 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v13.n0 1.35718
R997 rseg_4_routing_0/rseg_4_v3_0.v6 rseg_4_routing_0/rseg_4_v3_0.v6.t0 673.273
R998 rseg_4_routing_0/rseg_4_v3_0.v6.n0 rseg_4_routing_0/rseg_4_v3_0.v6.t2 10.7798
R999 rseg_4_routing_0/rseg_4_v3_0.v6.n0 rseg_4_routing_0/rseg_4_v3_0.v6.t1 10.6292
R1000 rseg_4_routing_0/rseg_4_v3_0.v6 rseg_4_routing_0/rseg_4_v3_0.v6.n0 3.43753
R1001 rseg_4_routing_0/rseg_4_v3_0.v9 rseg_4_routing_0/rseg_4_v3_0.v9.t0 675.929
R1002 rseg_4_routing_0/rseg_4_v3_0.v9.n0 rseg_4_routing_0/rseg_4_v3_0.v9.t2 10.8299
R1003 rseg_4_routing_0/rseg_4_v3_0.v9.n0 rseg_4_routing_0/rseg_4_v3_0.v9.t1 10.6741
R1004 rseg_4_routing_0/rseg_4_v3_0.v9 rseg_4_routing_0/rseg_4_v3_0.v9.n0 4.11253
R1005 rseg_4_routing_0/rseg_4_v3_0.v4 rseg_4_routing_0/rseg_4_v3_0.v4.t0 672.655
R1006 rseg_4_routing_0/rseg_4_v3_0.v4.n0 rseg_4_routing_0/rseg_4_v3_0.v4.t1 10.7124
R1007 rseg_4_routing_0/rseg_4_v3_0.v4.n0 rseg_4_routing_0/rseg_4_v3_0.v4.t2 10.6712
R1008 rseg_4_routing_0/rseg_4_v3_0.v4 rseg_4_routing_0/rseg_4_v3_0.v4.n0 2.05317
R1009 a_36136_n5474.n0 a_36136_n5474.t1 671.744
R1010 a_36136_n5474.n0 a_36136_n5474.t2 671.292
R1011 a_36136_n5474.t0 a_36136_n5474.n0 665.34
R1012 rseg_4_routing_0/rseg_4_v3_0.v5 rseg_4_routing_0/rseg_4_v3_0.v5.t0 673.212
R1013 rseg_4_routing_0/rseg_4_v3_0.v5.n0 rseg_4_routing_0/rseg_4_v3_0.v5.t2 10.7631
R1014 rseg_4_routing_0/rseg_4_v3_0.v5.n0 rseg_4_routing_0/rseg_4_v3_0.v5.t1 10.7147
R1015 rseg_4_routing_0/rseg_4_v3_0.v5 rseg_4_routing_0/rseg_4_v3_0.v5.n0 2.72674
R1016 rseg_4_routing_0/rseg_4_v3_0.v16.n0 rseg_4_routing_0/rseg_4_v3_0.v16.t2 668.13
R1017 rseg_4_routing_0/rseg_4_v3_0.v16.n0 rseg_4_routing_0/rseg_4_v3_0.v16.t1 12.1225
R1018 rseg_4_routing_0/rseg_4_v3_0.v16.t0 rseg_4_routing_0/rseg_4_v3_0.v16.n0 12.0768
R1019 a_34914_n5474.t0 a_34914_n5474.n0 670.336
R1020 a_34914_n5474.n0 a_34914_n5474.t2 670
R1021 a_34914_n5474.n0 a_34914_n5474.t1 666.258
R1022 rseg_4_routing_0/rseg_4_v3_0.v21 rseg_4_routing_0/rseg_4_v3_0.v21.t1 673.212
R1023 rseg_4_routing_0/rseg_4_v3_0.v21.n0 rseg_4_routing_0/rseg_4_v3_0.v21.t0 10.7601
R1024 rseg_4_routing_0/rseg_4_v3_0.v21.n0 rseg_4_routing_0/rseg_4_v3_0.v21.t2 10.7161
R1025 rseg_4_routing_0/rseg_4_v3_0.v21 rseg_4_routing_0/rseg_4_v3_0.v21.n0 2.72817
R1026 rseg_4_routing_0/rseg_4_v3_0.v59 rseg_4_routing_0/rseg_4_v3_0.v59.t1 675.533
R1027 rseg_4_routing_0/rseg_4_v3_0.v59.n0 rseg_4_routing_0/rseg_4_v3_0.v59.t2 10.7636
R1028 rseg_4_routing_0/rseg_4_v3_0.v59.n0 rseg_4_routing_0/rseg_4_v3_0.v59.t0 10.7261
R1029 rseg_4_routing_0/rseg_4_v3_0.v59 rseg_4_routing_0/rseg_4_v3_0.v59.n0 2.74248
R1030 bb0 bb0.t0 217.225
R1031 rseg_4_routing_0/rseg_4_v3_0.v22 rseg_4_routing_0/rseg_4_v3_0.v22.t2 673.34
R1032 rseg_4_routing_0/rseg_4_v3_0.v22.n0 rseg_4_routing_0/rseg_4_v3_0.v22.t1 10.7207
R1033 rseg_4_routing_0/rseg_4_v3_0.v22.n0 rseg_4_routing_0/rseg_4_v3_0.v22.t0 10.6941
R1034 rseg_4_routing_0/rseg_4_v3_0.v22 rseg_4_routing_0/rseg_4_v3_0.v22.n0 3.42321
C0 rseg_4_routing_0/rseg_4_v3_0.v35 rseg_4_routing_0/rseg_4_v3_0.v37 1.57341f
C1 rseg_4_routing_0/rseg_4_v3_0.v34 rseg_4_routing_0/rseg_4_v3_0.v37 0.04811f
C2 rseg_4_routing_0/rseg_4_v3_0.v26 rseg_4_routing_0/rseg_4_v3_0.v39 1.47954f
C3 rseg_4_routing_0/rseg_4_v3_0.v5 VPB 0.06953f
C4 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v12 1.24994f
C5 rseg_4_routing_0/rseg_4_v3_0.v57 rseg_4_routing_0/rseg_4_v3_0.v58 1.26639f
C6 V63 rseg_4_routing_0/rseg_4_v3_0.v56 0.066f
C7 rseg_4_routing_0/rseg_4_v3_0.v19 VPB 0.04638f
C8 b3 VPB 1.47496f
C9 rseg_4_routing_0/rseg_4_v3_0.v18 VPB 0.07072f
C10 VPB rseg_4_routing_0/rseg_4_v3_0.v45 0.15933f
C11 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v14 1.2479f
C12 rseg_4_routing_0/rseg_4_v3_0.v52 DEC3 0.03404f
C13 rseg_4_routing_0/rseg_4_v3_0.v54 rseg_4_routing_0/rseg_4_v3_0.v56 1.93547f
C14 DEC0 rseg_4_routing_0/rseg_4_v3_0.v6 0.0908f
C15 rseg_4_routing_0/rseg_4_v3_0.v36 VPB 0.04651f
C16 rseg_4_routing_0/rseg_4_v3_0.v21 rseg_4_routing_0/rseg_4_v3_0.v12 0.02615f
C17 V0 rseg_4_routing_0/rseg_4_v3_0.v6 0.01245f
C18 rseg_4_routing_0/rseg_4_v3_0.v24 VPB 0.23425f
C19 rseg_4_routing_0/rseg_4_v3_0.v50 DEC3 0.05882f
C20 VPB rseg_4_routing_0/rseg_4_v3_0.v20 0.04651f
C21 rseg_4_routing_0/rseg_4_v3_0.v23 VPB 0.13306f
C22 rseg_4_routing_0/rseg_4_v3_0.v5 rseg_4_routing_0/rseg_4_v3_0.v2 0.04809f
C23 rseg_4_routing_0/rseg_4_v3_0.v10 VPB 0.14937f
C24 rseg_4_routing_0/rseg_4_v3_0.v59 rseg_4_routing_0/rseg_4_v3_0.v57 1.9819f
C25 rseg_4_routing_0/rseg_4_v3_0.v11 rseg_4_routing_0/rseg_4_v3_0.v4 0.02254f
C26 rseg_4_routing_0/rseg_4_v3_0.v52 rseg_4_routing_0/rseg_4_v3_0.v50 1.36438f
C27 rseg_4_routing_0/rseg_4_v3_0.v25 rseg_4_routing_0/rseg_4_v3_0.v27 1.97317f
C28 rseg_4_routing_0/rseg_4_v3_0.v42 VPB 0.14894f
C29 rseg_4_routing_0/rseg_4_v3_0.v44 rseg_4_routing_0/rseg_4_v3_0.v45 1.18866f
C30 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v9 0.08427f
C31 rseg_4_routing_0/rseg_4_v3_0.v41 rseg_4_routing_0/rseg_4_v3_0.v38 0.04735f
C32 rseg_4_routing_0/rseg_4_v3_0.v28 rseg_4_routing_0/rseg_4_v3_0.v25 0.02715f
C33 rseg_4_routing_0/rseg_4_v3_0.v51 VPB 0.04529f
C34 rseg_4_routing_0/rseg_4_v3_0.v55 VPB 0.13379f
C35 DEC2 rseg_4_routing_0/rseg_4_v3_0.v35 0.02948f
C36 rseg_4_routing_0/rseg_4_v3_0.v30 rseg_4_routing_0/rseg_4_v3_0.v35 0.02493f
C37 DEC2 rseg_4_routing_0/rseg_4_v3_0.v34 0.05843f
C38 rseg_4_routing_0/rseg_4_v3_0.v28 rseg_4_routing_0/rseg_4_v3_0.v37 0.02615f
C39 rseg_4_routing_0/rseg_4_v3_0.v27 rseg_4_routing_0/rseg_4_v3_0.v29 1.85343f
C40 rseg_4_routing_0/rseg_4_v3_0.v61 rseg_4_routing_0/rseg_4_v3_0.v56 0.21461f
C41 rseg_4_routing_0/rseg_4_v3_0.v40 rseg_4_routing_0/rseg_4_v3_0.v38 1.94253f
C42 DEC2 rseg_4_routing_0/rseg_4_v3_0.v41 0.16929f
C43 b2 VPB 0.7129f
C44 rseg_4_routing_0/rseg_4_v3_0.v57 V63 0.02856f
C45 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v11 1.85017f
C46 DEC0 rseg_4_routing_0/rseg_4_v3_0.v7 0.14755f
C47 V0 rseg_4_routing_0/rseg_4_v3_0.v7 0.28896f
C48 rseg_4_routing_0/rseg_4_v3_0.v28 rseg_4_routing_0/rseg_4_v3_0.v29 1.21733f
C49 DEC0 rseg_4_routing_0/rseg_4_v3_0.v3 0.03386f
C50 DEC2 rseg_4_routing_0/rseg_4_v3_0.v46 0.15972f
C51 rseg_4_routing_0/rseg_4_v3_0.v39 rseg_4_routing_0/rseg_4_v3_0.v35 0.05244f
C52 rseg_4_routing_0/rseg_4_v3_0.v39 rseg_4_routing_0/rseg_4_v3_0.v34 0.05772f
C53 rseg_4_routing_0/rseg_4_v3_0.v41 rseg_4_routing_0/rseg_4_v3_0.v43 1.97214f
C54 rseg_4_routing_0/rseg_4_v3_0.v57 rseg_4_routing_0/rseg_4_v3_0.v54 0.04626f
C55 rseg_4_routing_0/rseg_4_v3_0.v44 rseg_4_routing_0/rseg_4_v3_0.v42 2.14311f
C56 rseg_4_routing_0/rseg_4_v3_0.v3 V0 0.32257f
C57 rseg_4_routing_0/rseg_4_v3_0.v40 DEC2 0.27737f
C58 VPB b0 0.1849f
C59 rseg_4_routing_0/rseg_4_v3_0.v43 rseg_4_routing_0/rseg_4_v3_0.v46 0.0119f
C60 rseg_4_routing_0/rseg_4_v3_0.v6 rseg_4_routing_0/rseg_4_v3_0.v9 0.04788f
C61 DEC0 rseg_4_routing_0/rseg_4_v3_0.v8 0.18308f
C62 rseg_4_routing_0/rseg_4_v3_0.v26 VPB 0.14911f
C63 rseg_4_routing_0/rseg_4_v3_0.v44 rseg_4_routing_0/rseg_4_v3_0.v51 0.03397f
C64 DEC1 VPB 3.01934f
C65 rseg_4_routing_0/rseg_4_v3_0.v40 rseg_4_routing_0/rseg_4_v3_0.v43 0.10119f
C66 rseg_4_routing_0/rseg_4_v3_0.v42 DEC3 0.01131f
C67 rseg_4_routing_0/rseg_4_v3_0.v22 VPB 0.1372f
C68 rseg_4_routing_0/rseg_4_v3_0.v40 rseg_4_routing_0/rseg_4_v3_0.v39 0.13214f
C69 VOUT b0 0.10734f
C70 rseg_4_routing_0/rseg_4_v3_0.v4 VPB 0.04526f
C71 rseg_4_routing_0/rseg_4_v3_0.v60 rseg_4_routing_0/rseg_4_v3_0.v58 2.29207f
C72 rseg_4_routing_0/rseg_4_v3_0.v11 rseg_4_routing_0/rseg_4_v3_0.v6 0.05322f
C73 rseg_4_routing_0/rseg_4_v3_0.v51 DEC3 0.03386f
C74 rseg_4_routing_0/rseg_4_v3_0.v55 DEC3 0.14747f
C75 rseg_4_routing_0/rseg_4_v3_0.v19 rseg_4_routing_0/rseg_4_v3_0.v18 0.69667f
C76 rseg_4_routing_0/rseg_4_v3_0.v51 rseg_4_routing_0/rseg_4_v3_0.v52 0.5508f
C77 rseg_4_routing_0/rseg_4_v3_0.v52 rseg_4_routing_0/rseg_4_v3_0.v55 0.06152f
C78 rseg_4_routing_0/rseg_4_v3_0.v30 rseg_4_routing_0/rseg_4_v3_0.v27 0.0119f
C79 VPB rseg_4_routing_0/rseg_4_v3_0.v58 0.08966f
C80 bb0 VPB 0.19301f
C81 rseg_4_routing_0/rseg_4_v3_0.v57 rseg_4_routing_0/rseg_4_v3_0.v61 0.0847f
C82 rseg_4_routing_0/rseg_4_v3_0.v36 rseg_4_routing_0/rseg_4_v3_0.v45 0.02213f
C83 rseg_4_routing_0/rseg_4_v3_0.v30 rseg_4_routing_0/rseg_4_v3_0.v28 1.27523f
C84 rseg_4_routing_0/rseg_4_v3_0.v51 rseg_4_routing_0/rseg_4_v3_0.v50 0.63972f
C85 rseg_4_routing_0/rseg_4_v3_0.v50 rseg_4_routing_0/rseg_4_v3_0.v55 0.05787f
C86 rseg_4_routing_0/rseg_4_v3_0.v13 VPB 0.16077f
C87 rseg_4_routing_0/rseg_4_v3_0.v19 rseg_4_routing_0/rseg_4_v3_0.v20 0.60845f
C88 rseg_4_routing_0/rseg_4_v3_0.v24 rseg_4_routing_0/rseg_4_v3_0.v18 0.0119f
C89 rseg_4_routing_0/rseg_4_v3_0.v59 rseg_4_routing_0/rseg_4_v3_0.v60 1.28515f
C90 bb0 VOUT 0.16947f
C91 rseg_4_routing_0/rseg_4_v3_0.v19 rseg_4_routing_0/rseg_4_v3_0.v23 0.05253f
C92 rseg_4_routing_0/rseg_4_v3_0.v18 rseg_4_routing_0/rseg_4_v3_0.v20 1.33533f
C93 rseg_4_routing_0/rseg_4_v3_0.v18 rseg_4_routing_0/rseg_4_v3_0.v23 0.05765f
C94 bb1 b1 0.04348f
C95 rseg_4_routing_0/rseg_4_v3_0.v4 rseg_4_routing_0/rseg_4_v3_0.v2 1.32352f
C96 rseg_4_routing_0/rseg_4_v3_0.v42 rseg_4_routing_0/rseg_4_v3_0.v45 0.09546f
C97 rseg_4_routing_0/rseg_4_v3_0.v59 VPB 0.05733f
C98 rseg_4_routing_0/rseg_4_v3_0.v9 rseg_4_routing_0/rseg_4_v3_0.v8 4.14551f
C99 rseg_4_routing_0/rseg_4_v3_0.v25 rseg_4_routing_0/rseg_4_v3_0.v29 0.08427f
C100 rseg_4_routing_0/rseg_4_v3_0.v24 rseg_4_routing_0/rseg_4_v3_0.v23 0.16418f
C101 rseg_4_routing_0/rseg_4_v3_0.v21 VPB 0.0691f
C102 rseg_4_routing_0/rseg_4_v3_0.v23 rseg_4_routing_0/rseg_4_v3_0.v20 0.06107f
C103 rseg_4_routing_0/rseg_4_v3_0.v10 rseg_4_routing_0/rseg_4_v3_0.v23 1.47977f
C104 V63 rseg_4_routing_0/rseg_4_v3_0.v60 0.4405f
C105 DEC3 rseg_4_routing_0/rseg_4_v3_0.v58 0.18689f
C106 rseg_4_routing_0/rseg_4_v3_0.v53 VPB 0.06876f
C107 rseg_4_routing_0/rseg_4_v3_0.v6 VPB 0.13684f
C108 rseg_4_routing_0/rseg_4_v3_0.v35 VPB 0.04651f
C109 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v2 0.02199f
C110 rseg_4_routing_0/rseg_4_v3_0.v11 rseg_4_routing_0/rseg_4_v3_0.v8 0.10095f
C111 rseg_4_routing_0/rseg_4_v3_0.v34 VPB 0.07006f
C112 V63 VPB 0.12476f
C113 rseg_4_routing_0/rseg_4_v3_0.v41 VPB 0.20005f
C114 rseg_4_routing_0/rseg_4_v3_0.v54 VPB 0.14253f
C115 rseg_4_routing_0/rseg_4_v3_0.v42 rseg_4_routing_0/rseg_4_v3_0.v55 1.48f
C116 rseg_4_routing_0/rseg_4_v3_0.v5 rseg_4_routing_0/rseg_4_v3_0.v4 0.61579f
C117 DEC1 rseg_4_routing_0/rseg_4_v3_0.v19 0.02948f
C118 VPB rseg_4_routing_0/rseg_4_v3_0.v46 0.21507f
C119 DEC1 rseg_4_routing_0/rseg_4_v3_0.v18 0.0583f
C120 rseg_4_routing_0/rseg_4_v3_0.v40 VPB 0.22957f
C121 rseg_4_routing_0/rseg_4_v3_0.v38 rseg_4_routing_0/rseg_4_v3_0.v37 0.4555f
C122 rseg_4_routing_0/rseg_4_v3_0.v59 DEC3 0.09426f
C123 rseg_4_routing_0/rseg_4_v3_0.v51 rseg_4_routing_0/rseg_4_v3_0.v55 0.05244f
C124 rseg_4_routing_0/rseg_4_v3_0.v59 rseg_4_routing_0/rseg_4_v3_0.v52 0.02139f
C125 rseg_4_routing_0/rseg_4_v3_0.v44 rseg_4_routing_0/rseg_4_v3_0.v53 0.02665f
C126 DEC2 rseg_4_routing_0/rseg_4_v3_0.v37 0.05823f
C127 DEC1 rseg_4_routing_0/rseg_4_v3_0.v24 0.31576f
C128 rseg_4_routing_0/rseg_4_v3_0.v26 rseg_4_routing_0/rseg_4_v3_0.v24 0.5557f
C129 DEC1 rseg_4_routing_0/rseg_4_v3_0.v20 0.03009f
C130 VPB rseg_4_routing_0/rseg_4_v3_0.v7 0.13207f
C131 DEC1 rseg_4_routing_0/rseg_4_v3_0.v23 0.14826f
C132 rseg_4_routing_0/rseg_4_v3_0.v44 rseg_4_routing_0/rseg_4_v3_0.v41 0.02715f
C133 DEC1 rseg_4_routing_0/rseg_4_v3_0.v10 0.01142f
C134 rseg_4_routing_0/rseg_4_v3_0.v61 rseg_4_routing_0/rseg_4_v3_0.v60 1.15198f
C135 rseg_4_routing_0/rseg_4_v3_0.v53 DEC3 0.05833f
C136 DEC0 V0 0.05523f
C137 rseg_4_routing_0/rseg_4_v3_0.v3 VPB 0.04526f
C138 rseg_4_routing_0/rseg_4_v3_0.v24 rseg_4_routing_0/rseg_4_v3_0.v22 1.95068f
C139 rseg_4_routing_0/rseg_4_v3_0.v22 rseg_4_routing_0/rseg_4_v3_0.v20 1.81035f
C140 rseg_4_routing_0/rseg_4_v3_0.v22 rseg_4_routing_0/rseg_4_v3_0.v23 0.64353f
C141 rseg_4_routing_0/rseg_4_v3_0.v52 rseg_4_routing_0/rseg_4_v3_0.v53 0.53572f
C142 V63 DEC3 0.14757f
C143 rseg_4_routing_0/rseg_4_v3_0.v44 rseg_4_routing_0/rseg_4_v3_0.v46 1.27501f
C144 rseg_4_routing_0/rseg_4_v3_0.v30 rseg_4_routing_0/rseg_4_v3_0.v29 1.22509f
C145 rseg_4_routing_0/rseg_4_v3_0.v27 VPB 0.11272f
C146 rseg_4_routing_0/rseg_4_v3_0.v61 VPB 0.09479f
C147 DEC0 rseg_4_routing_0/rseg_4_v3_0.v12 0.09244f
C148 rseg_4_routing_0/rseg_4_v3_0.v39 rseg_4_routing_0/rseg_4_v3_0.v37 2.15445f
C149 rseg_4_routing_0/rseg_4_v3_0.v57 rseg_4_routing_0/rseg_4_v3_0.v56 4.16288f
C150 VPB rseg_4_routing_0/rseg_4_v3_0.v8 0.27086f
C151 rseg_4_routing_0/rseg_4_v3_0.v54 DEC3 0.0997f
C152 rseg_4_routing_0/rseg_4_v3_0.v50 rseg_4_routing_0/rseg_4_v3_0.v53 0.04809f
C153 rseg_4_routing_0/rseg_4_v3_0.v28 VPB 0.11006f
C154 DEC3 rseg_4_routing_0/rseg_4_v3_0.v46 0.02072f
C155 rseg_4_routing_0/rseg_4_v3_0.v52 rseg_4_routing_0/rseg_4_v3_0.v54 1.83395f
C156 DEC0 rseg_4_routing_0/rseg_4_v3_0.v14 0.15976f
C157 V63 rseg_4_routing_0/rseg_4_v3_0.v50 0.02253f
C158 rseg_4_routing_0/rseg_4_v3_0.v7 rseg_4_routing_0/rseg_4_v3_0.v2 0.05759f
C159 rseg_4_routing_0/rseg_4_v3_0.v5 rseg_4_routing_0/rseg_4_v3_0.v6 0.5188f
C160 rseg_4_routing_0/rseg_4_v3_0.v21 rseg_4_routing_0/rseg_4_v3_0.v19 1.57642f
C161 rseg_4_routing_0/rseg_4_v3_0.v12 rseg_4_routing_0/rseg_4_v3_0.v14 1.27264f
C162 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v10 0.09544f
C163 rseg_4_routing_0/rseg_4_v3_0.v3 rseg_4_routing_0/rseg_4_v3_0.v2 0.71512f
C164 rseg_4_routing_0/rseg_4_v3_0.v21 rseg_4_routing_0/rseg_4_v3_0.v18 0.04843f
C165 DEC2 rseg_4_routing_0/rseg_4_v3_0.v38 0.09406f
C166 VPB bb2 0.73485f
C167 DEC1 rseg_4_routing_0/rseg_4_v3_0.v26 0.18677f
C168 rseg_4_routing_0/rseg_4_v3_0.v43 rseg_4_routing_0/rseg_4_v3_0.v38 0.05322f
C169 rseg_4_routing_0/rseg_4_v3_0.v34 rseg_4_routing_0/rseg_4_v3_0.v45 0.02163f
C170 rseg_4_routing_0/rseg_4_v3_0.v8 rseg_4_routing_0/rseg_4_v3_0.v2 0.0119f
C171 rseg_4_routing_0/rseg_4_v3_0.v30 DEC2 0.02141f
C172 DEC1 rseg_4_routing_0/rseg_4_v3_0.v22 0.09604f
C173 rseg_4_routing_0/rseg_4_v3_0.v61 DEC3 0.18664f
C174 DEC0 rseg_4_routing_0/rseg_4_v3_0.v9 0.16773f
C175 rseg_4_routing_0/rseg_4_v3_0.v39 rseg_4_routing_0/rseg_4_v3_0.v38 0.6218f
C176 rseg_4_routing_0/rseg_4_v3_0.v41 rseg_4_routing_0/rseg_4_v3_0.v45 0.08427f
C177 rseg_4_routing_0/rseg_4_v3_0.v21 rseg_4_routing_0/rseg_4_v3_0.v20 0.59731f
C178 rseg_4_routing_0/rseg_4_v3_0.v21 rseg_4_routing_0/rseg_4_v3_0.v23 2.15145f
C179 rseg_4_routing_0/rseg_4_v3_0.v61 rseg_4_routing_0/rseg_4_v3_0.v52 0.02116f
C180 rseg_4_routing_0/rseg_4_v3_0.v35 rseg_4_routing_0/rseg_4_v3_0.v36 0.578f
C181 rseg_4_routing_0/rseg_4_v3_0.v21 rseg_4_routing_0/rseg_4_v3_0.v10 0.02726f
C182 bb0 b0 0.04348f
C183 rseg_4_routing_0/rseg_4_v3_0.v36 rseg_4_routing_0/rseg_4_v3_0.v34 1.3376f
C184 DEC2 rseg_4_routing_0/rseg_4_v3_0.v43 0.09729f
C185 rseg_4_routing_0/rseg_4_v3_0.v46 rseg_4_routing_0/rseg_4_v3_0.v45 1.19314f
C186 rseg_4_routing_0/rseg_4_v3_0.v12 rseg_4_routing_0/rseg_4_v3_0.v9 0.02715f
C187 rseg_4_routing_0/rseg_4_v3_0.v40 rseg_4_routing_0/rseg_4_v3_0.v45 0.21475f
C188 DEC2 rseg_4_routing_0/rseg_4_v3_0.v39 0.14802f
C189 DEC0 rseg_4_routing_0/rseg_4_v3_0.v11 0.10225f
C190 rseg_4_routing_0/rseg_4_v3_0.v30 rseg_4_routing_0/rseg_4_v3_0.v39 0.01649f
C191 VPB b1 0.35495f
C192 rseg_4_routing_0/rseg_4_v3_0.v42 rseg_4_routing_0/rseg_4_v3_0.v53 0.02775f
C193 rseg_4_routing_0/rseg_4_v3_0.v61 rseg_4_routing_0/rseg_4_v3_0.v50 0.02163f
C194 rseg_4_routing_0/rseg_4_v3_0.v5 rseg_4_routing_0/rseg_4_v3_0.v7 2.15109f
C195 rseg_4_routing_0/rseg_4_v3_0.v5 rseg_4_routing_0/rseg_4_v3_0.v3 1.57251f
C196 rseg_4_routing_0/rseg_4_v3_0.v51 rseg_4_routing_0/rseg_4_v3_0.v53 1.5609f
C197 rseg_4_routing_0/rseg_4_v3_0.v11 rseg_4_routing_0/rseg_4_v3_0.v12 1.37192f
C198 rseg_4_routing_0/rseg_4_v3_0.v55 rseg_4_routing_0/rseg_4_v3_0.v53 2.1375f
C199 rseg_4_routing_0/rseg_4_v3_0.v42 rseg_4_routing_0/rseg_4_v3_0.v41 1.3027f
C200 rseg_4_routing_0/rseg_4_v3_0.v42 rseg_4_routing_0/rseg_4_v3_0.v46 0.3835f
C201 rseg_4_routing_0/rseg_4_v3_0.v25 VPB 0.20041f
C202 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v4 0.02197f
C203 rseg_4_routing_0/rseg_4_v3_0.v42 rseg_4_routing_0/rseg_4_v3_0.v40 0.5556f
C204 rseg_4_routing_0/rseg_4_v3_0.v11 rseg_4_routing_0/rseg_4_v3_0.v14 0.0119f
C205 rseg_4_routing_0/rseg_4_v3_0.v37 VPB 0.06876f
C206 rseg_4_routing_0/rseg_4_v3_0.v54 rseg_4_routing_0/rseg_4_v3_0.v55 0.58839f
C207 rseg_4_routing_0/rseg_4_v3_0.v51 rseg_4_routing_0/rseg_4_v3_0.v46 0.02537f
C208 rseg_4_routing_0/rseg_4_v3_0.v55 rseg_4_routing_0/rseg_4_v3_0.v46 0.01646f
C209 DEC1 rseg_4_routing_0/rseg_4_v3_0.v21 0.05816f
C210 rseg_4_routing_0/rseg_4_v3_0.v40 rseg_4_routing_0/rseg_4_v3_0.v55 0.0672f
C211 rseg_4_routing_0/rseg_4_v3_0.v29 VPB 0.16165f
C212 rseg_4_routing_0/rseg_4_v3_0.v56 VPB 0.17616f
C213 bb1 VPB 0.3629f
C214 rseg_4_routing_0/rseg_4_v3_0.v21 rseg_4_routing_0/rseg_4_v3_0.v22 0.48603f
C215 rseg_4_routing_0/rseg_4_v3_0.v59 rseg_4_routing_0/rseg_4_v3_0.v58 1.27914f
C216 rseg_4_routing_0/rseg_4_v3_0.v24 rseg_4_routing_0/rseg_4_v3_0.v27 0.10107f
C217 rseg_4_routing_0/rseg_4_v3_0.v27 rseg_4_routing_0/rseg_4_v3_0.v20 0.02218f
C218 DEC0 VPB 3.01878f
C219 rseg_4_routing_0/rseg_4_v3_0.v23 rseg_4_routing_0/rseg_4_v3_0.v8 0.06862f
C220 rseg_4_routing_0/rseg_4_v3_0.v4 rseg_4_routing_0/rseg_4_v3_0.v6 1.79741f
C221 rseg_4_routing_0/rseg_4_v3_0.v10 rseg_4_routing_0/rseg_4_v3_0.v8 0.55111f
C222 rseg_4_routing_0/rseg_4_v3_0.v11 rseg_4_routing_0/rseg_4_v3_0.v9 1.96808f
C223 V0 VPB 0.11923f
C224 rseg_4_routing_0/rseg_4_v3_0.v12 VPB 0.10974f
C225 V63 rseg_4_routing_0/rseg_4_v3_0.v58 0.2465f
C226 rseg_4_routing_0/rseg_4_v3_0.v38 VPB 0.13931f
C227 rseg_4_routing_0/rseg_4_v3_0.v57 rseg_4_routing_0/rseg_4_v3_0.v60 0.02715f
C228 rseg_4_routing_0/rseg_4_v3_0.v14 VPB 0.22406f
C229 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v6 0.02015f
C230 DEC2 VPB 3.02655f
C231 rseg_4_routing_0/rseg_4_v3_0.v56 DEC3 0.18009f
C232 rseg_4_routing_0/rseg_4_v3_0.v30 VPB 0.21415f
C233 rseg_4_routing_0/rseg_4_v3_0.v57 VPB 0.14518f
C234 DEC0 rseg_4_routing_0/rseg_4_v3_0.v2 0.05832f
C235 rseg_4_routing_0/rseg_4_v3_0.v43 VPB 0.11246f
C236 V0 rseg_4_routing_0/rseg_4_v3_0.v2 0.95873f
C237 rseg_4_routing_0/rseg_4_v3_0.v4 rseg_4_routing_0/rseg_4_v3_0.v7 0.06095f
C238 rseg_4_routing_0/rseg_4_v3_0.v26 rseg_4_routing_0/rseg_4_v3_0.v27 1.34745f
C239 DEC1 rseg_4_routing_0/rseg_4_v3_0.v27 0.09942f
C240 rseg_4_routing_0/rseg_4_v3_0.v59 V63 0.02312f
C241 rseg_4_routing_0/rseg_4_v3_0.v3 rseg_4_routing_0/rseg_4_v3_0.v4 0.64115f
C242 rseg_4_routing_0/rseg_4_v3_0.v39 VPB 0.13352f
C243 rseg_4_routing_0/rseg_4_v3_0.v50 rseg_4_routing_0/rseg_4_v3_0.v56 0.0119f
C244 rseg_4_routing_0/rseg_4_v3_0.v22 rseg_4_routing_0/rseg_4_v3_0.v27 0.05305f
C245 rseg_4_routing_0/rseg_4_v3_0.v26 rseg_4_routing_0/rseg_4_v3_0.v28 2.09546f
C246 b2 bb2 0.04424f
C247 DEC1 rseg_4_routing_0/rseg_4_v3_0.v28 0.09239f
C248 rseg_4_routing_0/rseg_4_v3_0.v59 rseg_4_routing_0/rseg_4_v3_0.v54 0.05213f
C249 VPB rseg_4_routing_0/rseg_4_v3_0.v9 0.20049f
C250 rseg_4_routing_0/rseg_4_v3_0.v44 DEC2 0.09236f
C251 rseg_4_routing_0/rseg_4_v3_0.v61 rseg_4_routing_0/rseg_4_v3_0.v58 0.0953f
C252 rseg_4_routing_0/rseg_4_v3_0.v35 rseg_4_routing_0/rseg_4_v3_0.v34 0.6765f
C253 rseg_4_routing_0/rseg_4_v3_0.v44 rseg_4_routing_0/rseg_4_v3_0.v43 1.32046f
C254 rseg_4_routing_0/rseg_4_v3_0.v18 rseg_4_routing_0/rseg_4_v3_0.v29 0.02156f
C255 rseg_4_routing_0/rseg_4_v3_0.v36 rseg_4_routing_0/rseg_4_v3_0.v37 0.57187f
C256 rseg_4_routing_0/rseg_4_v3_0.v54 rseg_4_routing_0/rseg_4_v3_0.v53 0.4235f
C257 DEC2 DEC3 0.01879f
C258 rseg_4_routing_0/rseg_4_v3_0.v11 VPB 0.11236f
C259 rseg_4_routing_0/rseg_4_v3_0.v25 rseg_4_routing_0/rseg_4_v3_0.v24 4.13148f
C260 rseg_4_routing_0/rseg_4_v3_0.v5 DEC0 0.0582f
C261 rseg_4_routing_0/rseg_4_v3_0.v57 DEC3 0.16656f
C262 rseg_4_routing_0/rseg_4_v3_0.v5 V0 0.23408f
C263 b2 b1 0.04424f
C264 rseg_4_routing_0/rseg_4_v3_0.v13 rseg_4_routing_0/rseg_4_v3_0.v8 0.21361f
C265 rseg_4_routing_0/rseg_4_v3_0.v40 rseg_4_routing_0/rseg_4_v3_0.v34 0.0119f
C266 rseg_4_routing_0/rseg_4_v3_0.v59 rseg_4_routing_0/rseg_4_v3_0.v61 1.8611f
C267 rseg_4_routing_0/rseg_4_v3_0.v24 rseg_4_routing_0/rseg_4_v3_0.v29 0.21451f
C268 rseg_4_routing_0/rseg_4_v3_0.v29 rseg_4_routing_0/rseg_4_v3_0.v20 0.02197f
C269 rseg_4_routing_0/rseg_4_v3_0.v40 rseg_4_routing_0/rseg_4_v3_0.v41 4.12073f
C270 rseg_4_routing_0/rseg_4_v3_0.v6 rseg_4_routing_0/rseg_4_v3_0.v7 0.66863f
C271 rseg_4_routing_0/rseg_4_v3_0.v19 rseg_4_routing_0/rseg_4_v3_0.v12 0.03375f
C272 rseg_4_routing_0/rseg_4_v3_0.v38 rseg_4_routing_0/rseg_4_v3_0.v45 0.02015f
C273 rseg_4_routing_0/rseg_4_v3_0.v55 rseg_4_routing_0/rseg_4_v3_0.v56 0.0921f
C274 rseg_4_routing_0/rseg_4_v3_0.v19 rseg_4_routing_0/rseg_4_v3_0.v14 0.02523f
C275 DEC0 rseg_4_routing_0/rseg_4_v3_0.v10 0.1869f
C276 rseg_4_routing_0/rseg_4_v3_0.v36 rseg_4_routing_0/rseg_4_v3_0.v38 1.81409f
C277 V63 rseg_4_routing_0/rseg_4_v3_0.v61 0.88774f
C278 DEC2 rseg_4_routing_0/rseg_4_v3_0.v45 0.18633f
C279 rseg_4_routing_0/rseg_4_v3_0.v6 rseg_4_routing_0/rseg_4_v3_0.v8 1.95031f
C280 rseg_4_routing_0/rseg_4_v3_0.v60 VPB 0.05229f
C281 rseg_4_routing_0/rseg_4_v3_0.v28 rseg_4_routing_0/rseg_4_v3_0.v35 0.03419f
C282 rseg_4_routing_0/rseg_4_v3_0.v26 rseg_4_routing_0/rseg_4_v3_0.v25 1.33058f
C283 DEC1 rseg_4_routing_0/rseg_4_v3_0.v25 0.16949f
C284 rseg_4_routing_0/rseg_4_v3_0.v12 rseg_4_routing_0/rseg_4_v3_0.v10 2.07729f
C285 rseg_4_routing_0/rseg_4_v3_0.v61 rseg_4_routing_0/rseg_4_v3_0.v54 0.02015f
C286 rseg_4_routing_0/rseg_4_v3_0.v43 rseg_4_routing_0/rseg_4_v3_0.v45 1.85532f
C287 DEC2 rseg_4_routing_0/rseg_4_v3_0.v36 0.03011f
C288 rseg_4_routing_0/rseg_4_v3_0.v26 rseg_4_routing_0/rseg_4_v3_0.v37 0.02748f
C289 rseg_4_routing_0/rseg_4_v3_0.v25 rseg_4_routing_0/rseg_4_v3_0.v22 0.04751f
C290 rseg_4_routing_0/rseg_4_v3_0.v14 rseg_4_routing_0/rseg_4_v3_0.v23 0.01651f
C291 bb1 b0 0.04348f
C292 rseg_4_routing_0/rseg_4_v3_0.v10 rseg_4_routing_0/rseg_4_v3_0.v14 0.31886f
C293 rseg_4_routing_0/rseg_4_v3_0.v43 rseg_4_routing_0/rseg_4_v3_0.v36 0.02218f
C294 DEC1 rseg_4_routing_0/rseg_4_v3_0.v29 0.18775f
C295 rseg_4_routing_0/rseg_4_v3_0.v26 rseg_4_routing_0/rseg_4_v3_0.v29 0.09546f
C296 rseg_4_routing_0/rseg_4_v3_0.v42 DEC2 0.18667f
C297 rseg_4_routing_0/rseg_4_v3_0.v3 rseg_4_routing_0/rseg_4_v3_0.v7 0.05244f
C298 rseg_4_routing_0/rseg_4_v3_0.v39 rseg_4_routing_0/rseg_4_v3_0.v36 0.06121f
C299 VOUT VPB 0.17791f
C300 rseg_4_routing_0/rseg_4_v3_0.v22 rseg_4_routing_0/rseg_4_v3_0.v29 0.02015f
C301 rseg_4_routing_0/rseg_4_v3_0.v39 rseg_4_routing_0/rseg_4_v3_0.v24 0.06886f
C302 rseg_4_routing_0/rseg_4_v3_0.v42 rseg_4_routing_0/rseg_4_v3_0.v43 1.3157f
C303 rseg_4_routing_0/rseg_4_v3_0.v8 rseg_4_routing_0/rseg_4_v3_0.v7 0.19295f
C304 rseg_4_routing_0/rseg_4_v3_0.v44 VPB 0.10926f
C305 rseg_4_routing_0/rseg_4_v3_0.v56 rseg_4_routing_0/rseg_4_v3_0.v58 0.54952f
C306 VPB rseg_4_routing_0/rseg_4_v3_0.v2 0.06872f
C307 rseg_4_routing_0/rseg_4_v3_0.v60 DEC3 0.09419f
C308 DEC0 rseg_4_routing_0/rseg_4_v3_0.v4 0.03422f
C309 rseg_4_routing_0/rseg_4_v3_0.v10 rseg_4_routing_0/rseg_4_v3_0.v9 1.3467f
C310 bb3 VPB 1.49092f
C311 rseg_4_routing_0/rseg_4_v3_0.v28 rseg_4_routing_0/rseg_4_v3_0.v27 1.34913f
C312 V0 rseg_4_routing_0/rseg_4_v3_0.v4 0.01764f
C313 DEC3 VPB 3.14208f
C314 rseg_4_routing_0/rseg_4_v3_0.v52 VPB 0.04529f
C315 DEC1 rseg_4_routing_0/rseg_4_v3_0.v14 0.02181f
C316 rseg_4_routing_0/rseg_4_v3_0.v26 DEC2 0.01138f
C317 rseg_4_routing_0/rseg_4_v3_0.v11 rseg_4_routing_0/rseg_4_v3_0.v10 1.3734f
C318 rseg_4_routing_0/rseg_4_v3_0.v30 rseg_4_routing_0/rseg_4_v3_0.v26 0.33918f
C319 rseg_4_routing_0/rseg_4_v3_0.v30 DEC1 0.15973f
C320 rseg_4_routing_0/rseg_4_v3_0.v59 rseg_4_routing_0/rseg_4_v3_0.v56 0.10213f
C321 rseg_4_routing_0/rseg_4_v3_0.v50 VPB 0.06892f
C322 DEC0 rseg_4_routing_0/rseg_4_v3_0.v13 0.19025f
C323 V0 GND 1.16344f
C324 V63 GND 2.20044f
C325 DEC3 GND 2.74984f
C326 DEC2 GND 1.9935f
C327 DEC1 GND 1.95634f
C328 DEC0 GND 2.30137f
C329 bb3 GND 0.95974f
C330 b3 GND 0.89639f
C331 VOUT GND 0.16049f
C332 bb2 GND 0.47591f
C333 b2 GND 0.4457f
C334 b1 GND 0.2124f
C335 bb1 GND 0.21534f
C336 b0 GND 0.11297f
C337 bb0 GND 0.13354f
C338 VPB GND 78.93223f
C339 rseg_4_routing_0/rseg_4_v3_0.v55 GND 1.89898f
C340 rseg_4_routing_0/rseg_4_v3_0.v54 GND 0.92879f
C341 rseg_4_routing_0/rseg_4_v3_0.v53 GND 1.14314f
C342 rseg_4_routing_0/rseg_4_v3_0.v52 GND 0.8323f
C343 rseg_4_routing_0/rseg_4_v3_0.v51 GND 0.71956f
C344 rseg_4_routing_0/rseg_4_v3_0.v50 GND 0.79316f
C345 rseg_4_routing_0/rseg_4_v3_0.v39 GND 1.88679f
C346 rseg_4_routing_0/rseg_4_v3_0.v38 GND 0.87481f
C347 rseg_4_routing_0/rseg_4_v3_0.v37 GND 1.12833f
C348 rseg_4_routing_0/rseg_4_v3_0.v36 GND 0.79452f
C349 rseg_4_routing_0/rseg_4_v3_0.v35 GND 0.69232f
C350 rseg_4_routing_0/rseg_4_v3_0.v34 GND 0.75887f
C351 rseg_4_routing_0/rseg_4_v3_0.v23 GND 1.868f
C352 rseg_4_routing_0/rseg_4_v3_0.v22 GND 0.85453f
C353 rseg_4_routing_0/rseg_4_v3_0.v21 GND 1.11257f
C354 rseg_4_routing_0/rseg_4_v3_0.v20 GND 0.77008f
C355 rseg_4_routing_0/rseg_4_v3_0.v19 GND 0.66926f
C356 rseg_4_routing_0/rseg_4_v3_0.v18 GND 0.73949f
C357 rseg_4_routing_0/rseg_4_v3_0.v7 GND 2.54397f
C358 rseg_4_routing_0/rseg_4_v3_0.v6 GND 0.84063f
C359 rseg_4_routing_0/rseg_4_v3_0.v5 GND 1.14719f
C360 rseg_4_routing_0/rseg_4_v3_0.v4 GND 0.77253f
C361 rseg_4_routing_0/rseg_4_v3_0.v3 GND 0.70326f
C362 rseg_4_routing_0/rseg_4_v3_0.v2 GND 0.72818f
C363 rseg_4_routing_0/rseg_4_v3_0.v61 GND 0.98585f
C364 rseg_4_routing_0/rseg_4_v3_0.v60 GND 1.48684f
C365 rseg_4_routing_0/rseg_4_v3_0.v59 GND 0.92749f
C366 rseg_4_routing_0/rseg_4_v3_0.v58 GND 2.26722f
C367 rseg_4_routing_0/rseg_4_v3_0.v57 GND 2.40805f
C368 rseg_4_routing_0/rseg_4_v3_0.v56 GND 3.42728f
C369 rseg_4_routing_0/rseg_4_v3_0.v46 GND 0.83546f
C370 rseg_4_routing_0/rseg_4_v3_0.v45 GND 0.83142f
C371 rseg_4_routing_0/rseg_4_v3_0.v44 GND 1.31433f
C372 rseg_4_routing_0/rseg_4_v3_0.v43 GND 0.8334f
C373 rseg_4_routing_0/rseg_4_v3_0.v42 GND 1.49005f
C374 rseg_4_routing_0/rseg_4_v3_0.v41 GND 2.32537f
C375 rseg_4_routing_0/rseg_4_v3_0.v40 GND 3.20861f
C376 rseg_4_routing_0/rseg_4_v3_0.v30 GND 0.79398f
C377 rseg_4_routing_0/rseg_4_v3_0.v29 GND 0.79447f
C378 rseg_4_routing_0/rseg_4_v3_0.v28 GND 1.27612f
C379 rseg_4_routing_0/rseg_4_v3_0.v27 GND 0.80491f
C380 rseg_4_routing_0/rseg_4_v3_0.v26 GND 1.44901f
C381 rseg_4_routing_0/rseg_4_v3_0.v25 GND 2.29648f
C382 rseg_4_routing_0/rseg_4_v3_0.v24 GND 3.14975f
C383 rseg_4_routing_0/rseg_4_v3_0.v14 GND 0.76536f
C384 rseg_4_routing_0/rseg_4_v3_0.v13 GND 0.79117f
C385 rseg_4_routing_0/rseg_4_v3_0.v12 GND 1.26691f
C386 rseg_4_routing_0/rseg_4_v3_0.v11 GND 0.79436f
C387 rseg_4_routing_0/rseg_4_v3_0.v10 GND 1.44302f
C388 rseg_4_routing_0/rseg_4_v3_0.v9 GND 2.29463f
C389 rseg_4_routing_0/rseg_4_v3_0.v8 GND 3.13866f
C390 rseg_4_routing_0/rseg_4_v3_0.v21.t1 GND 0.01292f
C391 rseg_4_routing_0/rseg_4_v3_0.v21.t2 GND 0.09788f
C392 rseg_4_routing_0/rseg_4_v3_0.v21.t0 GND 0.10105f
C393 rseg_4_routing_0/rseg_4_v3_0.v21.n0 GND 1.62825f
C394 a_34914_n5474.t2 GND 0.07342f
C395 a_34914_n5474.t1 GND 0.06664f
C396 a_34914_n5474.n0 GND 5.18539f
C397 a_34914_n5474.t0 GND 0.07455f
C398 rseg_4_routing_0/rseg_4_v3_0.v5.t0 GND 0.01294f
C399 rseg_4_routing_0/rseg_4_v3_0.v5.t2 GND 0.10145f
C400 rseg_4_routing_0/rseg_4_v3_0.v5.t1 GND 0.09797f
C401 rseg_4_routing_0/rseg_4_v3_0.v5.n0 GND 1.62712f
C402 a_36136_n5474.t2 GND 0.08054f
C403 a_36136_n5474.t1 GND 0.08241f
C404 a_36136_n5474.n0 GND 5.87337f
C405 a_36136_n5474.t0 GND 0.06369f
C406 rseg_4_routing_0/rseg_4_v3_0.v9.t0 GND 0.02752f
C407 rseg_4_routing_0/rseg_4_v3_0.v9.t1 GND 0.15141f
C408 rseg_4_routing_0/rseg_4_v3_0.v9.t2 GND 0.17047f
C409 rseg_4_routing_0/rseg_4_v3_0.v9.n0 GND 2.83038f
C410 rseg_4_routing_0/rseg_4_v3_0.v24.t1 GND 0.02265f
C411 rseg_4_routing_0/rseg_4_v3_0.v24.t2 GND 0.13251f
C412 rseg_4_routing_0/rseg_4_v3_0.v24.t0 GND 0.39728f
C413 rseg_4_routing_0/rseg_4_v3_0.v24.n0 GND 2.76757f
C414 a_29693_n8174.t1 GND 0.04948f
C415 a_29693_n8174.t4 GND 0.039f
C416 a_29693_n8174.n0 GND 2.59143f
C417 a_29693_n8174.t3 GND 0.05645f
C418 a_29693_n8174.n1 GND 2.38608f
C419 a_29693_n8174.t2 GND 0.039f
C420 a_29693_n8174.n2 GND 2.19006f
C421 a_29693_n8174.t0 GND 0.04849f
C422 rseg_4_routing_0/rseg_4_v3_0.v8.t0 GND 0.02279f
C423 rseg_4_routing_0/rseg_4_v3_0.v8.t1 GND 0.1333f
C424 rseg_4_routing_0/rseg_4_v3_0.v8.t2 GND 0.39585f
C425 rseg_4_routing_0/rseg_4_v3_0.v8.n0 GND 2.76319f
C426 rseg_4_routing_0/rseg_4_v3_0.v7.t0 GND 0.01248f
C427 rseg_4_routing_0/rseg_4_v3_0.v7.t1 GND 0.09062f
C428 rseg_4_routing_0/rseg_4_v3_0.v7.t2 GND 0.08856f
C429 rseg_4_routing_0/rseg_4_v3_0.v7.n0 GND 1.58095f
C430 a_31267_n6738.t1 GND 0.03957f
C431 a_31267_n6738.t3 GND 0.04498f
C432 a_31267_n6738.n0 GND 2.05844f
C433 a_31267_n6738.t4 GND 0.03831f
C434 a_31267_n6738.n1 GND 1.51138f
C435 a_31267_n6738.t2 GND 0.03831f
C436 a_31267_n6738.n2 GND 2.62168f
C437 a_31267_n6738.t0 GND 0.04733f
C438 a_35860_n5474.t2 GND 0.07897f
C439 a_35860_n5474.t1 GND 0.08079f
C440 a_35860_n5474.n0 GND 5.77629f
C441 a_35860_n5474.t0 GND 0.06395f
C442 rseg_4_routing_0/rseg_4_v3_0.v44.t1 GND 0.01506f
C443 rseg_4_routing_0/rseg_4_v3_0.v44.t2 GND 0.09069f
C444 rseg_4_routing_0/rseg_4_v3_0.v44.t0 GND 0.08797f
C445 rseg_4_routing_0/rseg_4_v3_0.v44.n0 GND 1.45497f
C446 rseg_4_routing_0/rseg_4_v3_0.v58.t1 GND 0.01583f
C447 rseg_4_routing_0/rseg_4_v3_0.v58.t2 GND 0.08108f
C448 rseg_4_routing_0/rseg_4_v3_0.v58.t0 GND 0.09013f
C449 rseg_4_routing_0/rseg_4_v3_0.v58.n0 GND 1.56677f
C450 a_32095_n6738.t1 GND 0.08006f
C451 a_32095_n6738.t3 GND 0.07704f
C452 a_32095_n6738.n0 GND 3.67426f
C453 a_32095_n6738.t4 GND 0.07394f
C454 a_32095_n6738.n1 GND 2.82116f
C455 a_32095_n6738.t2 GND 0.07394f
C456 a_32095_n6738.n2 GND 5.40641f
C457 a_32095_n6738.t0 GND 0.09319f
C458 a_35466_n5474.t2 GND 0.08071f
C459 a_35466_n5474.t1 GND 0.0698f
C460 a_35466_n5474.n0 GND 5.66782f
C461 a_35466_n5474.t0 GND 0.08167f
C462 rseg_4_routing_0/rseg_4_v3_0.v25.t2 GND 0.02742f
C463 rseg_4_routing_0/rseg_4_v3_0.v25.t1 GND 0.16899f
C464 rseg_4_routing_0/rseg_4_v3_0.v25.t0 GND 0.15083f
C465 rseg_4_routing_0/rseg_4_v3_0.v25.n0 GND 2.83612f
C466 rseg_4_routing_0/rseg_4_v3_0.v23.t1 GND 0.01247f
C467 rseg_4_routing_0/rseg_4_v3_0.v23.t2 GND 0.09059f
C468 rseg_4_routing_0/rseg_4_v3_0.v23.t0 GND 0.08855f
C469 rseg_4_routing_0/rseg_4_v3_0.v23.n0 GND 1.58122f
C470 a_31231_n8174.t1 GND 0.09555f
C471 a_31231_n8174.t4 GND 0.07299f
C472 a_31231_n8174.n0 GND 4.6643f
C473 a_31231_n8174.t3 GND 0.0965f
C474 a_31231_n8174.n1 GND 4.00369f
C475 a_31231_n8174.t2 GND 0.07299f
C476 a_31231_n8174.n2 GND 5.4004f
C477 a_31231_n8174.t0 GND 0.09358f
C478 a_35190_n5474.t2 GND 0.07488f
C479 a_35190_n5474.t1 GND 0.06634f
C480 a_35190_n5474.n0 GND 5.28272f
C481 a_35190_n5474.t0 GND 0.07606f
C482 rseg_4_routing_0/rseg_4_v3_0.v10.t0 GND 0.01438f
C483 rseg_4_routing_0/rseg_4_v3_0.v10.t2 GND 0.0778f
C484 rseg_4_routing_0/rseg_4_v3_0.v10.t1 GND 0.08736f
C485 rseg_4_routing_0/rseg_4_v3_0.v10.n0 GND 1.4371f
C486 a_31819_n6738.t1 GND 0.07983f
C487 a_31819_n6738.t3 GND 0.08121f
C488 a_31819_n6738.n0 GND 3.82467f
C489 a_31819_n6738.t4 GND 0.07505f
C490 a_31819_n6738.n1 GND 2.89621f
C491 a_31819_n6738.t2 GND 0.07505f
C492 a_31819_n6738.n2 GND 5.374f
C493 a_31819_n6738.t0 GND 0.09398f
C494 a_30245_n8174.t1 GND 0.0968f
C495 a_30245_n8174.t4 GND 0.07529f
C496 a_30245_n8174.n0 GND 5.41272f
C497 a_30245_n8174.t3 GND 0.1106f
C498 a_30245_n8174.n1 GND 4.73412f
C499 a_30245_n8174.t2 GND 0.07529f
C500 a_30245_n8174.n2 GND 4.30036f
C501 a_30245_n8174.t0 GND 0.09483f
C502 rseg_4_routing_0/rseg_4_v3_0.v12.t0 GND 0.01499f
C503 rseg_4_routing_0/rseg_4_v3_0.v12.t2 GND 0.09144f
C504 rseg_4_routing_0/rseg_4_v3_0.v12.t1 GND 0.08877f
C505 rseg_4_routing_0/rseg_4_v3_0.v12.n0 GND 1.46183f
C506 a_34638_n5474.t2 GND 0.03667f
C507 a_34638_n5474.t1 GND 0.0341f
C508 a_34638_n5474.n0 GND 2.59201f
C509 a_34638_n5474.t0 GND 0.03722f
C510 rseg_4_routing_0/rseg_4_v3_0.v28.t1 GND 0.01506f
C511 rseg_4_routing_0/rseg_4_v3_0.v28.t2 GND 0.08868f
C512 rseg_4_routing_0/rseg_4_v3_0.v28.t0 GND 0.09157f
C513 rseg_4_routing_0/rseg_4_v3_0.v28.n0 GND 1.45797f
C514 rseg_4_routing_0/rseg_4_v3_0.v53.t2 GND 0.01248f
C515 rseg_4_routing_0/rseg_4_v3_0.v53.t1 GND 0.09426f
C516 rseg_4_routing_0/rseg_4_v3_0.v53.t0 GND 0.09768f
C517 rseg_4_routing_0/rseg_4_v3_0.v53.n0 GND 1.54809f
C518 a_31507_n8174.t1 GND 0.09595f
C519 a_31507_n8174.t4 GND 0.07288f
C520 a_31507_n8174.n0 GND 4.84371f
C521 a_31507_n8174.t3 GND 0.09172f
C522 a_31507_n8174.n1 GND 3.72117f
C523 a_31507_n8174.t2 GND 0.07288f
C524 a_31507_n8174.n2 GND 5.40773f
C525 a_31507_n8174.t0 GND 0.09395f
C526 rseg_4_routing_0/rseg_4_v3_0.v26.t1 GND 0.01441f
C527 rseg_4_routing_0/rseg_4_v3_0.v26.t2 GND 0.07744f
C528 rseg_4_routing_0/rseg_4_v3_0.v26.t0 GND 0.08696f
C529 rseg_4_routing_0/rseg_4_v3_0.v26.n0 GND 1.43576f
C530 a_30521_n8174.t1 GND 0.08343f
C531 a_30521_n8174.t4 GND 0.06448f
C532 a_30521_n8174.n0 GND 4.80455f
C533 a_30521_n8174.t3 GND 0.0952f
C534 a_30521_n8174.n1 GND 4.09447f
C535 a_30521_n8174.t2 GND 0.06448f
C536 a_30521_n8174.n2 GND 3.71167f
C537 a_30521_n8174.t0 GND 0.08172f
C538 DEC0.t10 GND 0.06141f
C539 DEC0.t6 GND 0.06112f
C540 DEC0.n0 GND 0.19161f
C541 DEC0.t14 GND 0.06112f
C542 DEC0.n1 GND 0.09595f
C543 DEC0.t9 GND 0.06112f
C544 DEC0.n2 GND 0.07971f
C545 DEC0.t5 GND 0.06141f
C546 DEC0.t4 GND 0.06112f
C547 DEC0.n3 GND 0.19161f
C548 DEC0.t13 GND 0.06112f
C549 DEC0.n4 GND 0.09595f
C550 DEC0.t0 GND 0.06112f
C551 DEC0.n5 GND 0.07971f
C552 DEC0.n6 GND 0.09764f
C553 DEC0.t2 GND 0.06141f
C554 DEC0.t12 GND 0.06112f
C555 DEC0.n7 GND 0.19161f
C556 DEC0.t11 GND 0.06112f
C557 DEC0.n8 GND 0.09595f
C558 DEC0.t1 GND 0.06112f
C559 DEC0.n9 GND 0.09595f
C560 DEC0.t8 GND 0.06112f
C561 DEC0.n10 GND 0.09595f
C562 DEC0.t3 GND 0.06112f
C563 DEC0.n11 GND 0.09595f
C564 DEC0.t15 GND 0.06112f
C565 DEC0.n12 GND 0.09595f
C566 DEC0.t7 GND 0.06112f
C567 DEC0.n13 GND 0.21388f
C568 DEC0.n14 GND 0.29901f
C569 a_30955_n8174.t1 GND 0.08408f
C570 a_30955_n8174.t4 GND 0.0646f
C571 a_30955_n8174.n0 GND 3.95828f
C572 a_30955_n8174.t3 GND 0.08975f
C573 a_30955_n8174.n1 GND 3.79219f
C574 a_30955_n8174.t2 GND 0.0646f
C575 a_30955_n8174.n2 GND 4.76416f
C576 a_30955_n8174.t0 GND 0.08235f
C577 a_29969_n8174.t1 GND 0.09741f
C578 a_29969_n8174.t4 GND 0.07626f
C579 a_29969_n8174.n0 GND 5.27749f
C580 a_29969_n8174.t3 GND 0.11145f
C581 a_29969_n8174.n1 GND 4.74566f
C582 a_29969_n8174.t2 GND 0.07626f
C583 a_29969_n8174.n2 GND 4.32003f
C584 a_29969_n8174.t0 GND 0.09544f
C585 a_33357_n6738.t1 GND 0.04297f
C586 a_33357_n6738.t3 GND 0.0365f
C587 a_33357_n6738.n0 GND 2.11432f
C588 a_33357_n6738.t4 GND 0.03583f
C589 a_33357_n6738.n1 GND 1.26954f
C590 a_33357_n6738.t2 GND 0.03583f
C591 a_33357_n6738.n2 GND 2.81878f
C592 a_33357_n6738.t0 GND 0.04624f
C593 rseg_4_routing_0/rseg_4_v3_0.v37.t2 GND 0.01293f
C594 rseg_4_routing_0/rseg_4_v3_0.v37.t1 GND 0.09801f
C595 rseg_4_routing_0/rseg_4_v3_0.v37.t0 GND 0.10101f
C596 rseg_4_routing_0/rseg_4_v3_0.v37.n0 GND 1.62769f
C597 rseg_4_routing_0/rseg_4_v3_0.v42.t2 GND 0.01441f
C598 rseg_4_routing_0/rseg_4_v3_0.v42.t1 GND 0.07654f
C599 rseg_4_routing_0/rseg_4_v3_0.v42.t0 GND 0.0857f
C600 rseg_4_routing_0/rseg_4_v3_0.v42.n0 GND 1.43497f
C601 rseg_4_routing_0/rseg_4_v3_0.v56.t1 GND 0.0223f
C602 rseg_4_routing_0/rseg_4_v3_0.v56.t2 GND 0.12905f
C603 rseg_4_routing_0/rseg_4_v3_0.v56.t0 GND 0.42097f
C604 rseg_4_routing_0/rseg_4_v3_0.v56.n0 GND 2.85985f
C605 rseg_4_routing_0/rseg_4_v3_0.v55.t1 GND 0.01209f
C606 rseg_4_routing_0/rseg_4_v3_0.v55.t2 GND 0.08753f
C607 rseg_4_routing_0/rseg_4_v3_0.v55.t0 GND 0.08547f
C608 rseg_4_routing_0/rseg_4_v3_0.v55.n0 GND 1.50136f
C609 a_35584_n5474.t2 GND 0.0805f
C610 a_35584_n5474.t1 GND 0.08183f
C611 a_35584_n5474.n0 GND 5.8709f
C612 a_35584_n5474.t0 GND 0.06677f
C613 rseg_4_routing_0/rseg_4_v3_0.v41.t2 GND 0.02728f
C614 rseg_4_routing_0/rseg_4_v3_0.v41.t1 GND 0.16768f
C615 rseg_4_routing_0/rseg_4_v3_0.v41.t0 GND 0.1501f
C616 rseg_4_routing_0/rseg_4_v3_0.v41.n0 GND 2.84284f
C617 DEC2.t7 GND 0.06493f
C618 DEC2.t0 GND 0.06462f
C619 DEC2.n0 GND 0.20259f
C620 DEC2.t12 GND 0.06462f
C621 DEC2.n1 GND 0.10145f
C622 DEC2.t6 GND 0.06462f
C623 DEC2.n2 GND 0.10145f
C624 DEC2.t14 GND 0.06462f
C625 DEC2.n3 GND 0.10145f
C626 DEC2.t5 GND 0.06462f
C627 DEC2.n4 GND 0.10145f
C628 DEC2.t1 GND 0.06462f
C629 DEC2.n5 GND 0.16031f
C630 DEC2.t13 GND 0.0639f
C631 DEC2.n6 GND 0.08395f
C632 DEC2.t11 GND 0.06493f
C633 DEC2.t10 GND 0.06493f
C634 DEC2.t2 GND 0.06462f
C635 DEC2.n7 GND 0.20259f
C636 DEC2.t8 GND 0.06462f
C637 DEC2.n8 GND 0.10145f
C638 DEC2.t15 GND 0.06462f
C639 DEC2.n9 GND 0.10145f
C640 DEC2.t3 GND 0.06462f
C641 DEC2.n10 GND 0.10145f
C642 DEC2.t9 GND 0.06462f
C643 DEC2.n11 GND 0.10145f
C644 DEC2.n12 GND 0.16868f
C645 DEC2.t4 GND 0.0639f
C646 DEC2.n13 GND 0.16403f
C647 a_32805_n6738.t3 GND 0.08331f
C648 a_32805_n6738.t1 GND 0.07429f
C649 a_32805_n6738.n0 GND 3.92477f
C650 a_32805_n6738.t2 GND 0.09293f
C651 a_32805_n6738.t4 GND 0.07283f
C652 a_32805_n6738.n1 GND 5.53481f
C653 a_32805_n6738.n2 GND 2.64425f
C654 a_32805_n6738.t0 GND 0.07283f
C655 a_32529_n6738.t1 GND 0.0819f
C656 a_32529_n6738.t3 GND 0.07479f
C657 a_32529_n6738.n0 GND 3.75672f
C658 a_32529_n6738.t4 GND 0.09282f
C659 a_32529_n6738.t2 GND 0.07318f
C660 a_32529_n6738.n1 GND 5.4585f
C661 a_32529_n6738.n2 GND 2.6889f
C662 a_32529_n6738.t0 GND 0.07318f
C663 rseg_4_routing_0/rseg_4_v3_0.v60.t1 GND 0.01662f
C664 rseg_4_routing_0/rseg_4_v3_0.v60.t2 GND 0.09404f
C665 rseg_4_routing_0/rseg_4_v3_0.v60.t0 GND 0.09697f
C666 rseg_4_routing_0/rseg_4_v3_0.v60.n0 GND 1.57947f
C667 rseg_4_routing_0/rseg_4_v3_0.v57.t2 GND 0.02716f
C668 rseg_4_routing_0/rseg_4_v3_0.v57.t1 GND 0.1492f
C669 rseg_4_routing_0/rseg_4_v3_0.v57.t0 GND 0.16449f
C670 rseg_4_routing_0/rseg_4_v3_0.v57.n0 GND 2.95161f
C671 a_31543_n6738.t3 GND 0.07971f
C672 a_31543_n6738.t2 GND 0.0947f
C673 a_31543_n6738.t4 GND 0.07612f
C674 a_31543_n6738.n0 GND 5.33217f
C675 a_31543_n6738.t1 GND 0.07612f
C676 a_31543_n6738.n1 GND 2.97065f
C677 a_31543_n6738.n2 GND 3.98477f
C678 a_31543_n6738.t0 GND 0.08576f
C679 DEC3.t3 GND 0.06266f
C680 DEC3.t2 GND 0.06236f
C681 DEC3.n0 GND 0.19549f
C682 DEC3.t8 GND 0.06236f
C683 DEC3.n1 GND 0.09789f
C684 DEC3.t1 GND 0.06236f
C685 DEC3.n2 GND 0.09789f
C686 DEC3.t12 GND 0.06236f
C687 DEC3.n3 GND 0.09789f
C688 DEC3.t6 GND 0.06236f
C689 DEC3.n4 GND 0.09789f
C690 DEC3.t0 GND 0.06236f
C691 DEC3.n5 GND 0.09789f
C692 DEC3.t9 GND 0.06236f
C693 DEC3.n6 GND 0.25521f
C694 DEC3.t15 GND 0.06266f
C695 DEC3.t11 GND 0.06236f
C696 DEC3.n7 GND 0.19549f
C697 DEC3.t5 GND 0.06236f
C698 DEC3.n8 GND 0.09789f
C699 DEC3.t14 GND 0.06236f
C700 DEC3.n9 GND 0.08132f
C701 DEC3.t13 GND 0.06266f
C702 DEC3.t7 GND 0.06236f
C703 DEC3.n10 GND 0.19549f
C704 DEC3.t10 GND 0.06236f
C705 DEC3.n11 GND 0.09789f
C706 DEC3.t4 GND 0.06236f
C707 DEC3.n12 GND 0.08132f
C708 DEC3.n13 GND 0.07851f
C709 a_33081_n6738.t4 GND 0.08487f
C710 a_33081_n6738.t1 GND 0.07389f
C711 a_33081_n6738.n0 GND 4.0948f
C712 a_33081_n6738.t2 GND 0.09304f
C713 a_33081_n6738.t3 GND 0.07249f
C714 a_33081_n6738.n1 GND 5.60801f
C715 a_33081_n6738.n2 GND 2.60041f
C716 a_33081_n6738.t0 GND 0.07249f
C717 DEC1.t8 GND 0.06373f
C718 DEC1.t0 GND 0.06342f
C719 DEC1.n0 GND 0.19883f
C720 DEC1.t1 GND 0.06342f
C721 DEC1.n1 GND 0.09957f
C722 DEC1.t7 GND 0.06342f
C723 DEC1.n2 GND 0.09957f
C724 DEC1.t15 GND 0.06342f
C725 DEC1.n3 GND 0.09957f
C726 DEC1.t9 GND 0.06342f
C727 DEC1.n4 GND 0.09957f
C728 DEC1.t6 GND 0.06342f
C729 DEC1.n5 GND 0.15733f
C730 DEC1.t14 GND 0.06272f
C731 DEC1.n6 GND 0.08681f
C732 DEC1.t5 GND 0.06373f
C733 DEC1.t11 GND 0.06392f
C734 DEC1.t2 GND 0.0636f
C735 DEC1.n7 GND 0.21516f
C736 DEC1.t3 GND 0.0636f
C737 DEC1.n8 GND 0.10774f
C738 DEC1.t12 GND 0.0636f
C739 DEC1.n9 GND 0.10774f
C740 DEC1.t4 GND 0.0636f
C741 DEC1.n10 GND 0.10774f
C742 DEC1.t10 GND 0.0636f
C743 DEC1.n11 GND 0.10774f
C744 DEC1.n12 GND 0.16555f
C745 DEC1.t13 GND 0.06272f
C746 DEC1.n13 GND 0.16147f
C747 VPB.n0 GND 0.01416f
C748 VPB.n1 GND 0.01402f
C749 VPB.n2 GND 0.02309f
C750 VPB.n3 GND 0.09183f
C751 VPB.n4 GND 0.09183f
C752 VPB.t21 GND 0.07936f
C753 VPB.t91 GND 0.0814f
C754 VPB.t7 GND 0.0814f
C755 VPB.t47 GND 0.06105f
C756 VPB.n7 GND 0.01783f
C757 VPB.n8 GND 0.09183f
C758 VPB.n9 GND 0.09183f
C759 VPB.t51 GND 0.07936f
C760 VPB.t89 GND 0.0814f
C761 VPB.t78 GND 0.0814f
C762 VPB.t42 GND 0.06105f
C763 VPB.t2 GND 0.07936f
C764 VPB.t35 GND 0.0814f
C765 VPB.t13 GND 0.0814f
C766 VPB.t4 GND 0.06105f
C767 VPB.n10 GND 0.01724f
C768 VPB.n12 GND 0.02506f
C769 VPB.n13 GND 0.09183f
C770 VPB.n14 GND 0.09183f
C771 VPB.t12 GND 0.07936f
C772 VPB.t52 GND 0.0814f
C773 VPB.t46 GND 0.0814f
C774 VPB.t81 GND 0.06105f
C775 VPB.t11 GND 0.07936f
C776 VPB.t61 GND 0.0814f
C777 VPB.t48 GND 0.0814f
C778 VPB.t40 GND 0.06105f
C779 VPB.n15 GND 0.01701f
C780 VPB.n16 GND 0.03845f
C781 VPB.n17 GND 0.03845f
C782 VPB.n18 GND 0.01863f
C783 VPB.n19 GND 0.01212f
C784 VPB.n20 GND 0.01724f
C785 VPB.n21 GND 0.01724f
C786 VPB.n23 GND 0.02691f
C787 VPB.n24 GND 0.09183f
C788 VPB.n25 GND 0.09183f
C789 VPB.t36 GND 0.07936f
C790 VPB.t0 GND 0.0814f
C791 VPB.t19 GND 0.0814f
C792 VPB.t50 GND 0.06105f
C793 VPB.t16 GND 0.07936f
C794 VPB.t34 GND 0.0814f
C795 VPB.t37 GND 0.0814f
C796 VPB.t92 GND 0.06105f
C797 VPB.n26 GND 0.01701f
C798 VPB.n28 GND 0.03795f
C799 VPB.n29 GND 0.01888f
C800 VPB.n30 GND 0.09183f
C801 VPB.n31 GND 0.09183f
C802 VPB.t77 GND 0.07936f
C803 VPB.t74 GND 0.0814f
C804 VPB.t73 GND 0.0814f
C805 VPB.t70 GND 0.06105f
C806 VPB.t76 GND 0.07936f
C807 VPB.t71 GND 0.0814f
C808 VPB.t72 GND 0.0814f
C809 VPB.t75 GND 0.06105f
C810 VPB.n32 GND 0.03066f
C811 VPB.n33 GND 0.02055f
C812 VPB.n34 GND 0.01948f
C813 VPB.n35 GND 0.03845f
C814 VPB.n36 GND 0.03845f
C815 VPB.n37 GND 0.01579f
C816 VPB.n38 GND 0.01862f
C817 VPB.n39 GND 0.01724f
C818 VPB.n40 GND 0.09183f
C819 VPB.n41 GND 0.09183f
C820 VPB.t30 GND 0.07936f
C821 VPB.t31 GND 0.0814f
C822 VPB.t65 GND 0.0814f
C823 VPB.t57 GND 0.06105f
C824 VPB.n43 GND 0.01512f
C825 VPB.n44 GND 0.01494f
C826 VPB.n46 GND 0.01783f
C827 VPB.n47 GND 0.09183f
C828 VPB.n49 GND 0.01431f
C829 VPB.n50 GND 0.01483f
C830 VPB.n52 GND 0.09183f
C831 VPB.t69 GND 0.07936f
C832 VPB.t93 GND 0.0814f
C833 VPB.t49 GND 0.0814f
C834 VPB.t17 GND 0.06105f
C835 VPB.t20 GND 0.07936f
C836 VPB.t38 GND 0.0814f
C837 VPB.t26 GND 0.0814f
C838 VPB.t25 GND 0.06105f
C839 VPB.n54 GND 0.03845f
C840 VPB.n55 GND 0.0407f
C841 VPB.n56 GND 0.03845f
C842 VPB.n57 GND 0.01945f
C843 VPB.n58 GND 0.01875f
C844 VPB.n59 GND 0.01875f
C845 VPB.n60 GND 0.02107f
C846 VPB.n61 GND 0.03845f
C847 VPB.t14 GND 0.07936f
C848 VPB.t5 GND 0.0814f
C849 VPB.t87 GND 0.0814f
C850 VPB.t32 GND 0.06105f
C851 VPB.n62 GND 0.0407f
C852 VPB.n63 GND 0.03845f
C853 VPB.n65 GND 0.01889f
C854 VPB.n66 GND 0.02691f
C855 VPB.n67 GND 0.03845f
C856 VPB.n68 GND 0.03845f
C857 VPB.n69 GND 0.02107f
C858 VPB.n70 GND 0.02309f
C859 VPB.n71 GND 0.09183f
C860 VPB.t62 GND 0.07936f
C861 VPB.t88 GND 0.0814f
C862 VPB.t58 GND 0.0814f
C863 VPB.t44 GND 0.06105f
C864 VPB.n72 GND 0.0407f
C865 VPB.t64 GND 0.06105f
C866 VPB.t15 GND 0.0814f
C867 VPB.t59 GND 0.0814f
C868 VPB.t43 GND 0.07936f
C869 VPB.n73 GND 0.09183f
C870 VPB.n76 GND 0.01575f
C871 VPB.n77 GND 0.01494f
C872 VPB.n78 GND 0.01701f
C873 VPB.n79 GND 0.01945f
C874 VPB.n80 GND 0.01888f
C875 VPB.n81 GND 0.01313f
C876 VPB.n82 GND 0.09183f
C877 VPB.t6 GND 0.07936f
C878 VPB.t33 GND 0.0814f
C879 VPB.t45 GND 0.0814f
C880 VPB.t79 GND 0.06105f
C881 VPB.n83 GND 0.0407f
C882 VPB.t60 GND 0.06105f
C883 VPB.t18 GND 0.0814f
C884 VPB.t1 GND 0.0814f
C885 VPB.t86 GND 0.07936f
C886 VPB.n84 GND 0.09183f
C887 VPB.n86 GND 0.02253f
C888 VPB.n87 GND 0.01491f
C889 VPB.n88 GND 0.02418f
C890 VPB.n89 GND 0.11718f
C891 VPB.n90 GND 0.11718f
C892 VPB.t53 GND 0.07936f
C893 VPB.t22 GND 0.0814f
C894 VPB.t82 GND 0.0814f
C895 VPB.t23 GND 0.08553f
C896 VPB.t84 GND 0.08553f
C897 VPB.t10 GND 0.0814f
C898 VPB.t9 GND 0.06724f
C899 VPB.t24 GND 0.08349f
C900 VPB.t83 GND 0.08966f
C901 VPB.t28 GND 0.08553f
C902 VPB.t8 GND 0.08553f
C903 VPB.t66 GND 0.08553f
C904 VPB.t67 GND 0.08553f
C905 VPB.t54 GND 0.05899f
C906 VPB.n91 GND 0.02055f
C907 VPB.n92 GND 0.03747f
C908 VPB.n93 GND 0.06363f
C909 VPB.n94 GND 0.0407f
C910 VPB.n95 GND 0.06363f
C911 VPB.n96 GND 0.03426f
C912 VPB.n97 GND 0.02418f
C913 VPB.n99 GND 0.01655f
C914 VPB.n100 GND 0.01331f
C915 VPB.n101 GND 0.03845f
C916 VPB.n102 GND 0.0407f
C917 VPB.n103 GND 0.03845f
C918 VPB.n104 GND 0.01945f
C919 VPB.n105 GND 0.03795f
C920 VPB.n106 GND 0.0141f
C921 VPB.n107 GND 0.0173f
C922 VPB.n108 GND 0.01336f
C923 VPB.n109 GND 0.03845f
C924 VPB.n110 GND 0.0407f
C925 VPB.n111 GND 0.03845f
C926 VPB.n112 GND 0.01945f
C927 VPB.n113 GND 0.02564f
C928 VPB.n114 GND 0.01945f
C929 VPB.n115 GND 0.02564f
C930 VPB.n117 GND 0.09183f
C931 VPB.t63 GND 0.07936f
C932 VPB.t85 GND 0.0814f
C933 VPB.t68 GND 0.0814f
C934 VPB.t29 GND 0.06105f
C935 VPB.n118 GND 0.0407f
C936 VPB.t41 GND 0.06105f
C937 VPB.t90 GND 0.0814f
C938 VPB.t56 GND 0.0814f
C939 VPB.t39 GND 0.07936f
C940 VPB.n119 GND 0.09183f
C941 VPB.n122 GND 0.01754f
C942 VPB.n123 GND 0.01313f
C943 VPB.n124 GND 0.02107f
C944 VPB.n125 GND 0.03845f
C945 VPB.n126 GND 0.0407f
C946 VPB.n127 GND 0.03845f
C947 VPB.n128 GND 0.01945f
C948 VPB.n129 GND 0.02506f
C949 VPB.n130 GND 0.01456f
C950 VPB.n131 GND 0.01724f
C951 VPB.n133 GND 0.03845f
C952 VPB.n134 GND 0.0407f
C953 VPB.n135 GND 0.03845f
C954 VPB.n136 GND 0.01945f
C955 VPB.n137 GND 0.01728f
C956 VPB.n138 GND 0.01728f
C957 VPB.n139 GND 0.02107f
C958 VPB.n140 GND 0.03845f
C959 VPB.t3 GND 0.07936f
C960 VPB.t55 GND 0.0814f
C961 VPB.t80 GND 0.0814f
C962 VPB.t27 GND 0.06105f
C963 VPB.n141 GND 0.0407f
C964 VPB.n142 GND 0.03845f
C965 VPB.n143 GND 0.0146f
C966 VPB.n144 GND 0.01467f
C967 a_31783_n8174.t1 GND 0.04927f
C968 a_31783_n8174.t3 GND 0.03722f
C969 a_31783_n8174.n0 GND 2.56635f
C970 a_31783_n8174.t4 GND 0.04443f
C971 a_31783_n8174.n1 GND 1.74851f
C972 a_31783_n8174.t2 GND 0.03722f
C973 a_31783_n8174.n2 GND 2.76876f
C974 a_31783_n8174.t0 GND 0.04824f
C975 a_36412_n5474.t2 GND 0.04203f
C976 a_36412_n5474.t1 GND 0.03172f
C977 a_36412_n5474.n0 GND 2.9852f
C978 a_36412_n5474.t0 GND 0.04106f
C979 rseg_4_routing_0/rseg_4_v3_0.v40.t0 GND 0.02245f
C980 rseg_4_routing_0/rseg_4_v3_0.v40.t2 GND 0.13085f
C981 rseg_4_routing_0/rseg_4_v3_0.v40.t1 GND 0.40073f
C982 rseg_4_routing_0/rseg_4_v3_0.v40.n0 GND 2.77279f
C983 rseg_4_routing_0/rseg_4_v3_0.v39.t1 GND 0.0125f
C984 rseg_4_routing_0/rseg_4_v3_0.v39.t2 GND 0.0907f
C985 rseg_4_routing_0/rseg_4_v3_0.v39.t0 GND 0.08878f
C986 rseg_4_routing_0/rseg_4_v3_0.v39.n0 GND 1.58019f
.ends

