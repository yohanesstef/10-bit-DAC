magic
tech sky130A
magscale 1 2
timestamp 1751042016
<< error_p >>
rect -223 321 223 355
rect -253 106 253 321
rect -223 72 223 106
rect -253 -143 253 72
rect -253 -389 -223 -177
rect -187 -323 -157 -243
rect 157 -323 187 -243
rect -187 -327 187 -323
rect 223 -389 253 -177
rect -253 -393 253 -389
<< nwell >>
rect -223 109 223 355
rect -223 -140 223 106
rect -223 -389 223 -143
<< mvpmos >>
rect -129 171 -29 255
rect 29 171 129 255
rect -129 -78 -29 6
rect 29 -78 129 6
rect -129 -327 -29 -243
rect 29 -327 129 -243
<< mvpdiff >>
rect -187 243 -129 255
rect -187 183 -175 243
rect -141 183 -129 243
rect -187 171 -129 183
rect -29 243 29 255
rect -29 183 -17 243
rect 17 183 29 243
rect -29 171 29 183
rect 129 243 187 255
rect 129 183 141 243
rect 175 183 187 243
rect 129 171 187 183
rect -187 -6 -129 6
rect -187 -66 -175 -6
rect -141 -66 -129 -6
rect -187 -78 -129 -66
rect -29 -6 29 6
rect -29 -66 -17 -6
rect 17 -66 29 -6
rect -29 -78 29 -66
rect 129 -6 187 6
rect 129 -66 141 -6
rect 175 -66 187 -6
rect 129 -78 187 -66
rect -187 -255 -129 -243
rect -187 -315 -175 -255
rect -141 -315 -129 -255
rect -187 -327 -129 -315
rect -29 -255 29 -243
rect -29 -315 -17 -255
rect 17 -315 29 -255
rect -29 -327 29 -315
rect 129 -255 187 -243
rect 129 -315 141 -255
rect 175 -315 187 -255
rect 129 -327 187 -315
<< mvpdiffc >>
rect -175 183 -141 243
rect -17 183 17 243
rect 141 183 175 243
rect -175 -66 -141 -6
rect -17 -66 17 -6
rect 141 -66 175 -6
rect -175 -315 -141 -255
rect -17 -315 17 -255
rect 141 -315 175 -255
<< poly >>
rect -129 336 -29 352
rect -129 302 -113 336
rect -45 302 -29 336
rect -129 255 -29 302
rect 29 336 129 352
rect 29 302 45 336
rect 113 302 129 336
rect 29 255 129 302
rect -129 145 -29 171
rect 29 145 129 171
rect -129 87 -29 103
rect -129 53 -113 87
rect -45 53 -29 87
rect -129 6 -29 53
rect 29 87 129 103
rect 29 53 45 87
rect 113 53 129 87
rect 29 6 129 53
rect -129 -104 -29 -78
rect 29 -104 129 -78
rect -129 -162 -29 -146
rect -129 -196 -113 -162
rect -45 -196 -29 -162
rect -129 -243 -29 -196
rect 29 -162 129 -146
rect 29 -196 45 -162
rect 113 -196 129 -162
rect 29 -243 129 -196
rect -129 -353 -29 -327
rect 29 -353 129 -327
<< polycont >>
rect -113 302 -45 336
rect 45 302 113 336
rect -113 53 -45 87
rect 45 53 113 87
rect -113 -196 -45 -162
rect 45 -196 113 -162
<< locali >>
rect -129 302 -113 336
rect -45 302 -29 336
rect 29 302 45 336
rect 113 302 129 336
rect -175 243 -141 259
rect -175 167 -141 183
rect -17 243 17 259
rect -17 167 17 183
rect 141 243 175 259
rect 141 167 175 183
rect -129 53 -113 87
rect -45 53 -29 87
rect 29 53 45 87
rect 113 53 129 87
rect -175 -6 -141 10
rect -175 -82 -141 -66
rect -17 -6 17 10
rect -17 -82 17 -66
rect 141 -6 175 10
rect 141 -82 175 -66
rect -129 -196 -113 -162
rect -45 -196 -29 -162
rect 29 -196 45 -162
rect 113 -196 129 -162
rect -175 -255 -141 -239
rect -175 -331 -141 -315
rect -17 -255 17 -239
rect -17 -331 17 -315
rect 141 -255 175 -239
rect 141 -331 175 -315
<< viali >>
rect -105 302 -53 336
rect 53 302 105 336
rect -175 183 -141 243
rect -17 183 17 243
rect 141 183 175 243
rect -105 53 -53 87
rect 53 53 105 87
rect -175 -66 -141 -6
rect -17 -66 17 -6
rect 141 -66 175 -6
rect -105 -196 -53 -162
rect 53 -196 105 -162
rect -175 -315 -141 -255
rect -17 -315 17 -255
rect 141 -315 175 -255
<< metal1 >>
rect -117 336 -41 342
rect -117 302 -105 336
rect -53 302 -41 336
rect -117 296 -41 302
rect 41 336 117 342
rect 41 302 53 336
rect 105 302 117 336
rect 41 296 117 302
rect -181 243 -135 255
rect -181 183 -175 243
rect -141 183 -135 243
rect -181 171 -135 183
rect -23 243 23 255
rect -23 183 -17 243
rect 17 183 23 243
rect -23 171 23 183
rect 135 243 181 255
rect 135 183 141 243
rect 175 183 181 243
rect 135 171 181 183
rect -117 87 -41 93
rect -117 53 -105 87
rect -53 53 -41 87
rect -117 47 -41 53
rect 41 87 117 93
rect 41 53 53 87
rect 105 53 117 87
rect 41 47 117 53
rect -181 -6 -135 6
rect -181 -66 -175 -6
rect -141 -66 -135 -6
rect -181 -78 -135 -66
rect -23 -6 23 6
rect -23 -66 -17 -6
rect 17 -66 23 -6
rect -23 -78 23 -66
rect 135 -6 181 6
rect 135 -66 141 -6
rect 175 -66 181 -6
rect 135 -78 181 -66
rect -117 -162 -41 -156
rect -117 -196 -105 -162
rect -53 -196 -41 -162
rect -117 -202 -41 -196
rect 41 -162 117 -156
rect 41 -196 53 -162
rect 105 -196 117 -162
rect 41 -202 117 -196
rect -181 -255 -135 -243
rect -181 -315 -175 -255
rect -141 -315 -135 -255
rect -181 -327 -135 -315
rect -23 -255 23 -243
rect -23 -315 -17 -255
rect 17 -315 23 -255
rect -23 -327 23 -315
rect 135 -255 181 -243
rect 135 -315 141 -255
rect 175 -315 181 -255
rect 135 -327 181 -315
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 0.50 m 3 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
