magic
tech sky130A
magscale 1 2
timestamp 1749654170
<< nwell >>
rect -601 499 955 1949
<< mvnsubdiff >>
rect -535 1870 889 1883
rect -535 1836 -475 1870
rect 829 1836 889 1870
rect -535 1823 889 1836
rect -535 612 889 625
rect -535 578 -475 612
rect 829 578 889 612
rect -535 565 889 578
<< mvnsubdiffcont >>
rect -475 1836 829 1870
rect -475 578 829 612
<< locali >>
rect -535 1836 -475 1870
rect 829 1836 889 1870
rect -535 578 -475 612
rect 829 578 889 612
<< viali >>
rect -475 1836 829 1870
rect -377 1723 -233 1757
rect -35 1723 109 1757
rect 307 1723 451 1757
rect 649 1723 793 1757
<< metal1 >>
rect -535 1870 889 1883
rect -535 1836 -475 1870
rect 829 1836 889 1870
rect -535 1823 889 1836
rect -389 1757 -221 1823
rect -389 1723 -377 1757
rect -233 1723 -221 1757
rect -389 1711 -221 1723
rect -47 1757 121 1823
rect -47 1723 -35 1757
rect 109 1723 121 1757
rect -47 1711 121 1723
rect 295 1757 463 1823
rect 295 1723 307 1757
rect 451 1723 463 1757
rect 295 1711 463 1723
rect 637 1757 805 1823
rect 637 1723 649 1757
rect 793 1723 805 1757
rect 637 1711 805 1723
rect -535 1581 889 1641
rect -229 1427 -169 1452
rect -483 1339 -423 1345
rect -483 1273 -423 1279
rect -483 1081 -417 1087
rect -483 1015 -417 1021
rect -483 823 -417 829
rect -483 757 -417 763
rect -229 731 -169 1367
rect -141 1427 -81 1433
rect -141 1361 -81 1367
rect 113 1339 173 1438
rect 201 1427 261 1433
rect 201 1361 261 1367
rect 113 1169 173 1279
rect -141 1081 -75 1087
rect -141 1015 -75 1021
rect -141 823 -75 829
rect -141 757 -75 763
rect 113 731 173 1109
rect 201 1169 261 1175
rect 201 1103 261 1109
rect 455 1081 515 1438
rect 543 1427 603 1433
rect 543 1361 603 1367
rect 543 1169 603 1175
rect 543 1103 603 1109
rect 455 911 515 1021
rect 455 851 603 911
rect 201 823 267 829
rect 201 757 267 763
rect 455 731 515 851
rect 797 823 857 1438
rect 797 731 857 763
rect -257 685 -169 731
rect 85 685 173 731
rect 427 685 515 731
rect 769 685 857 731
<< via1 >>
rect -229 1367 -169 1427
rect -483 1279 -423 1339
rect -483 1021 -417 1081
rect -483 763 -417 823
rect -141 1367 -81 1427
rect 201 1367 261 1427
rect 113 1279 173 1339
rect 113 1109 173 1169
rect -141 1021 -75 1081
rect -141 763 -75 823
rect 201 1109 261 1169
rect 543 1367 603 1427
rect 543 1109 603 1169
rect 455 1021 515 1081
rect 201 763 267 823
rect 797 763 857 823
<< metal2 >>
rect -235 1367 -229 1427
rect -169 1367 -141 1427
rect -81 1367 201 1427
rect 261 1367 543 1427
rect 603 1367 609 1427
rect -489 1279 -483 1339
rect -423 1279 113 1339
rect 173 1279 179 1339
rect 107 1109 113 1169
rect 173 1109 201 1169
rect 261 1109 543 1169
rect 603 1109 609 1169
rect -489 1021 -483 1081
rect -417 1021 -141 1081
rect -75 1021 455 1081
rect 515 1021 521 1081
rect -489 763 -483 823
rect -417 763 -141 823
rect -75 763 201 823
rect 267 763 797 823
rect 857 763 863 823
use sky130_fd_pr__pfet_g5v0d10v5_4VG7B4  sky130_fd_pr__pfet_g5v0d10v5_4VG7B4_0
timestamp 1749638674
transform 0 -1 1 1 0 1224
box -611 -186 611 148
use sky130_fd_pr__pfet_g5v0d10v5_4VG7B4  sky130_fd_pr__pfet_g5v0d10v5_4VG7B4_1
timestamp 1749638674
transform 0 -1 685 1 0 1224
box -611 -186 611 148
use sky130_fd_pr__pfet_g5v0d10v5_4VG7B4  sky130_fd_pr__pfet_g5v0d10v5_4VG7B4_2
timestamp 1749638674
transform 0 -1 343 1 0 1224
box -611 -186 611 148
use sky130_fd_pr__pfet_g5v0d10v5_4VG7B4  XM1
timestamp 1749638674
transform 0 -1 -341 1 0 1224
box -611 -186 611 148
<< end >>
