magic
tech sky130A
magscale 1 2
timestamp 1750900893
<< locali >>
rect 5620 4517 5654 6150
rect 10462 4517 10496 6150
rect 11374 4517 11408 6150
rect 13698 4517 13732 6116
rect 1885 3585 1919 4075
rect 4365 3585 4399 4075
rect 6675 3585 6709 4075
rect 9198 3585 9232 4075
rect 11565 3585 11599 4075
rect 14049 3585 14083 4075
<< metal1 >>
rect 906 4195 966 4307
rect -535 4135 966 4195
rect -535 3243 -475 4135
rect 1182 4107 1242 4307
rect -447 4047 1242 4107
rect -447 3243 -387 4047
rect 1458 4019 1518 4307
rect -359 3959 1518 4019
rect -359 3243 -299 3959
rect 1734 3931 1794 4307
rect -271 3871 1794 3931
rect -271 3243 -211 3871
rect 2010 3843 2070 4307
rect 2286 3931 2346 4307
rect 2562 4019 2622 4307
rect 2838 4107 2898 4307
rect 3114 4195 3174 4307
rect 3390 4195 3450 4307
rect 3114 4135 3215 4195
rect 2838 4047 3127 4107
rect 2562 3959 3039 4019
rect 2286 3871 2951 3931
rect 2010 3783 2863 3843
rect 2803 3243 2863 3783
rect 2891 3243 2951 3871
rect 2979 3243 3039 3959
rect 3067 3243 3127 4047
rect 3155 3244 3215 4135
rect 3243 4135 3450 4195
rect 3243 3244 3303 4135
rect 3666 4107 3726 4307
rect 3331 4047 3726 4107
rect 3331 3244 3391 4047
rect 3942 4019 4002 4307
rect 3419 3959 4002 4019
rect 3419 3244 3479 3959
rect 4218 3931 4278 4307
rect 3507 3871 4278 3931
rect 4494 3931 4554 4307
rect 4770 4019 4830 4307
rect 5046 4107 5106 4307
rect 5322 4195 5382 4307
rect 5748 4195 5808 4307
rect 5322 4135 5640 4195
rect 5046 4047 5552 4107
rect 4770 3959 5464 4019
rect 4494 3871 5376 3931
rect 3507 3244 3567 3871
rect 5316 3243 5376 3871
rect 5404 3243 5464 3959
rect 5492 3243 5552 4047
rect 5580 3243 5640 4135
rect 5668 4135 5808 4195
rect 5668 3243 5728 4135
rect 6024 4107 6084 4307
rect 5756 4047 6084 4107
rect 5756 3243 5816 4047
rect 6300 4019 6360 4307
rect 5844 3959 6360 4019
rect 5844 3243 5904 3959
rect 6576 3931 6636 4307
rect 5932 3871 6636 3931
rect 5932 3243 5992 3871
rect 6852 3843 6912 4307
rect 7128 3931 7188 4307
rect 7404 4019 7464 4307
rect 7680 4107 7740 4307
rect 7956 4195 8016 4307
rect 8232 4195 8292 4307
rect 7956 4135 8128 4195
rect 7680 4047 8040 4107
rect 7404 3959 7952 4019
rect 7128 3871 7864 3931
rect 6852 3783 7776 3843
rect 7716 3243 7776 3783
rect 7804 3243 7864 3871
rect 7892 3243 7952 3959
rect 7980 3243 8040 4047
rect 8068 3244 8128 4135
rect 8156 4135 8292 4195
rect 8156 3244 8216 4135
rect 8508 4107 8568 4307
rect 8244 4047 8568 4107
rect 8244 3244 8304 4047
rect 8784 4019 8844 4307
rect 8332 3959 8844 4019
rect 8332 3244 8392 3959
rect 9060 3931 9120 4307
rect 8420 3871 9120 3931
rect 9336 3931 9396 4307
rect 9612 4019 9672 4307
rect 9888 4107 9948 4307
rect 10164 4195 10224 4307
rect 10590 4195 10650 4307
rect 10164 4135 10446 4195
rect 9888 4047 10358 4107
rect 9612 3959 10270 4019
rect 9336 3871 10182 3931
rect 8420 3244 8480 3871
rect 10122 3243 10182 3871
rect 10210 3243 10270 3959
rect 10298 3243 10358 4047
rect 10386 3243 10446 4135
rect 10477 4135 10650 4195
rect 10477 3243 10537 4135
rect 10866 4107 10926 4307
rect 10565 4047 10926 4107
rect 10565 3243 10625 4047
rect 11142 4019 11202 4307
rect 10653 3959 11202 4019
rect 10653 3243 10713 3959
rect 11418 3931 11478 4307
rect 10741 3871 11478 3931
rect 10741 3243 10801 3871
rect 11694 3843 11754 4307
rect 11970 3931 12030 4307
rect 12246 4019 12306 4307
rect 12522 4107 12582 4307
rect 12798 4195 12858 4307
rect 13074 4195 13134 4307
rect 12798 4135 12865 4195
rect 12522 4047 12777 4107
rect 12246 3959 12689 4019
rect 11970 3871 12601 3931
rect 11694 3783 12513 3843
rect 12453 3243 12513 3783
rect 12541 3243 12601 3871
rect 12629 3243 12689 3959
rect 12717 3243 12777 4047
rect 12805 3244 12865 4135
rect 12894 4135 13134 4195
rect 12894 3244 12954 4135
rect 13350 4107 13410 4307
rect 12982 4047 13410 4107
rect 12982 3244 13042 4047
rect 13626 4019 13686 4307
rect 13070 3959 13686 4019
rect 13070 3244 13130 3959
rect 13902 3931 13962 4307
rect 13158 3871 13962 3931
rect 14178 3931 14238 4307
rect 14454 4019 14514 4307
rect 14730 4107 14790 4307
rect 15006 4195 15066 4307
rect 15006 4135 15512 4195
rect 14730 4047 15424 4107
rect 14454 3959 15336 4019
rect 14178 3871 15248 3931
rect 13158 3244 13218 3871
rect 15188 3243 15248 3871
rect 15276 3243 15336 3959
rect 15364 3243 15424 4047
rect 15452 3243 15512 4135
<< metal2 >>
rect 11318 6985 13562 7045
rect 11042 6897 13286 6957
rect 10766 6809 12706 6869
rect 10490 6721 12126 6781
rect 10214 6633 11546 6693
rect 4664 6000 14420 6060
rect 4388 5912 14144 5972
rect 4940 5824 14696 5884
rect 4112 5736 13868 5796
rect 5216 5648 14972 5708
rect 3836 5560 13592 5620
rect 5492 5472 15248 5532
rect 3560 5384 13316 5444
rect 3284 5296 13040 5356
rect 1076 5208 10832 5268
rect 3008 5120 12764 5180
rect 1352 5032 11108 5092
rect 2732 4944 12488 5004
rect 1628 4856 11384 4916
rect 2456 4768 12212 4828
rect 1904 4680 11660 4740
rect 2180 4592 11936 4652
use rseg_2_v3  rseg_2_v3_0
timestamp 1749563245
transform 1 0 -23537 0 1 13286
box 22810 -13247 39241 -9665
use tps2_sw_stage_1  tps2_sw_stage_1_0
timestamp 1750900893
transform 1 0 899 0 1 4200
box -169 -173 4803 1866
use tps2_sw_stage_1  tps2_sw_stage_1_1
timestamp 1750900893
transform 1 0 5741 0 1 4200
box -169 -173 4803 1866
use tps2_sw_stage_1  tps2_sw_stage_1_2
timestamp 1750900893
transform 1 0 10583 0 1 4200
box -169 -173 4803 1866
use tps2_sw_stage_2  tps2_sw_stage_2_0
timestamp 1750900893
transform 1 0 5734 0 1 6234
box -162 -1648 5722 817
use tps2_sw_stage_3  tps2_sw_stage_3_0
timestamp 1750900893
transform 1 0 11482 0 1 6257
box -156 -189 2416 794
<< labels >>
flabel metal2 s -566 2941 -566 2941 6 FreeSans 320 0 0 0 V0
port 0 sw
flabel metal2 s 15574 2966 15574 2966 6 FreeSans 480 0 0 0 V48
port 1 sw
flabel metal2 s 921 4358 921 4358 6 FreeSans 480 0 0 0 DEC0[0]
port 2 sw
flabel metal2 s 5751 4361 5751 4361 6 FreeSans 480 0 0 0 DEC0[1]
port 3 sw
flabel metal2 s 11704 4361 11704 4361 6 FreeSans 480 0 0 0 DEC0[2]
port 4 sw
flabel metal2 s 11746 6400 11746 6400 6 FreeSans 480 0 0 0 DEC2[0]
port 9 sw
flabel metal2 s 12327 6403 12327 6403 6 FreeSans 480 0 0 0 DEC2[1]
port 10 sw
flabel metal2 s 12902 6399 12902 6399 6 FreeSans 480 0 0 0 DEC2[2]
port 11 sw
flabel metal2 s 13473 6409 13473 6409 6 FreeSans 480 0 0 0 DEC2[3]
port 12 sw
flabel metal2 s 13661 6751 13661 6751 6 FreeSans 480 0 0 0 VH
port 13 sw
flabel metal2 s 13311 6666 13311 6666 6 FreeSans 480 0 0 0 VL
port 14 sw
flabel locali s 13711 5311 13711 5311 6 FreeSans 800 0 0 0 GND
port 15 sw
flabel metal2 s 10501 6413 10501 6413 6 FreeSans 480 0 0 0 DEC1[0]
port 5 sw
flabel metal2 s 6031 6413 6031 6413 6 FreeSans 480 0 0 0 DEC1[1]
port 6 sw
flabel metal2 s 7436 6392 7436 6392 6 FreeSans 480 0 0 0 DEC1[2]
port 7 sw
flabel metal2 s 9028 6412 9028 6412 6 FreeSans 480 0 0 0 DEC1[3]
port 8 sw
<< end >>
