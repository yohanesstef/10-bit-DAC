magic
tech sky130A
magscale 1 2
timestamp 1751045299
<< pwell >>
rect 14692 13579 15422 14791
<< mvpsubdiff >>
rect 14728 14697 15386 14755
rect 14728 13673 14786 14697
rect 15328 13673 15386 14697
rect 14728 13615 15386 13673
<< locali >>
rect 14740 14709 15374 14743
rect 14740 13661 14774 14709
rect 15340 13661 15374 14709
rect 14740 13627 15374 13661
<< metal1 >>
rect 14952 14730 15004 14736
rect 14952 14644 15004 14678
rect 15110 14592 15162 14598
rect 14866 13747 14912 14578
rect 14952 14481 15004 14487
rect 14952 14395 15004 14429
rect 15110 14343 15162 14349
rect 14952 14232 15004 14238
rect 14952 14149 15004 14180
rect 15110 14094 15162 14100
rect 14952 13983 15004 13989
rect 14952 13900 15004 13931
rect 15110 13845 15162 13851
rect 15202 13747 15248 14578
<< via1 >>
rect 14952 14678 15004 14730
rect 15110 14598 15162 14650
rect 14952 14429 15004 14481
rect 15110 14349 15162 14401
rect 14952 14180 15004 14232
rect 15110 14100 15162 14152
rect 14952 13931 15004 13983
rect 15110 13851 15162 13903
<< metal2 >>
rect 14946 14678 14952 14730
rect 15004 14678 15010 14730
rect 15104 14598 15110 14650
rect 15162 14598 15168 14650
rect 14946 14429 14952 14481
rect 15004 14429 15010 14481
rect 15104 14349 15110 14401
rect 15162 14349 15168 14401
rect 14946 14180 14952 14232
rect 15004 14180 15010 14232
rect 15104 14100 15110 14152
rect 15162 14100 15168 14152
rect 14946 13931 14952 13983
rect 15004 13931 15010 13983
rect 15104 13851 15110 13903
rect 15162 13851 15168 13903
use sky130_fd_pr__nfet_g5v0d10v5_CSEDJZ  sky130_fd_pr__nfet_g5v0d10v5_CSEDJZ_0
timestamp 1751042016
transform 1 0 15057 0 1 13820
box -187 -99 187 99
use sky130_fd_pr__nfet_g5v0d10v5_CSEDJZ  sky130_fd_pr__nfet_g5v0d10v5_CSEDJZ_1
timestamp 1751042016
transform 1 0 15057 0 1 14069
box -187 -99 187 99
use sky130_fd_pr__nfet_g5v0d10v5_CSEDJZ  sky130_fd_pr__nfet_g5v0d10v5_CSEDJZ_2
timestamp 1751042016
transform 1 0 15057 0 1 14318
box -187 -99 187 99
use sky130_fd_pr__nfet_g5v0d10v5_CSEDJZ  sky130_fd_pr__nfet_g5v0d10v5_CSEDJZ_3
timestamp 1751042016
transform 1 0 15057 0 1 14567
box -187 -99 187 99
<< end >>
