.include /home/yohanes/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.subckt nand_hvl A B X GND VDDH
x1 A B GND GND VDDH VDDH X sky130_fd_sc_hvl__nand2_1
.ends

