** sch_path: /mnt/disk1/home/yohanes/10-bit-DAC/xschem/logic_shift_seg2.sch
**.subckt logic_shift_seg2 b[6],b[7],b[8],b[9] bb[6],bb[7],bb[8] BS[8],BS[9] VDD GND
*.ipin b[6],b[7],b[8],b[9]
*.opin BS[8],BS[9]
*.ipin GND
*.ipin VDD
*.ipin bb[6],bb[7],bb[8]
x1 b[9] b[8] GND GND VDD VDD n1 sky130_fd_sc_hd__nand2_1
x2 b[9] b[7] GND GND VDD VDD n2 sky130_fd_sc_hd__nand2_1
x3 b[9] b[6] GND GND VDD VDD n3 sky130_fd_sc_hd__nand2_1
x5 bb[8] bb[7] bb[6] GND GND VDD VDD n6 sky130_fd_sc_hd__nand3_1
x4 n3 n2 n1 GND GND VDD VDD BS[9] sky130_fd_sc_hd__nand3_1
x6 b[6] b[8] GND GND VDD VDD n4 sky130_fd_sc_hd__nand2_1
x7 b[7] b[8] GND GND VDD VDD n5 sky130_fd_sc_hd__nand2_1
x8 n6 n5 n4 GND GND VDD VDD BS[8] sky130_fd_sc_hd__nand3_1
**.ends
.end
