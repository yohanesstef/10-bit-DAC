magic
tech sky130A
magscale 1 2
timestamp 1749548291
<< error_s >>
rect 38897 -4596 38903 -4590
rect 38951 -4596 38957 -4590
rect 38891 -4602 38897 -4596
rect 38957 -4602 38963 -4596
rect 38891 -4656 38897 -4650
rect 38957 -4656 38963 -4650
rect 38897 -4662 38903 -4656
rect 38951 -4662 38957 -4656
rect 38621 -4684 38627 -4678
rect 38675 -4684 38681 -4678
rect 38615 -4690 38621 -4684
rect 38681 -4690 38687 -4684
rect 38615 -4744 38621 -4738
rect 38681 -4744 38687 -4738
rect 38621 -4750 38627 -4744
rect 38675 -4750 38681 -4744
rect 38345 -4772 38351 -4766
rect 38399 -4772 38405 -4766
rect 38339 -4778 38345 -4772
rect 38405 -4778 38411 -4772
rect 38339 -4832 38345 -4826
rect 38405 -4832 38411 -4826
rect 38345 -4838 38351 -4832
rect 38399 -4838 38405 -4832
rect 38069 -4860 38075 -4854
rect 38123 -4860 38129 -4854
rect 38063 -4866 38069 -4860
rect 38129 -4866 38135 -4860
rect 38063 -4920 38069 -4914
rect 38129 -4920 38135 -4914
rect 38069 -4926 38075 -4920
rect 38123 -4926 38129 -4920
rect 37765 -4948 37771 -4942
rect 37819 -4948 37825 -4942
rect 37759 -4954 37765 -4948
rect 37825 -4954 37831 -4948
rect 37759 -5008 37765 -5002
rect 37825 -5008 37831 -5002
rect 37765 -5014 37771 -5008
rect 37819 -5014 37825 -5008
rect 37489 -5036 37495 -5030
rect 37543 -5036 37549 -5030
rect 37483 -5042 37489 -5036
rect 37549 -5042 37555 -5036
rect 37483 -5096 37489 -5090
rect 37549 -5096 37555 -5090
rect 37489 -5102 37495 -5096
rect 37543 -5102 37549 -5096
rect 37213 -5124 37219 -5118
rect 37267 -5124 37273 -5118
rect 37207 -5130 37213 -5124
rect 37273 -5130 37279 -5124
rect 37207 -5184 37213 -5178
rect 37273 -5184 37279 -5178
rect 37213 -5190 37219 -5184
rect 37267 -5190 37273 -5184
rect 36937 -5212 36943 -5206
rect 36991 -5212 36997 -5206
rect 36931 -5218 36937 -5212
rect 36997 -5218 37003 -5212
rect 36931 -5272 36937 -5266
rect 36997 -5272 37003 -5266
rect 36937 -5278 36943 -5272
rect 36991 -5278 36997 -5272
<< pwell >>
rect 35000 -4677 39284 -4139
<< mvpsubdiff >>
rect 35036 -4187 39248 -4175
rect 35036 -4221 35144 -4187
rect 39140 -4221 39248 -4187
rect 35036 -4233 39248 -4221
rect 35036 -4283 35094 -4233
rect 35036 -4533 35048 -4283
rect 35082 -4533 35094 -4283
rect 35036 -4583 35094 -4533
rect 39190 -4283 39248 -4233
rect 39190 -4533 39202 -4283
rect 39236 -4533 39248 -4283
rect 39190 -4583 39248 -4533
rect 35036 -4595 39248 -4583
rect 35036 -4629 35144 -4595
rect 39140 -4629 39248 -4595
rect 35036 -4641 39248 -4629
<< mvpsubdiffcont >>
rect 35144 -4221 39140 -4187
rect 35048 -4533 35082 -4283
rect 39202 -4533 39236 -4283
rect 35144 -4629 39140 -4595
<< locali >>
rect 35048 -4221 35144 -4187
rect 39140 -4221 39236 -4187
rect 35048 -4283 35082 -4221
rect 35048 -4595 35082 -4533
rect 39202 -4283 39236 -4221
rect 39202 -4595 39236 -4533
rect 35048 -4629 35144 -4595
rect 39140 -4629 39236 -4595
<< metal1 >>
rect 35950 -3867 36010 -3861
rect 35352 -4043 35412 -4037
rect 35144 -4131 35204 -4125
rect 35144 -4481 35204 -4191
rect 35352 -4481 35412 -4103
rect 35752 -4043 35812 -4037
rect 35448 -4131 35508 -4125
rect 35448 -4481 35508 -4191
rect 35656 -4131 35716 -4125
rect 35656 -4481 35716 -4191
rect 35752 -4481 35812 -4103
rect 35950 -4282 36010 -3927
rect 36236 -3955 36296 -3949
rect 35960 -4393 36010 -4282
rect 35950 -4481 36010 -4393
rect 36038 -4131 36098 -4125
rect 36038 -4282 36098 -4191
rect 36038 -4393 36088 -4282
rect 36038 -4481 36098 -4393
rect 36236 -4481 36296 -4015
rect 36332 -4043 36392 -4037
rect 36332 -4481 36392 -4103
rect 36530 -4043 36590 -4037
rect 36530 -4282 36590 -4103
rect 36540 -4393 36590 -4282
rect 36530 -4481 36590 -4393
rect 36618 -4131 36678 -4125
rect 36618 -4282 36678 -4191
rect 36816 -4131 36876 -4125
rect 36618 -4393 36668 -4282
rect 36618 -4481 36678 -4393
rect 36816 -4481 36876 -4191
<< via1 >>
rect 35950 -3927 36010 -3867
rect 35352 -4103 35412 -4043
rect 35144 -4191 35204 -4131
rect 35752 -4103 35812 -4043
rect 35448 -4191 35508 -4131
rect 35656 -4191 35716 -4131
rect 36236 -4015 36296 -3955
rect 36038 -4191 36098 -4131
rect 36332 -4103 36392 -4043
rect 36530 -4103 36590 -4043
rect 36618 -4191 36678 -4131
rect 36816 -4191 36876 -4131
<< metal2 >>
rect 35944 -3927 35950 -3867
rect 36010 -3927 39146 -3867
rect 36230 -4015 36236 -3955
rect 36296 -4015 38870 -3955
rect 35346 -4103 35352 -4043
rect 35412 -4103 35752 -4043
rect 35812 -4103 36332 -4043
rect 36392 -4103 36398 -4043
rect 36524 -4103 36530 -4043
rect 36590 -4103 38594 -4043
rect 35138 -4191 35144 -4131
rect 35204 -4191 35448 -4131
rect 35508 -4191 35514 -4131
rect 35650 -4191 35656 -4131
rect 35716 -4191 36038 -4131
rect 36098 -4191 36618 -4131
rect 36678 -4191 36684 -4131
rect 36810 -4191 36816 -4131
rect 36876 -4191 38318 -4131
use hnmos_1  hnmos_1_0
timestamp 1749548291
transform 1 0 35485 0 1 -4510
box -41 3 235 201
use hnmos_1  hnmos_1_1
timestamp 1749548291
transform 1 0 35181 0 1 -4510
box -41 3 235 201
use hnmos_2  hnmos_2_0
timestamp 1749548291
transform 1 0 36332 0 1 -4508
box -4 1 548 199
use hnmos_2  hnmos_2_1
timestamp 1749548291
transform 1 0 35752 0 1 -4508
box -4 1 548 199
use nswitch_4_stage_3  nswitch_4_stage_3_0
timestamp 1749548291
transform 1 0 36874 0 1 -4551
box 34 -727 1140 690
use nswitch_4_stage_3_H  nswitch_4_stage_3_H_0
timestamp 1749548291
transform 1 0 38006 0 1 -4551
box 34 -375 1140 690
<< end >>
