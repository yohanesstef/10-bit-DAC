magic
tech sky130A
magscale 1 2
timestamp 1750166649
<< nwell >>
rect 1957 1661 4889 2977
<< metal1 >>
rect 3017 2525 3077 2531
rect 2559 2408 2701 2468
rect 2641 2173 2701 2408
rect 2770 2261 2830 2267
rect 3017 2230 3077 2465
rect 3146 2437 3206 2443
rect 3146 2371 3206 2377
rect 3271 2349 3317 2420
rect 3258 2289 3264 2349
rect 3324 2289 3330 2349
rect 2770 2195 2830 2201
rect 2941 2170 3077 2230
rect 2641 2107 2701 2113
rect 3393 1825 3453 2776
rect 3898 2525 3958 2531
rect 3898 2459 3958 2465
rect 3769 2437 3829 2443
rect 4063 2408 4205 2468
rect 3516 2289 3522 2349
rect 3582 2289 3588 2349
rect 3529 2230 3575 2289
rect 3769 2230 3829 2377
rect 4145 2261 4205 2408
rect 3693 2170 3829 2230
rect 3899 2170 3911 2230
rect 4145 2195 4205 2201
rect 4274 2173 4334 2179
rect 4274 2107 4334 2113
<< via1 >>
rect 3017 2465 3077 2525
rect 2770 2201 2830 2261
rect 3146 2377 3206 2437
rect 3264 2289 3324 2349
rect 2641 2113 2701 2173
rect 3898 2465 3958 2525
rect 3769 2377 3829 2437
rect 3522 2289 3582 2349
rect 4145 2201 4205 2261
rect 4274 2113 4334 2173
<< metal2 >>
rect 3011 2465 3017 2525
rect 3077 2465 3898 2525
rect 3958 2465 3964 2525
rect 3140 2377 3146 2437
rect 3206 2377 3769 2437
rect 3829 2377 3835 2437
rect 3258 2289 3264 2349
rect 3324 2289 3522 2349
rect 3582 2289 3588 2349
rect 2764 2201 2770 2261
rect 2830 2201 4145 2261
rect 4205 2201 4211 2261
rect 2635 2113 2641 2173
rect 2701 2113 4274 2173
rect 4334 2113 4340 2173
use cm2_pcell1_5  cm2_pcell1_5_0 ~/10-bit-DAC/mag
timestamp 1750158893
transform 1 0 3325 0 1 2116
box -1368 137 1564 861
use cm2_pcell1_5  cm2_pcell1_5_1
timestamp 1750158893
transform -1 0 3521 0 -1 2522
box -1368 137 1564 861
<< end >>
