magic
tech sky130A
magscale 1 2
timestamp 1749731508
<< magnet >>
rect 9 706 69 734
rect 1269 706 1329 734
rect 69 650 135 706
rect 195 650 261 706
rect 321 650 387 706
rect 447 650 513 706
rect 573 650 639 706
rect 699 650 765 706
rect 825 650 891 706
rect 951 650 1017 706
rect 1077 650 1143 706
rect 1203 650 1269 706
rect 135 622 195 650
rect 261 622 321 650
rect 387 622 447 650
rect 513 622 573 650
rect 639 622 699 650
rect 765 622 825 650
rect 891 622 951 650
rect 1017 622 1077 650
rect 1143 622 1203 650
rect 69 566 135 622
rect 195 566 261 622
rect 321 566 387 622
rect 447 566 513 622
rect 573 566 639 622
rect 699 566 765 622
rect 825 566 891 622
rect 951 566 1017 622
rect 1077 566 1143 622
rect 1203 566 1269 622
rect 135 538 195 566
rect 261 538 321 566
rect 387 538 447 566
rect 513 538 573 566
rect 639 538 699 566
rect 765 538 825 566
rect 891 538 951 566
rect 1017 538 1077 566
rect 1143 538 1203 566
rect 69 482 135 538
rect 195 482 261 538
rect 321 482 387 538
rect 447 482 513 538
rect 573 482 639 538
rect 699 482 765 538
rect 825 482 891 538
rect 951 482 1017 538
rect 1077 482 1143 538
rect 1203 482 1269 538
rect 135 454 195 482
rect 261 454 321 482
rect 387 454 447 482
rect 513 454 573 482
rect 639 454 699 482
rect 765 454 825 482
rect 891 454 951 482
rect 1017 454 1077 482
rect 1143 454 1203 482
rect 69 398 135 454
rect 195 398 261 454
rect 321 398 387 454
rect 447 398 513 454
rect 573 398 639 454
rect 699 398 765 454
rect 825 398 891 454
rect 951 398 1017 454
rect 1077 398 1143 454
rect 1203 398 1269 454
rect 135 370 195 398
rect 261 370 321 398
rect 387 370 447 398
rect 513 370 573 398
rect 639 370 699 398
rect 765 370 825 398
rect 891 370 951 398
rect 1017 370 1077 398
rect 1143 370 1203 398
rect 69 314 135 370
rect 195 314 261 370
rect 321 314 387 370
rect 447 314 513 370
rect 573 314 639 370
rect 699 314 765 370
rect 825 314 891 370
rect 951 314 1017 370
rect 1077 314 1143 370
rect 1203 314 1269 370
rect 135 286 195 314
rect 261 286 321 314
rect 387 286 447 314
rect 513 286 573 314
rect 639 286 699 314
rect 765 286 825 314
rect 891 286 951 314
rect 1017 286 1077 314
rect 1143 286 1203 314
rect 69 230 135 286
rect 195 230 261 286
rect 321 230 387 286
rect 447 230 513 286
rect 573 230 639 286
rect 699 230 765 286
rect 825 230 891 286
rect 951 230 1017 286
rect 1077 230 1143 286
rect 1203 230 1269 286
rect 135 202 195 230
rect 261 202 321 230
rect 387 202 447 230
rect 513 202 573 230
rect 639 202 699 230
rect 765 202 825 230
rect 891 202 951 230
rect 1017 202 1077 230
rect 1143 202 1203 230
rect 69 146 135 202
rect 195 146 261 202
rect 321 146 387 202
rect 447 146 513 202
rect 573 146 639 202
rect 699 146 765 202
rect 825 146 891 202
rect 951 146 1017 202
rect 1077 146 1143 202
rect 1203 146 1269 202
rect 135 118 195 146
rect 261 118 321 146
rect 387 118 447 146
rect 513 118 573 146
rect 639 118 699 146
rect 765 118 825 146
rect 891 118 951 146
rect 1017 118 1077 146
rect 1143 118 1203 146
rect 69 62 135 118
rect 195 62 261 118
rect 321 62 387 118
rect 447 62 513 118
rect 573 62 639 118
rect 699 62 765 118
rect 825 62 891 118
rect 951 62 1017 118
rect 1077 62 1143 118
rect 1203 62 1269 118
rect 135 34 195 62
rect 261 34 321 62
rect 387 34 447 62
rect 513 34 573 62
rect 639 34 699 62
rect 765 34 825 62
rect 891 34 951 62
rect 1017 34 1077 62
rect 1143 34 1203 62
rect 69 -22 135 34
rect 195 -22 261 34
rect 321 -22 387 34
rect 447 -22 513 34
rect 573 -22 639 34
rect 699 -22 765 34
rect 825 -22 891 34
rect 951 -22 1017 34
rect 1077 -22 1143 34
rect 1203 -22 1269 34
rect 135 -50 195 -22
rect 261 -50 321 -22
rect 387 -50 447 -22
rect 513 -50 573 -22
rect 639 -50 699 -22
rect 765 -50 825 -22
rect 891 -50 951 -22
rect 1017 -50 1077 -22
rect 1143 -50 1203 -22
rect 69 -106 135 -50
rect 195 -106 261 -50
rect 321 -106 387 -50
rect 447 -106 513 -50
rect 573 -106 639 -50
rect 699 -106 765 -50
rect 825 -106 891 -50
rect 951 -106 1017 -50
rect 1077 -106 1143 -50
rect 1203 -106 1269 -50
rect 9 -134 69 -106
rect 1269 -134 1329 -106
<< end >>
