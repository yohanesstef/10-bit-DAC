magic
tech sky130A
magscale 1 2
timestamp 1751058216
<< pwell >>
rect 18478 19848 18606 23430
rect 25955 1186 26083 4768
<< viali >>
rect 15822 23334 16210 23394
rect 26626 23334 27014 23394
rect 13365 18634 13399 19086
rect 12204 5090 12238 5542
rect 18999 1222 19387 1282
rect 32950 1222 33338 1282
<< metal1 >>
rect 38434 26130 38645 26136
rect 38434 25930 38439 26130
rect 38639 25930 38645 26130
rect 38434 25924 38645 25930
rect 15816 24930 16216 24936
rect 13352 24230 13412 24236
rect 13352 23624 13412 23630
rect 13359 19086 13405 23624
rect 15816 23394 16216 24330
rect 15816 23334 15822 23394
rect 16210 23334 16216 23394
rect 15816 23322 16216 23334
rect 26620 24930 27020 24936
rect 26620 23394 27020 24330
rect 26620 23334 26626 23394
rect 27014 23334 27020 23394
rect 35433 24230 35668 24236
rect 35433 23391 35668 23630
rect 38172 24230 38407 24236
rect 38172 23371 38407 23630
rect 38489 23486 38589 25924
rect 45994 25630 46194 25636
rect 38489 23428 38589 23434
rect 42561 24230 42796 24236
rect 42561 23367 42796 23630
rect 26620 23322 27020 23334
rect 38489 23266 38589 23272
rect 38489 23160 38589 23166
rect 45994 19913 46194 25030
rect 46623 24930 46823 24936
rect 46623 21213 46823 24330
rect 13359 18634 13365 19086
rect 13399 18634 13405 19086
rect 13359 18622 13405 18634
rect 13975 16863 14035 17640
rect 15217 16951 15277 17632
rect 15217 16885 15277 16891
rect 16314 16951 16374 16957
rect 13975 16797 14035 16803
rect 16072 16863 16132 16869
rect 16072 13025 16132 16803
rect 16072 12959 16132 12965
rect 16187 13377 16247 13383
rect 16187 6636 16247 13317
rect 16314 13113 16374 16891
rect 16314 13047 16374 13053
rect 16471 12937 16531 17646
rect 16471 12871 16531 12877
rect 16787 13465 16847 13471
rect 16787 8083 16847 13405
rect 17327 12849 17387 17646
rect 17327 12783 17387 12789
rect 17467 12761 17527 12767
rect 16781 8031 16787 8083
rect 16847 8031 16853 8083
rect 17467 8060 17527 12701
rect 18173 12761 18233 17645
rect 18173 12695 18233 12701
rect 18764 12673 18824 17646
rect 20660 13993 20720 17092
rect 20660 13927 20720 13933
rect 21240 13905 21300 17092
rect 21240 13839 21300 13845
rect 21820 13817 21880 17092
rect 21820 13751 21880 13757
rect 22400 13729 22460 17092
rect 23654 14081 23714 17092
rect 25062 14345 25122 17092
rect 25062 14279 25122 14285
rect 26470 14257 26530 17092
rect 26470 14191 26530 14197
rect 27878 14169 27938 17092
rect 31892 14433 31952 19133
rect 46175 15635 46423 16035
rect 46523 15635 46529 16035
rect 46917 15635 46923 16035
rect 47023 15635 48623 16035
rect 49223 15635 49229 16035
rect 46623 15035 47923 15435
rect 48523 15035 48529 15435
rect 31892 14367 31952 14373
rect 49518 14500 49729 14506
rect 49518 14357 49523 14500
rect 46907 14297 46913 14357
rect 47013 14300 49523 14357
rect 49723 14300 49729 14500
rect 47013 14297 49729 14300
rect 49518 14294 49729 14297
rect 27878 14103 27938 14109
rect 23654 14015 23714 14021
rect 49518 13900 49729 13906
rect 31468 13817 31528 13823
rect 22400 13663 22460 13669
rect 26935 13729 26995 13735
rect 18764 12607 18824 12613
rect 22995 12673 23055 12679
rect 19967 12585 20027 12591
rect 19122 12409 19182 12415
rect 18543 12321 18603 12327
rect 18239 12233 18299 12239
rect 17938 12145 17998 12151
rect 17938 9141 17998 12085
rect 18239 9141 18299 12173
rect 18543 9142 18603 12261
rect 19122 9144 19182 12349
rect 19967 9143 20027 12525
rect 21112 12497 21172 12503
rect 21112 9141 21172 12437
rect 22995 8062 23055 12613
rect 16781 7587 16787 7639
rect 16847 7587 16853 7639
rect 16187 6578 16247 6584
rect 16787 6636 16847 7587
rect 26935 6659 26995 13669
rect 31468 8086 31528 13757
rect 49518 13713 49523 13900
rect 46907 13653 46913 13713
rect 47013 13700 49523 13713
rect 49723 13700 49729 13900
rect 47013 13694 49729 13700
rect 47013 13653 49578 13694
rect 49518 13300 49729 13306
rect 49518 13100 49523 13300
rect 49723 13100 49729 13300
rect 49518 13094 49729 13100
rect 49518 13069 49578 13094
rect 46907 13009 46913 13069
rect 47013 13009 49578 13069
rect 37333 12761 37393 12767
rect 32093 12673 32153 12679
rect 31462 8026 31468 8086
rect 31528 8026 31534 8086
rect 32093 8056 32153 12613
rect 36213 12585 36273 12591
rect 35068 12497 35128 12503
rect 33644 12409 33704 12415
rect 33039 12233 33099 12239
rect 33039 9132 33099 12173
rect 33340 12145 33400 12151
rect 33340 9132 33400 12085
rect 33644 9133 33704 12349
rect 34223 12321 34283 12327
rect 34223 9136 34283 12261
rect 35068 9134 35128 12437
rect 36213 9132 36273 12525
rect 37333 8071 37393 12701
rect 49518 12700 49729 12706
rect 49518 12500 49523 12700
rect 49723 12500 49729 12700
rect 49518 12494 49729 12500
rect 49518 12425 49578 12494
rect 46907 12365 46913 12425
rect 47013 12365 49578 12425
rect 49518 12100 49729 12106
rect 49518 11900 49523 12100
rect 49723 11900 49729 12100
rect 49518 11894 49729 11900
rect 49518 11781 49578 11894
rect 46907 11721 46913 11781
rect 47013 11721 49578 11781
rect 49518 11500 49729 11506
rect 49518 11300 49523 11500
rect 49723 11300 49729 11500
rect 49518 11294 49729 11300
rect 49518 11137 49578 11294
rect 46907 11077 46913 11137
rect 47013 11077 49578 11137
rect 49518 10900 49729 10906
rect 49518 10754 49523 10900
rect 49297 10700 49523 10754
rect 49723 10700 49729 10900
rect 49297 10694 49729 10700
rect 49297 10493 49357 10694
rect 46907 10433 46913 10493
rect 47013 10433 49357 10493
rect 49518 10300 49729 10306
rect 49518 10154 49523 10300
rect 49297 10100 49523 10154
rect 49723 10100 49729 10300
rect 49297 10094 49729 10100
rect 49297 9849 49357 10094
rect 46907 9789 46913 9849
rect 47013 9789 49357 9849
rect 49518 9700 49729 9706
rect 49518 9554 49523 9700
rect 49297 9500 49523 9554
rect 49723 9500 49729 9700
rect 49297 9494 49729 9500
rect 49297 9205 49357 9494
rect 46907 9145 46913 9205
rect 47013 9145 49357 9205
rect 49517 9100 49729 9106
rect 49517 8900 49523 9100
rect 49723 8900 49729 9100
rect 49517 8894 49729 8900
rect 49517 8561 49577 8894
rect 46907 8501 46913 8561
rect 47013 8501 49577 8561
rect 46623 7914 47923 8314
rect 48523 7914 48529 8314
rect 31462 7586 31468 7646
rect 31528 7586 31534 7646
rect 31468 6645 31528 7586
rect 46015 7314 46423 7714
rect 46523 7314 46529 7714
rect 46623 7314 46823 7714
rect 46917 7314 46923 7714
rect 47023 7314 48623 7714
rect 49223 7314 49229 7714
rect 31468 6593 31763 6645
rect 16787 6578 16847 6584
rect 12198 5542 12244 5554
rect 12198 5090 12204 5542
rect 12238 5090 12244 5542
rect 12198 993 12244 5090
rect 18993 1282 19393 1294
rect 18993 1222 18999 1282
rect 19387 1222 19393 1282
rect 12191 987 12251 993
rect 12191 381 12251 387
rect 18993 287 19393 1222
rect 18993 -319 19393 -313
rect 32944 1282 33344 1294
rect 32944 1222 32950 1282
rect 33338 1222 33344 1282
rect 32944 287 33344 1222
rect 40759 987 40959 6592
rect 40759 381 40959 387
rect 32944 -319 33344 -313
rect 46015 -413 46175 2384
rect 46623 287 46823 2838
rect 46623 -319 46823 -313
rect 46015 -1019 46175 -1013
<< via1 >>
rect 38439 25930 38639 26130
rect 15816 24330 16216 24930
rect 13352 23630 13412 24230
rect 26620 24330 27020 24930
rect 35433 23630 35668 24230
rect 38172 23630 38407 24230
rect 45994 25030 46194 25630
rect 38489 23434 38589 23486
rect 42561 23630 42796 24230
rect 38489 23166 38589 23266
rect 46623 24330 46823 24930
rect 15217 16891 15277 16951
rect 16314 16891 16374 16951
rect 13975 16803 14035 16863
rect 16072 16803 16132 16863
rect 16072 12965 16132 13025
rect 16187 13317 16247 13377
rect 16314 13053 16374 13113
rect 16471 12877 16531 12937
rect 16787 13405 16847 13465
rect 17327 12789 17387 12849
rect 17467 12701 17527 12761
rect 16787 8031 16847 8083
rect 18173 12701 18233 12761
rect 20660 13933 20720 13993
rect 21240 13845 21300 13905
rect 21820 13757 21880 13817
rect 25062 14285 25122 14345
rect 26470 14197 26530 14257
rect 46423 15635 46523 16035
rect 46923 15635 47023 16035
rect 48623 15635 49223 16035
rect 47923 15035 48523 15435
rect 31892 14373 31952 14433
rect 46913 14297 47013 14357
rect 49523 14300 49723 14500
rect 27878 14109 27938 14169
rect 23654 14021 23714 14081
rect 31468 13757 31528 13817
rect 22400 13669 22460 13729
rect 26935 13669 26995 13729
rect 18764 12613 18824 12673
rect 22995 12613 23055 12673
rect 19967 12525 20027 12585
rect 19122 12349 19182 12409
rect 18543 12261 18603 12321
rect 18239 12173 18299 12233
rect 17938 12085 17998 12145
rect 21112 12437 21172 12497
rect 16787 7587 16847 7639
rect 16187 6584 16247 6636
rect 46913 13653 47013 13713
rect 49523 13700 49723 13900
rect 49523 13100 49723 13300
rect 46913 13009 47013 13069
rect 37333 12701 37393 12761
rect 32093 12613 32153 12673
rect 31468 8026 31528 8086
rect 36213 12525 36273 12585
rect 35068 12437 35128 12497
rect 33644 12349 33704 12409
rect 33039 12173 33099 12233
rect 33340 12085 33400 12145
rect 34223 12261 34283 12321
rect 49523 12500 49723 12700
rect 46913 12365 47013 12425
rect 49523 11900 49723 12100
rect 46913 11721 47013 11781
rect 49523 11300 49723 11500
rect 46913 11077 47013 11137
rect 49523 10700 49723 10900
rect 46913 10433 47013 10493
rect 49523 10100 49723 10300
rect 46913 9789 47013 9849
rect 49523 9500 49723 9700
rect 46913 9145 47013 9205
rect 49523 8900 49723 9100
rect 46913 8501 47013 8561
rect 47923 7914 48523 8314
rect 31468 7586 31528 7646
rect 16787 6584 16847 6636
rect 46423 7314 46523 7714
rect 46923 7314 47023 7714
rect 48623 7314 49223 7714
rect 12191 387 12251 987
rect 18993 -313 19393 287
rect 40759 387 40959 987
rect 32944 -313 33344 287
rect 46623 -313 46823 287
rect 46015 -1013 46175 -413
<< metal2 >>
rect 38339 26130 38739 26230
rect 38339 25930 38439 26130
rect 38639 25930 38739 26130
rect 38339 25830 38739 25930
rect -1226 25030 45994 25630
rect 46194 25030 49223 25630
rect -1226 24330 15816 24930
rect 16216 24330 26620 24930
rect 27020 24330 46623 24930
rect 46823 24330 48523 24930
rect -1226 23630 13352 24230
rect 13412 23630 35433 24230
rect 35668 23630 38172 24230
rect 38407 23630 42561 24230
rect 42796 23630 47823 24230
rect 38489 23486 38589 23492
rect 38489 23266 38589 23434
rect 38489 23160 38589 23166
rect 18478 20374 18616 20636
rect 21430 19079 21440 19135
rect 21496 19079 21506 19135
rect 26262 19079 26272 19135
rect 26328 19079 26338 19135
rect 15886 18762 15896 18818
rect 15952 18762 15962 18818
rect 18405 18762 18415 18818
rect 18471 18762 18481 18818
rect 15211 16891 15217 16951
rect 15277 16891 16314 16951
rect 16374 16891 16380 16951
rect 13969 16803 13975 16863
rect 14035 16803 16072 16863
rect 16132 16803 16138 16863
rect 46417 15635 46423 16035
rect 46523 15635 46923 16035
rect 47023 15635 47029 16035
rect 21430 14551 21440 14607
rect 21496 14551 21506 14607
rect 26263 14463 26273 14519
rect 26329 14463 26339 14519
rect 46719 14297 46913 14357
rect 47013 14297 47019 14357
rect 38148 13936 38158 13992
rect 38214 13936 38224 13992
rect 34815 13845 34825 13901
rect 34881 13845 34891 13901
rect 46719 13653 46913 13713
rect 47013 13653 47019 13713
rect 23482 13583 23492 13639
rect 23548 13583 23558 13639
rect 20149 13495 20159 13551
rect 20215 13495 20225 13551
rect 15886 13231 15896 13287
rect 15952 13231 15962 13287
rect 18405 13143 18415 13199
rect 18471 13143 18481 13199
rect 46719 13009 46913 13069
rect 47013 13009 47019 13069
rect 46719 12365 46913 12425
rect 47013 12365 47019 12425
rect 15856 11997 19628 12057
rect 15856 11909 19628 11969
rect 15856 11821 19628 11881
rect 15856 11733 19628 11793
rect 46719 11721 46913 11781
rect 47013 11721 47019 11781
rect 46719 11077 46913 11137
rect 47013 11077 47019 11137
rect 46719 10433 46913 10493
rect 47013 10433 47019 10493
rect 46719 9789 46913 9849
rect 47013 9789 47019 9849
rect 46719 9145 46913 9205
rect 47013 9145 47019 9205
rect 46719 8501 46913 8561
rect 47013 8501 47019 8561
rect 16781 8031 16787 8083
rect 16847 8031 16853 8083
rect 16787 7639 16847 8031
rect 31462 8026 31468 8086
rect 31528 8026 31534 8086
rect 31468 7646 31528 8026
rect 16781 7587 16787 7639
rect 16847 7587 16853 7639
rect 31462 7586 31468 7646
rect 31528 7586 31534 7646
rect 46417 7314 46423 7714
rect 46523 7314 46923 7714
rect 47023 7314 47029 7714
rect 16078 6584 16187 6636
rect 16247 6584 16253 6636
rect 16781 6584 16787 6636
rect 16847 6584 17024 6636
rect 20147 6584 20157 6640
rect 20213 6584 20223 6640
rect 23482 6584 23492 6640
rect 23548 6584 23558 6640
rect 34818 6591 34828 6647
rect 34884 6645 34894 6647
rect 34884 6593 35057 6645
rect 34884 6591 34894 6593
rect 38151 6591 38161 6647
rect 38217 6591 38227 6647
rect 47223 987 47823 23630
rect -1226 387 12191 987
rect 12251 387 24183 987
rect 24773 387 40759 987
rect 40959 387 47823 987
rect 47923 15435 48523 24330
rect 47923 8314 48523 15035
rect 47923 287 48523 7914
rect -1226 -313 18993 287
rect 19393 -313 27737 287
rect 28327 -313 32944 287
rect 33344 -313 46623 287
rect 46823 -313 48523 287
rect 48623 16035 49223 25030
rect 48623 7714 49223 15635
rect 49423 14500 49823 14600
rect 49423 14300 49523 14500
rect 49723 14300 49823 14500
rect 49423 14200 49823 14300
rect 49423 13900 49823 14000
rect 49423 13700 49523 13900
rect 49723 13700 49823 13900
rect 49423 13600 49823 13700
rect 49423 13300 49823 13400
rect 49423 13100 49523 13300
rect 49723 13100 49823 13300
rect 49423 13000 49823 13100
rect 49423 12700 49823 12800
rect 49423 12500 49523 12700
rect 49723 12500 49823 12700
rect 49423 12400 49823 12500
rect 49423 12100 49823 12200
rect 49423 11900 49523 12100
rect 49723 11900 49823 12100
rect 49423 11800 49823 11900
rect 49423 11500 49823 11600
rect 49423 11300 49523 11500
rect 49723 11300 49823 11500
rect 49423 11200 49823 11300
rect 49423 10900 49823 11000
rect 49423 10700 49523 10900
rect 49723 10700 49823 10900
rect 49423 10600 49823 10700
rect 49423 10300 49823 10400
rect 49423 10100 49523 10300
rect 49723 10100 49823 10300
rect 49423 10000 49823 10100
rect 49423 9700 49823 9800
rect 49423 9500 49523 9700
rect 49723 9500 49823 9700
rect 49423 9400 49823 9500
rect 49423 9100 49823 9200
rect 49423 8900 49523 9100
rect 49723 8900 49823 9100
rect 49423 8800 49823 8900
rect 48623 -413 49223 7314
rect -1226 -1013 46015 -413
rect 46175 -1013 49223 -413
<< via2 >>
rect 13850 20385 14009 20626
rect 34162 20383 34535 20626
rect 21440 19079 21496 19135
rect 26272 19079 26328 19135
rect 15896 18762 15952 18818
rect 18415 18762 18471 18818
rect 21440 14551 21496 14607
rect 26273 14463 26329 14519
rect 38158 13936 38214 13992
rect 34825 13845 34881 13901
rect 23492 13583 23548 13639
rect 20159 13495 20215 13551
rect 15896 13231 15952 13287
rect 18415 13143 18471 13199
rect 20157 6584 20213 6640
rect 23492 6584 23548 6640
rect 34828 6591 34884 6647
rect 38161 6591 38217 6647
rect 13764 3987 13895 4236
rect 24187 3980 24765 4234
rect 27741 3980 28319 4234
rect 39860 3981 39997 4234
rect 24183 387 24773 987
rect 27737 -313 28327 287
<< metal3 >>
rect 13838 20626 17211 20636
rect 13838 20385 13850 20626
rect 14009 20385 17211 20626
rect 13838 20374 17211 20385
rect 15891 18818 15957 18828
rect 15891 18762 15896 18818
rect 15952 18762 15957 18818
rect 15891 18752 15957 18762
rect 15894 13297 15954 18752
rect 15891 13287 15957 13297
rect 15891 13231 15896 13287
rect 15952 13231 15957 13287
rect 15891 13221 15957 13231
rect 16811 4242 17211 20374
rect 34150 20626 34550 20636
rect 34150 20383 34162 20626
rect 34535 20383 34550 20626
rect 21435 19135 21501 19145
rect 21435 19079 21440 19135
rect 21496 19079 21501 19135
rect 21435 19069 21501 19079
rect 26267 19135 26333 19145
rect 26267 19079 26272 19135
rect 26328 19079 26333 19135
rect 26267 19069 26333 19079
rect 18410 18818 18476 18828
rect 18410 18762 18415 18818
rect 18471 18762 18476 18818
rect 18410 18752 18476 18762
rect 18413 17617 18473 18752
rect 18413 14343 18474 17617
rect 21438 14617 21498 19069
rect 21435 14607 21501 14617
rect 21435 14551 21440 14607
rect 21496 14551 21501 14607
rect 21435 14541 21501 14551
rect 26271 14529 26331 19069
rect 26268 14519 26334 14529
rect 26268 14463 26273 14519
rect 26329 14463 26334 14519
rect 26268 14453 26334 14463
rect 18413 13209 18473 14343
rect 23487 13639 23553 13649
rect 23487 13583 23492 13639
rect 23548 13583 23553 13639
rect 23487 13573 23553 13583
rect 20154 13551 20220 13561
rect 20154 13495 20159 13551
rect 20215 13495 20220 13551
rect 20154 13485 20220 13495
rect 18410 13199 18476 13209
rect 18410 13143 18415 13199
rect 18471 13143 18476 13199
rect 18410 13133 18476 13143
rect 20157 6650 20217 13485
rect 23490 6650 23550 13573
rect 20152 6640 20218 6650
rect 20152 6584 20157 6640
rect 20213 6584 20218 6640
rect 20152 6574 20218 6584
rect 23487 6640 23553 6650
rect 23487 6584 23492 6640
rect 23548 6584 23553 6640
rect 23487 6574 23553 6584
rect 34150 4242 34550 20383
rect 38153 13992 38219 14002
rect 38153 13936 38158 13992
rect 38214 13936 38219 13992
rect 38153 13926 38219 13936
rect 34820 13901 34886 13911
rect 34820 13845 34825 13901
rect 34881 13845 34886 13901
rect 34820 13835 34886 13845
rect 34823 6657 34883 13835
rect 38156 6657 38216 13926
rect 34823 6647 34889 6657
rect 34823 6591 34828 6647
rect 34884 6591 34889 6647
rect 34823 6581 34889 6591
rect 38156 6647 38222 6657
rect 38156 6591 38161 6647
rect 38217 6591 38222 6647
rect 38156 6581 38222 6591
rect 13756 4236 17211 4242
rect 13756 3987 13764 4236
rect 13895 3987 17211 4236
rect 13756 3980 17211 3987
rect 24178 4234 24778 4242
rect 24178 3980 24187 4234
rect 24765 3980 24778 4234
rect 24178 987 24778 3980
rect 24178 387 24183 987
rect 24773 387 24778 987
rect 24178 382 24778 387
rect 27732 4234 28332 4242
rect 27732 3980 27741 4234
rect 28319 3980 28332 4234
rect 27732 287 28332 3980
rect 34150 4234 40015 4242
rect 34150 3981 39860 4234
rect 39997 3981 40015 4234
rect 34150 3970 40015 3981
rect 27732 -313 27737 287
rect 28327 -313 28332 287
rect 27732 -318 28332 -313
use top_dcell_routing  top_dcell_routing_0
timestamp 1751042016
transform 1 0 0 0 1 0
box 15856 1202 46823 23447
use top_segment_1  top_segment_1_0
timestamp 1750900893
transform 1 0 26106 0 1 1210
box -385 -24 14453 8429
use top_segment_2  top_segment_2_0
timestamp 1750900893
transform -1 0 34310 0 -1 23469
box -727 39 15704 7051
use top_segment_3  top_segment_3_0
timestamp 1749552768
transform -1 0 24112 0 -1 23696
box 5007 266 11251 6636
use top_segment_4  top_segment_4_1
timestamp 1749664768
transform 1 0 -17367 0 1 13412
box 29493 -12226 43322 -3773
<< labels >>
flabel metal2 s 38339 25830 38739 26230 0 FreeSans 800 0 0 0 ROUT
port 10 nsew
flabel metal2 s 49423 14200 49823 14600 0 FreeSans 800 0 0 0 DIN0
port 0 nsew
flabel metal2 s 49423 13600 49823 14000 0 FreeSans 800 0 0 0 DIN1
port 1 nsew
flabel metal2 s 49423 13000 49823 13400 0 FreeSans 800 0 0 0 DIN2
port 2 nsew
flabel metal2 s 49423 12400 49823 12800 0 FreeSans 800 0 0 0 DIN3
port 3 nsew
flabel metal2 s 49423 11800 49823 12200 0 FreeSans 800 0 0 0 DIN4
port 4 nsew
flabel metal2 s 49423 11200 49823 11600 0 FreeSans 800 0 0 0 DIN5
port 5 nsew
flabel metal2 s 49423 10600 49823 11000 0 FreeSans 800 0 0 0 DIN6
port 6 nsew
flabel metal2 s 49423 10000 49823 10400 0 FreeSans 800 0 0 0 DIN7
port 7 nsew
flabel metal2 s 49423 9400 49823 9800 0 FreeSans 800 0 0 0 DIN8
port 8 nsew
flabel metal2 s 49423 8800 49823 9200 0 FreeSans 800 0 0 0 DIN9
port 9 nsew
flabel metal2 s 32932 9309 32992 9369 0 FreeSans 800 0 0 0 VS1
port 11 nsew
flabel metal2 s 20842 16776 20902 16836 0 FreeSans 800 0 0 0 VL2
port 12 nsew
flabel metal2 s 20566 16688 20626 16748 0 FreeSans 800 0 0 0 VH2
port 13 nsew
flabel metal2 s 18575 17506 18635 17566 0 FreeSans 800 0 0 0 VL3
port 14 nsew
flabel metal2 s 18852 17418 18912 17478 0 FreeSans 800 0 0 0 VH3
port 15 nsew
flabel metal2 s -916 -1013 284 -413 0 FreeSans 4800 0 0 0 VDD
port 21 nsew
flabel metal2 s -916 387 284 987 0 FreeSans 4800 0 0 0 VDDH
port 22 nsew
flabel metal2 s -916 -313 284 287 0 FreeSans 4800 0 0 0 GND
port 23 nsew
flabel metal2 s 17831 9309 17891 9369 0 FreeSans 800 0 0 0 VS4
port 16 nsew
flabel metal2 s 15856 11733 15916 11793 0 FreeSans 480 0 0 0 SH[1]
port 17 nsew
flabel metal2 s 15856 11821 15916 11881 0 FreeSans 480 0 0 0 SH[2]
port 18 nsew
flabel metal2 s 15856 11909 15916 11969 0 FreeSans 480 0 0 0 SH[3]
port 19 nsew
flabel metal2 s 15856 11997 15916 12057 0 FreeSans 480 0 0 0 SH[4]
port 20 nsew
<< end >>
