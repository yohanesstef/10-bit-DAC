magic
tech sky130A
magscale 1 2
timestamp 1751053439
<< mvpsubdiffcont >>
rect 14515 14507 15029 14541
rect 14455 13219 14489 14481
rect 15055 14275 15089 14481
rect 15055 14241 15629 14275
rect 15055 13193 15089 14241
rect 15655 13219 15689 14215
rect 14515 13159 15630 13193
<< mvnsubdiffcont >>
rect 16517 14496 17023 14530
rect 16457 14044 16491 14470
rect 15925 14010 16491 14044
rect 15865 13227 15899 13984
rect 16457 13201 16491 14010
rect 17049 13227 17083 14470
rect 15925 13167 17023 13201
<< viali >>
rect 14515 14507 15029 14541
rect 16517 14496 17023 14530
<< metal1 >>
rect 14509 14541 15035 14553
rect 14509 14507 14515 14541
rect 15029 14507 15035 14541
rect 14509 14495 15035 14507
rect 14744 14345 14800 14351
rect 14744 14283 14800 14289
rect 14915 14287 14921 14339
rect 14973 14287 14979 14339
rect 14567 13111 14627 13279
rect 14679 13111 14707 14111
rect 14744 14096 14800 14102
rect 14744 14034 14800 14040
rect 14744 13847 14800 13853
rect 14744 13785 14800 13791
rect 14744 13598 14800 13604
rect 14744 13536 14800 13542
rect 14744 13349 14800 13355
rect 14744 13287 14800 13293
rect 14837 13111 14865 14111
rect 15167 14110 15227 14608
rect 15517 14110 15577 14608
rect 14915 14038 14921 14090
rect 14973 14038 14979 14090
rect 15340 14038 15346 14090
rect 15398 14038 15404 14090
rect 15973 13861 16033 14608
rect 16323 13869 16383 14608
rect 16511 14530 17037 14542
rect 16511 14496 16517 14530
rect 17023 14496 17037 14530
rect 16511 14484 17037 14496
rect 16742 14345 16798 14351
rect 16431 14263 16589 14293
rect 16742 14283 16798 14289
rect 16323 13861 16369 13869
rect 16431 13841 16461 14263
rect 16742 14096 16798 14102
rect 14915 13789 14921 13841
rect 14973 13789 14979 13841
rect 15340 13789 15346 13841
rect 15398 13789 15404 13841
rect 16146 13789 16152 13841
rect 16204 13789 16210 13841
rect 16397 13789 16403 13841
rect 16455 13789 16461 13841
rect 16489 14014 16589 14044
rect 16489 13761 16519 14014
rect 16431 13731 16519 13761
rect 16431 13592 16461 13731
rect 16589 13703 16619 13849
rect 14915 13540 14921 13592
rect 14973 13540 14979 13592
rect 15340 13540 15346 13592
rect 15398 13540 15404 13592
rect 16146 13540 16152 13592
rect 16204 13540 16210 13592
rect 16397 13540 16403 13592
rect 16455 13540 16461 13592
rect 16489 13673 16619 13703
rect 16489 13343 16519 13673
rect 16589 13351 16619 13516
rect 15340 13291 15346 13343
rect 15398 13291 15404 13343
rect 16146 13291 16152 13343
rect 16204 13291 16210 13343
rect 16397 13291 16403 13343
rect 16455 13313 16519 13343
rect 16455 13291 16461 13313
rect 14907 13251 14953 13279
rect 15507 13251 15553 13279
rect 14907 13221 15553 13251
rect 16339 13263 16369 13283
rect 16589 13263 16619 13283
rect 16339 13233 16619 13263
rect 16677 13089 16705 14089
rect 16742 14034 16798 14040
rect 16742 13847 16798 13853
rect 16742 13785 16798 13791
rect 16742 13598 16798 13604
rect 16742 13536 16798 13542
rect 16742 13349 16798 13355
rect 16742 13287 16798 13293
rect 16835 13089 16863 14089
rect 16915 13089 16975 13267
<< via1 >>
rect 14744 14289 14800 14345
rect 14921 14287 14973 14339
rect 14744 14040 14800 14096
rect 14744 13791 14800 13847
rect 14744 13542 14800 13598
rect 14744 13293 14800 13349
rect 14921 14038 14973 14090
rect 15346 14038 15398 14090
rect 16742 14289 16798 14345
rect 14921 13789 14973 13841
rect 15346 13789 15398 13841
rect 16152 13789 16204 13841
rect 16403 13789 16455 13841
rect 14921 13540 14973 13592
rect 15346 13540 15398 13592
rect 16152 13540 16204 13592
rect 16403 13540 16455 13592
rect 15346 13291 15398 13343
rect 16152 13291 16204 13343
rect 16403 13291 16455 13343
rect 16742 14040 16798 14096
rect 16742 13791 16798 13847
rect 16742 13542 16798 13598
rect 16742 13293 16798 13349
<< metal2 >>
rect 14744 14345 14800 14355
rect 16742 14345 16798 14355
rect 14744 14279 14800 14289
rect 14915 14287 14921 14339
rect 14973 14309 15233 14339
rect 14973 14287 14979 14309
rect 14744 14096 14800 14106
rect 15203 14090 15233 14309
rect 16742 14279 16798 14289
rect 16125 14210 17161 14240
rect 16073 14152 17161 14182
rect 16742 14096 16798 14106
rect 14744 14030 14800 14040
rect 14915 14038 14921 14090
rect 14973 14060 15175 14090
rect 15203 14060 15346 14090
rect 14973 14038 14979 14060
rect 14744 13847 14800 13857
rect 15145 13841 15175 14060
rect 15340 14038 15346 14060
rect 15398 14038 15404 14090
rect 16742 14030 16798 14040
rect 16125 13961 17161 13991
rect 16125 13903 17161 13933
rect 16742 13847 16798 13857
rect 14744 13781 14800 13791
rect 14915 13789 14921 13841
rect 14973 13811 15117 13841
rect 15145 13811 15346 13841
rect 14973 13789 14979 13811
rect 14744 13598 14800 13608
rect 15087 13592 15117 13811
rect 15340 13789 15346 13811
rect 15398 13789 15404 13841
rect 16146 13789 16152 13841
rect 16204 13811 16403 13841
rect 16204 13789 16210 13811
rect 16397 13789 16403 13811
rect 16455 13789 16461 13841
rect 16742 13781 16798 13791
rect 16125 13712 17161 13742
rect 16125 13654 17161 13684
rect 16742 13598 16798 13608
rect 14744 13532 14800 13542
rect 14915 13540 14921 13592
rect 14973 13562 15059 13592
rect 15087 13562 15346 13592
rect 14973 13540 14979 13562
rect 14744 13349 14800 13359
rect 15029 13343 15059 13562
rect 15340 13540 15346 13562
rect 15398 13540 15404 13592
rect 16146 13540 16152 13592
rect 16204 13562 16403 13592
rect 16204 13540 16210 13562
rect 16397 13540 16403 13562
rect 16455 13540 16461 13592
rect 16742 13532 16798 13542
rect 16125 13463 17161 13493
rect 16131 13405 17161 13435
rect 16742 13349 16798 13359
rect 15029 13313 15346 13343
rect 14744 13283 14800 13293
rect 15340 13291 15346 13313
rect 15398 13291 15404 13343
rect 16146 13291 16152 13343
rect 16204 13313 16403 13343
rect 16204 13291 16210 13313
rect 16397 13291 16403 13313
rect 16455 13291 16461 13343
rect 16742 13283 16798 13293
<< via2 >>
rect 14744 14289 14800 14345
rect 14744 14040 14800 14096
rect 16742 14289 16798 14345
rect 14744 13791 14800 13847
rect 16742 14040 16798 14096
rect 14744 13542 14800 13598
rect 16742 13791 16798 13847
rect 14744 13293 14800 13349
rect 16742 13542 16798 13598
rect 16742 13293 16798 13349
<< metal3 >>
rect 14407 14350 16349 14351
rect 14407 14345 16808 14350
rect 14407 14289 14744 14345
rect 14800 14289 16742 14345
rect 16798 14289 16808 14345
rect 14407 14285 16808 14289
rect 14734 14284 16808 14285
rect 14407 14096 16808 14101
rect 14407 14040 14744 14096
rect 14800 14040 16742 14096
rect 16798 14040 16808 14096
rect 14407 14035 16808 14040
rect 14407 13847 16808 13852
rect 14407 13791 14744 13847
rect 14800 13791 16742 13847
rect 16798 13791 16808 13847
rect 14407 13786 16808 13791
rect 14407 13598 16808 13603
rect 14407 13542 14744 13598
rect 14800 13542 16742 13598
rect 16798 13542 16808 13598
rect 14407 13537 16808 13542
rect 14407 13349 16808 13354
rect 14407 13293 14744 13349
rect 14800 13293 16742 13349
rect 16798 13293 16808 13349
rect 14407 13288 16808 13293
use interpolation_switch  interpolation_switch_0 ~/10-bit-DAC/mag
timestamp 1751047215
transform 1 0 15195 0 1 13261
box -188 -172 1374 1062
use seg_sel_nmos  seg_sel_nmos_0
timestamp 1751047180
transform 1 0 15337 0 1 13280
box -930 -169 -200 1309
use seg_sel_pmos  seg_sel_pmos_0
timestamp 1751047404
transform 1 0 10148 0 1 12795
box 6231 294 7013 1813
<< labels >>
flabel metal2 s 17133 13463 17161 13491 0 FreeSans 160 0 0 0 b[0]
port 0 nsew
flabel metal2 s 17129 13712 17157 13740 0 FreeSans 160 0 0 0 b[1]
port 1 nsew
flabel metal2 s 17128 13961 17156 13989 0 FreeSans 160 0 0 0 b[2]
port 2 nsew
flabel metal2 s 17131 14210 17159 14238 0 FreeSans 160 0 0 0 b[3]
port 3 nsew
flabel metal2 s 17133 13405 17161 13433 0 FreeSans 160 0 0 0 bb[0]
port 4 nsew
flabel metal2 s 17129 13654 17157 13682 0 FreeSans 160 0 0 0 bb[1]
port 5 nsew
flabel metal2 s 17128 13903 17156 13931 0 FreeSans 160 0 0 0 bb[2]
port 6 nsew
flabel metal2 s 17131 14152 17159 14180 0 FreeSans 160 0 0 0 bb[3]
port 7 nsew
flabel metal1 s 14679 13111 14707 13139 0 FreeSans 160 0 0 0 SH[1]
port 8 nsew
flabel metal1 s 14837 13111 14865 13139 0 FreeSans 160 0 0 0 SH[2]
port 9 nsew
flabel metal1 s 16677 13089 16705 13117 0 FreeSans 160 0 0 0 SH[3]
port 10 nsew
flabel metal1 s 16835 13089 16863 13117 0 FreeSans 160 0 0 0 SH[4]
port 11 nsew
flabel metal1 s 14567 13111 14627 13171 0 FreeSans 160 0 0 0 VS1
port 12 nsew
flabel metal1 s 15973 14548 16033 14608 0 FreeSans 160 0 0 0 VH3
port 16 nsew
flabel metal1 s 16323 14548 16383 14608 0 FreeSans 160 0 0 0 VL3
port 15 nsew
flabel metal1 s 15517 14548 15577 14608 0 FreeSans 160 0 0 0 VL2
port 13 nsew
flabel metal1 s 15167 14548 15227 14608 0 FreeSans 160 0 0 0 VH2
port 14 nsew
flabel metal1 s 16915 13089 16975 13149 0 FreeSans 160 0 0 0 VS4
port 17 nsew
flabel metal3 s 14407 13537 14467 13603 0 FreeSans 160 0 0 0 VOUT[1]
port 19 nsew
flabel metal3 s 14407 13786 14467 13852 0 FreeSans 160 0 0 0 VOUT[2]
port 20 nsew
flabel metal3 s 14407 14035 14467 14101 0 FreeSans 160 0 0 0 VOUT[3]
port 21 nsew
flabel metal3 s 14407 14285 14467 14351 0 FreeSans 160 0 0 0 VOUT[4]
port 22 nsew
flabel metal3 s 14407 13288 14467 13354 0 FreeSans 160 0 0 0 VOUT[0]
port 18 nsew
flabel metal1 s 16511 14484 16571 14542 0 FreeSans 160 0 0 0 VDDH
port 23 nsew
flabel metal1 s 14509 14495 14569 14553 0 FreeSans 160 0 0 0 GND
port 24 nsew
<< end >>
