magic
tech sky130A
magscale 1 2
timestamp 1749844197
<< metal2 >>
rect 31 -25 1536 35
rect 31 -113 1536 -53
rect 31 -201 1536 -141
rect 31 -289 1536 -229
rect 31 -377 1536 -317
rect 31 -465 1536 -405
rect 31 -553 1536 -493
rect 31 -641 1536 -581
use cm_pcell1_4  cm_pcell1_4_0
timestamp 1749844197
transform 1 0 -14 0 1 -323
box -21 1 1625 678
use cm_pcell1_4  cm_pcell1_4_1
timestamp 1749844197
transform 1 0 -14 0 -1 -283
box -21 1 1625 678
<< end >>
