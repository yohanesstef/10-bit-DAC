magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -955 307 955
<< psubdiff >>
rect -271 885 -175 919
rect 175 885 271 919
rect -271 823 -237 885
rect 237 823 271 885
rect -271 -885 -237 -823
rect 237 -885 271 -823
rect -271 -919 -175 -885
rect 175 -919 271 -885
<< psubdiffcont >>
rect -175 885 175 919
rect -271 -823 -237 823
rect 237 -823 271 823
rect -175 -919 175 -885
<< xpolycontact >>
rect -141 357 141 789
rect -141 -789 141 -357
<< xpolyres >>
rect -141 -357 141 357
<< locali >>
rect -271 885 -175 919
rect 175 885 271 919
rect -271 823 -237 885
rect 237 823 271 885
rect -271 -885 -237 -823
rect 237 -885 271 -823
rect -271 -919 -175 -885
rect 175 -919 271 -885
<< viali >>
rect -125 374 125 771
rect -125 -771 125 -374
<< metal1 >>
rect -131 771 131 783
rect -131 374 -125 771
rect 125 374 131 771
rect -131 362 131 374
rect -131 -374 131 -362
rect -131 -771 -125 -374
rect 125 -771 131 -374
rect -131 -783 131 -771
<< properties >>
string FIXED_BBOX -254 -902 254 902
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 3.731 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 5.559k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
