magic
tech sky130A
magscale 1 2
timestamp 1750060524
<< metal1 >>
rect 3390 259 3436 365
rect 3508 259 3554 365
rect 3377 199 3383 259
rect 3443 199 3449 259
rect 3495 199 3501 259
rect 3561 199 3567 259
rect 3495 -85 3501 -25
rect 3561 -85 3567 -25
rect 3377 -173 3383 -113
rect 3443 -173 3449 -113
rect 3390 -279 3436 -173
rect 3508 -291 3554 -85
<< via1 >>
rect 3383 199 3443 259
rect 3501 199 3561 259
rect 3501 -85 3561 -25
rect 3383 -173 3443 -113
<< metal2 >>
rect 3119 817 3129 873
rect 3185 817 3195 873
rect 2993 729 3003 785
rect 3059 729 3069 785
rect 3875 641 3885 697
rect 3941 641 3951 697
rect 2936 609 3699 611
rect 2936 553 3633 609
rect 3689 553 3699 609
rect 2936 551 3699 553
rect 3749 465 3759 521
rect 3815 465 3825 521
rect 3245 377 3255 433
rect 3311 377 3321 433
rect 2993 289 3003 345
rect 3059 289 3069 345
rect 3371 257 3383 259
rect 3371 201 3381 257
rect 3371 199 3383 201
rect 3443 199 3449 259
rect 3495 199 3501 259
rect 3561 257 3573 259
rect 3563 201 3573 257
rect 3561 199 3573 201
rect 3375 -27 3501 -25
rect 3371 -83 3381 -27
rect 3437 -83 3501 -27
rect 3375 -85 3501 -83
rect 3561 -85 3567 -25
rect 3377 -173 3383 -113
rect 3443 -115 3573 -113
rect 3443 -171 3507 -115
rect 3563 -171 3573 -115
rect 3443 -173 3573 -171
rect 2993 -259 3003 -203
rect 3059 -259 3069 -203
rect 3245 -347 3255 -291
rect 3311 -347 3321 -291
rect 3749 -435 3759 -379
rect 3815 -435 3825 -379
rect 3624 -467 4006 -465
rect 3624 -523 3633 -467
rect 3689 -523 4006 -467
rect 3624 -525 4006 -523
rect 3875 -611 3885 -555
rect 3941 -611 3951 -555
rect 2993 -699 3003 -643
rect 3059 -699 3069 -643
rect 3119 -787 3129 -731
rect 3185 -787 3195 -731
<< via2 >>
rect 3129 817 3185 873
rect 3003 729 3059 785
rect 3885 641 3941 697
rect 3633 553 3689 609
rect 3759 465 3815 521
rect 3255 377 3311 433
rect 3003 289 3059 345
rect 3381 201 3383 257
rect 3383 201 3437 257
rect 3507 201 3561 257
rect 3561 201 3563 257
rect 3381 -83 3437 -27
rect 3507 -171 3563 -115
rect 3003 -259 3059 -203
rect 3255 -347 3311 -291
rect 3759 -435 3815 -379
rect 3633 -523 3689 -467
rect 3885 -611 3941 -555
rect 3003 -699 3059 -643
rect 3129 -787 3185 -731
<< metal3 >>
rect 2998 785 3064 1071
rect 2998 729 3003 785
rect 3059 729 3064 785
rect 2998 345 3064 729
rect 2998 289 3003 345
rect 3059 289 3064 345
rect 2998 -203 3064 289
rect 2998 -259 3003 -203
rect 3059 -259 3064 -203
rect 2998 -643 3064 -259
rect 2998 -699 3003 -643
rect 3059 -699 3064 -643
rect 2998 -704 3064 -699
rect 3124 873 3190 1071
rect 3124 817 3129 873
rect 3185 817 3190 873
rect 3124 -731 3190 817
rect 3250 433 3316 1071
rect 3250 377 3255 433
rect 3311 377 3316 433
rect 3250 -291 3316 377
rect 3376 257 3442 1071
rect 3376 201 3381 257
rect 3437 201 3442 257
rect 3376 -27 3442 201
rect 3376 -83 3381 -27
rect 3437 -83 3442 -27
rect 3376 -176 3442 -83
rect 3502 257 3568 1071
rect 3502 201 3507 257
rect 3563 201 3568 257
rect 3502 -115 3568 201
rect 3502 -171 3507 -115
rect 3563 -171 3568 -115
rect 3502 -176 3568 -171
rect 3628 609 3694 1071
rect 3628 553 3633 609
rect 3689 553 3694 609
rect 3250 -347 3255 -291
rect 3311 -347 3316 -291
rect 3250 -352 3316 -347
rect 3628 -467 3694 553
rect 3754 521 3820 1071
rect 3754 465 3759 521
rect 3815 465 3820 521
rect 3754 -379 3820 465
rect 3754 -435 3759 -379
rect 3815 -435 3820 -379
rect 3754 -440 3820 -435
rect 3880 697 3946 1071
rect 3880 641 3885 697
rect 3941 641 3946 697
rect 3628 -523 3633 -467
rect 3689 -523 3694 -467
rect 3628 -528 3694 -523
rect 3880 -555 3946 641
rect 3880 -611 3885 -555
rect 3941 -611 3946 -555
rect 3880 -616 3946 -611
rect 3124 -787 3129 -731
rect 3185 -787 3190 -731
rect 3124 -792 3190 -787
use cm_ncell1_half  cm_ncell1_half_0
timestamp 1750060524
transform 1 0 -26 0 1 3
box -12 0 7008 1068
use cm_ncell1_half  cm_ncell1_half_1
timestamp 1750060524
transform -1 0 6970 0 -1 83
box -12 0 7008 1068
<< labels >>
flabel metal3 s 2998 1001 3064 1071 0 FreeSans 320 0 0 0 G1
port 0 nsew
flabel metal3 s 3124 1001 3190 1071 0 FreeSans 320 0 0 0 io0
port 1 nsew
flabel metal3 s 3250 1001 3316 1071 0 FreeSans 320 0 0 0 io1
port 2 nsew
flabel metal3 s 3376 1001 3442 1071 0 FreeSans 320 0 0 0 to0
port 3 nsew
flabel metal3 s 3502 1001 3568 1071 0 FreeSans 320 0 0 0 to1
port 4 nsew
flabel metal3 s 3628 1001 3694 1071 0 FreeSans 320 0 0 0 to2
port 5 nsew
flabel metal3 s 3754 1001 3820 1071 0 FreeSans 320 0 0 0 to3
port 6 nsew
flabel metal3 s 3880 1001 3946 1071 0 FreeSans 320 0 0 0 to4
port 7 nsew
flabel metal1 s 2825 1001 2891 1071 0 FreeSans 320 0 0 0 GND
port 8 nsew
<< end >>
