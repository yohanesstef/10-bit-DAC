magic
tech sky130A
timestamp 1749667264
use sky130_fd_sc_hd__nand2_1  x1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 315 0 1 -980
box -19 -24 157 296
use sky130_fd_sc_hd__nand2_1  x2
timestamp 1704896540
transform 1 0 453 0 1 -980
box -19 -24 157 296
use sky130_fd_sc_hd__nor2_1  x3 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 591 0 1 -980
box -19 -24 157 296
<< end >>
