magic
tech sky130A
magscale 1 2
timestamp 1750900893
<< error_s >>
rect 36386 -4420 36392 -4414
rect 36440 -4420 36446 -4414
rect 36380 -4426 36386 -4420
rect 36446 -4426 36452 -4420
rect 36380 -4480 36386 -4474
rect 36446 -4480 36452 -4474
rect 36386 -4486 36392 -4480
rect 36440 -4486 36446 -4480
rect 36110 -4508 36116 -4502
rect 36164 -4508 36170 -4502
rect 36104 -4514 36110 -4508
rect 36170 -4514 36176 -4508
rect 36104 -4568 36110 -4562
rect 36170 -4568 36176 -4562
rect 36110 -4574 36116 -4568
rect 36164 -4574 36170 -4568
rect 35834 -4596 35840 -4590
rect 35888 -4596 35894 -4590
rect 35828 -4602 35834 -4596
rect 35894 -4602 35900 -4596
rect 35828 -4656 35834 -4650
rect 35894 -4656 35900 -4650
rect 35834 -4662 35840 -4656
rect 35888 -4662 35894 -4656
rect 35568 -4684 35574 -4678
rect 35622 -4684 35628 -4678
rect 35562 -4690 35568 -4684
rect 35628 -4690 35634 -4684
rect 35562 -4744 35568 -4738
rect 35628 -4744 35634 -4738
rect 35568 -4750 35574 -4744
rect 35622 -4750 35628 -4744
rect 35480 -4772 35486 -4766
rect 35534 -4772 35540 -4766
rect 35474 -4778 35480 -4772
rect 35540 -4778 35546 -4772
rect 35474 -4832 35480 -4826
rect 35540 -4832 35546 -4826
rect 35480 -4838 35486 -4832
rect 35534 -4838 35540 -4832
rect 35214 -4860 35220 -4854
rect 35268 -4860 35274 -4854
rect 35208 -4866 35214 -4860
rect 35274 -4866 35280 -4860
rect 35208 -4920 35214 -4914
rect 35274 -4920 35280 -4914
rect 35214 -4926 35220 -4920
rect 35268 -4926 35274 -4920
rect 34938 -4948 34944 -4942
rect 34992 -4948 34998 -4942
rect 34932 -4954 34938 -4948
rect 34998 -4954 35004 -4948
rect 34932 -5008 34938 -5002
rect 34998 -5008 35004 -5002
rect 34938 -5014 34944 -5008
rect 34992 -5014 34998 -5008
rect 34662 -5036 34668 -5030
rect 34716 -5036 34722 -5030
rect 34656 -5042 34662 -5036
rect 34722 -5042 34728 -5036
rect 34656 -5096 34662 -5090
rect 34722 -5096 34728 -5090
rect 34662 -5102 34668 -5096
rect 34716 -5102 34722 -5096
<< metal1 >>
rect 36386 -4420 36446 -4414
rect 36110 -4508 36170 -4502
rect 35834 -4596 35894 -4590
rect 35568 -4684 35628 -4678
rect 35480 -4772 35540 -4766
rect 35214 -4860 35274 -4854
rect 34938 -4948 34998 -4942
rect 34662 -5036 34722 -5030
rect 34291 -5386 34486 -5326
rect 34662 -5386 34722 -5096
rect 34938 -5386 34998 -5008
rect 35214 -5386 35274 -4920
rect 35480 -5187 35540 -4832
rect 35490 -5298 35540 -5187
rect 35480 -5386 35540 -5298
rect 35568 -5187 35628 -4744
rect 35568 -5298 35618 -5187
rect 35568 -5386 35628 -5298
rect 35834 -5386 35894 -4656
rect 36110 -5386 36170 -4568
rect 36386 -5386 36446 -4480
rect 36622 -5386 36817 -5326
rect 34755 -5414 34815 -5386
rect 34291 -5474 34815 -5414
rect 35031 -5502 35091 -5386
rect 34291 -5562 35091 -5502
rect 35307 -5590 35367 -5386
rect 34291 -5650 35367 -5590
rect 35741 -5590 35801 -5386
rect 36017 -5502 36077 -5386
rect 36293 -5414 36353 -5386
rect 36293 -5474 36817 -5414
rect 36017 -5562 36817 -5502
rect 35741 -5650 36817 -5590
<< via1 >>
rect 36386 -4480 36446 -4420
rect 36110 -4568 36170 -4508
rect 35834 -4656 35894 -4596
rect 35568 -4744 35628 -4684
rect 35480 -4832 35540 -4772
rect 35214 -4920 35274 -4860
rect 34938 -5008 34998 -4948
rect 34662 -5096 34722 -5036
use hnmos_8  hnmos_8_8
timestamp 1750900893
transform 1 0 34447 0 1 -5402
box -137 -180 2351 358
<< end >>
