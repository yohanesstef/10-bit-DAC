magic
tech sky130A
magscale 1 2
timestamp 1749057406
<< pwell >>
rect -307 -1042 307 1042
<< psubdiff >>
rect -271 972 -175 1006
rect 175 972 271 1006
rect -271 910 -237 972
rect 237 910 271 972
rect -271 -972 -237 -910
rect 237 -972 271 -910
rect -271 -1006 -175 -972
rect 175 -1006 271 -972
<< psubdiffcont >>
rect -175 972 175 1006
rect -271 -910 -237 910
rect 237 -910 271 910
rect -175 -1006 175 -972
<< xpolycontact >>
rect -141 444 141 876
rect -141 -876 141 -444
<< xpolyres >>
rect -141 -444 141 444
<< locali >>
rect -271 972 -175 1006
rect 175 972 271 1006
rect -271 910 -237 972
rect 237 910 271 972
rect -271 -972 -237 -910
rect 237 -972 271 -910
rect -271 -1006 -175 -972
rect 175 -1006 271 -972
<< viali >>
rect -125 461 125 858
rect -125 -858 125 -461
<< metal1 >>
rect -131 858 131 870
rect -131 461 -125 858
rect 125 461 131 858
rect -131 449 131 461
rect -131 -461 131 -449
rect -131 -858 -125 -461
rect 125 -858 131 -461
rect -131 -870 131 -858
<< properties >>
string FIXED_BBOX -254 -989 254 989
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 4.603 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 6.796k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
