magic
tech sky130A
magscale 1 2
timestamp 1749017082
<< metal1 >>
rect 19701 -21505 19761 -21181
rect 19678 -21767 19761 -21505
rect 19257 -21829 19761 -21767
rect 19789 -22153 19849 -21181
rect 19678 -22415 19849 -22153
rect 19257 -22477 19849 -22415
rect 19877 -22801 19937 -21181
rect 19678 -23063 19937 -22801
rect 19257 -23125 19937 -23063
use rseg_1_pin_4  rseg_1_pin_4_0 ~/10-bit-DAC/mag
timestamp 1748967404
transform 1 0 18073 0 1 1583
box 1540 -22764 1864 -22364
<< end >>
