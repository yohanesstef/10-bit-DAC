magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< xpolycontact >>
rect -141 234 141 666
rect -141 -666 141 -234
<< xpolyres >>
rect -141 -234 141 234
<< viali >>
rect -125 251 125 648
rect -125 -648 125 -251
<< metal1 >>
rect -131 648 131 660
rect -131 251 -125 648
rect 125 251 131 648
rect -131 239 131 251
rect -131 -251 131 -239
rect -131 -648 -125 -251
rect 125 -648 131 -251
rect -131 -660 131 -648
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 2.501 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 3.814k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
