* PEX produced on Sat Jun 28 04:59:43 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from DAC_10b_top.ext - technology: sky130A

.subckt DAC_10b_posim_top DIN0 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 DIN9 ROUT1 ROUT2
+ VDD VDDH GND VOUT
X0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t4 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_45343_4538.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t4 GND.t178 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t6 top_DAC_0/top_final_switch_0.VOUT[1].t4 a_6778_12595.t3 GND.t418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 GND.t970 GND.t971 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t2 a_30056_7686.t3 GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X5 GND.t360 GND.t358 GND.t359 GND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X6 a_44062_19517.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t0 GND.t913 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t2 a_14331_6250.t3 VDDH.t491 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X8 a_21927_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t2 a_23629_18133.t0 GND.t901 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.t1 GND.t167 sky130_fd_pr__res_xhigh_po_1p41 l=10.24
X10 a_44234_9966.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t0 GND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t22 GND.t29 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X12 a_44234_17252.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t4 GND.t740 GND.t504 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t22 VDDH.t571 VDDH.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X14 GND.t379 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t1 GND.t378 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_45023_21964.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t4 GND.t372 GND.t371 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 GND.t357 GND.t355 GND.t356 GND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X17 VDDH.t572 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t7 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t4 a_43167_4358.t0 GND.t937 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t24 VDDH.t507 VDDH.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X20 GND.t820 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t3 GND.t819 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t2 GND.t387 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X22 VDDH.t508 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t18 VDDH.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X23 VDD.t120 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t3 VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X24 a_14615_13536.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t2 top_DAC_0/top_rseg_n_dcell_0.VH2.t2 GND.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X25 a_20656_10031.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t2 a_19946_8950.t1 VDDH.t378 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X26 a_43698_8776.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t2 a_43724_9372.t1 VDDH.t515 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X27 a_23307_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t2 a_22193_18133.t1 GND.t403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X28 a_14948_18696.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t2 a_14790_18696.t0 VDDH.t493 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t24 VOUT.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t4 a_43167_3162.t1 GND.t955 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t0 DIN2.t0 VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 GND.t353 GND.t354 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t7 VDDH.t345 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.t1 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t2 GND.t41 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X36 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t2 a_43240_20580.t1 VDDH.t382 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X37 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t2 a_23307_20174.t3 GND.t591 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X38 GND.t423 GND.t424 GND.t167 sky130_fd_pr__res_xhigh_po_1p41 l=11.57
X39 GND.t31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t32 GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X40 a_6923_9707.t23 VOUT.t48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t19 GND.t813 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X41 VDDH.t469 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t6 a_43724_8936.t1 VDDH.t468 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X42 a_18284_18696.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t2 a_15618_18696.t0 VDDH.t405 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X43 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33.t2 GND.t22 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X44 a_31042_7686.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28.t0 GND.t527 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X45 a_36888_19550.t3 a_36888_19786.t6 GND.t700 GND.t698 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X46 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t5 VDD.t218 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X47 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31.t2 GND.t60 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X48 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t2 a_24963_20174.t3 GND.t737 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t20 top_DAC_0/top_final_switch_0.VOUT[0].t4 a_5050_12595.t3 GND.t887 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X50 a_43698_14716.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t2 a_43724_15312.t0 VDDH.t351 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.t0 GND.t57 sky130_fd_pr__res_xhigh_po_1p41 l=1.99
X52 VDDH.t509 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t6 VDDH.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X53 a_6923_9707.t11 top_DAC_0/top_final_switch_0.VOUT[4].t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t16 GND.t813 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t24 GND.t33 GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X55 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t3 a_21927_20174.t3 GND.t787 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X56 VDDH.t510 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t3 VDDH.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t2 a_29780_7686.t1 GND.t928 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X58 a_31870_7686.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31.t1 GND.t528 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X59 top_DAC_0/top_final_switch_0.VOUT[1].t3 top_DAC_0/top_rseg_n_dcell_0.SH[3].t2 top_DAC_0/top_rseg_n_dcell_0.VL3.t2 VDDH.t562 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X60 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38.t0 GND.t364 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X61 VDD.t211 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t4 VDD.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t28 VDDH.t511 VDDH.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X63 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t3 a_44255_4614.t0 GND.t954 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X64 a_23629_18133.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t4 top_DAC_0/top_rseg_n_dcell_0.VL2.t1 GND.t529 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X65 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4.t0 GND.t368 sky130_fd_pr__res_xhigh_po_1p41 l=3.37
X66 VDD.t220 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t2 VDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t23 VOUT.t49 a_5050_12595.t9 GND.t887 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t23 GND.t539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.087 pd=0.89 as=0.174 ps=1.78 w=0.6 l=20
X69 a_14615_14034.t1 top_DAC_0/top_rseg_n_dcell_0.SH[2].t2 top_DAC_0/top_final_switch_0.VOUT[3].t0 GND.t496 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X70 a_20932_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t2 a_18724_8950.t1 VDDH.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X71 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t4 a_45023_18840.t0 GND.t155 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X72 a_24135_20174.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t3 a_23629_18133.t5 GND.t404 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X73 a_15098_19866.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t3 a_15618_18696.t1 VDDH.t494 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X74 a_43167_4358.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t5 GND.t822 GND.t821 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X75 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.t0 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=4.81
X76 VDDH.t237 VDDH.t235 VDDH.t236 VDDH.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X77 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t4 a_43391_3326.t0 GND.t140 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t22 VDDH.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X79 VDDH.t234 VDDH.t232 VDDH.t233 VDDH.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X80 GND.t35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t3 GND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X81 a_42982_21320.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t2 a_42724_21320.t1 VDDH.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X82 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t29 VDDH.t512 VDDH.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X83 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t4 a_24135_20174.t1 GND.t788 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X84 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t2 GND.t889 GND.t888 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X85 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t5 VDD.t122 VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X86 VDDH.t231 VDDH.t229 VDDH.t230 VDDH.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X87 VDDH.t513 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t18 VDDH.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X88 GND.t352 GND.t350 GND.t351 GND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X89 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t9 GND.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X90 VDDH.t313 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t17 VDDH.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X91 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t4 VDD.t164 VDD.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X92 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t26 GND.t37 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X93 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t2 VDDH.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X94 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60.t0 GND.t81 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X95 a_15224_18696.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.t0 VDDH.t498 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X96 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t3 DIN1.t0 VDD.t52 VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X97 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t28 VOUT.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 a_44234_11946.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t1 GND.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X99 GND.t348 GND.t349 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 GND.t734 DIN2.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t1 GND.t733 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X101 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t0 GND.t18 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X102 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t2 a_15629_7686.t4 VDDH.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X103 a_31594_7686.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30.t1 GND.t530 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X104 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47.t1 GND.t80 sky130_fd_pr__res_xhigh_po_1p41 l=6.09
X105 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t4 a_44255_3438.t0 GND.t547 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X106 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t5 a_44479_3254.t0 GND.t141 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X107 a_43698_9766.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t8 a_44234_10322.t1 GND.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X108 a_14514_18696.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t2 a_17148_18696.t2 VDDH.t440 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X109 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15.t0 GND.t79 sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X110 GND.t935 DIN5.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t3 GND.t934 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X111 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t32 VDDH.t314 VDDH.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X112 top_DAC_0/top_rseg_n_dcell_0.VL2.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t3 a_14615_14034.t2 GND.t487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X113 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t18 VDDH.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X114 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.t2 GND.t79 sky130_fd_pr__res_xhigh_po_1p41 l=4.45
X115 VDDH.t315 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t7 VDDH.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X116 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t1 a_38672_20477.t1 GND.t799 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X117 GND.t898 GND.t899 GND.t19 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X118 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t3 a_21375_20174.t2 GND.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X119 GND.t441 DIN8.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t0 GND.t440 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X120 VDDH.t316 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t6 VDDH.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X121 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t25 VOUT.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 a_16615_7686.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t2 VDDH.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X123 VDDH.t471 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t7 a_43724_15866.t1 VDDH.t470 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X124 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t35 VDDH.t317 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X125 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t36 VDDH.t318 VDDH.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X126 a_45023_21136.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t2 GND.t386 GND.t385 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X127 GND.t346 GND.t347 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t4 GND.t518 GND.t517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X129 GND.t344 GND.t345 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 a_33634_8950.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t2 a_27620_6250.t3 GND.t463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X131 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28.t2 GND.t9 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X132 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t4 GND.t523 GND.t522 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X133 a_24687_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t3 a_23629_18133.t3 GND.t571 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X134 VDDH.t228 VDDH.t226 VDDH.t227 VDDH.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X135 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t2 GND.t18 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X136 a_43391_3878.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t5 a_43391_3794.t0 GND.t862 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X137 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t29 VOUT.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t2 VDDH.t529 VDDH.t528 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X139 VDDH.t319 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t5 VDDH.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X140 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t23 VDDH.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X141 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t2 GND.t54 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X142 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t27 GND.t62 GND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X143 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t7 VOUT.t50 a_8506_12595.t11 GND.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X144 a_28606_6250.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t3 a_34304_8950.t2 GND.t464 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X145 a_5111_10963.t3 a_5111_10963.t2 GND.t927 GND.t462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.464 ps=3.78 w=1.6 l=1
X146 GND.t762 GND.t763 GND.t9 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X147 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t24 VDDH.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X148 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t22 VOUT.t51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t8 VDDH.t337 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X149 GND.t342 GND.t343 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t16 VDDH.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X151 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t8 VDDH.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X152 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t28 GND.t64 GND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X153 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13.t0 GND.t38 sky130_fd_pr__res_xhigh_po_1p41 l=5.58
X154 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34.t2 GND.t364 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X155 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t13 top_DAC_0/top_final_switch_0.VOUT[1].t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t3 VDDH.t337 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X156 a_42724_21320.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t6 VDDH.t367 VDDH.t365 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X157 GND.t341 GND.t338 GND.t340 GND.t339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X158 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t1 GND.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X159 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t5 a_23859_20174.t1 GND.t789 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X160 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t0 top_DAC_0/top_final_switch_0.VOUT[2].t4 a_8506_12595.t0 GND.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X161 GND.t572 GND.t573 GND.t60 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X162 a_29434_6250.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t4 a_35132_8950.t2 GND.t465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X163 GND.t964 GND.t965 GND.t167 sky130_fd_pr__res_xhigh_po_1p41 l=6.65
X164 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t20 GND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X165 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t6 GND.t427 GND.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X166 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t3 VDD.t92 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X167 a_43240_22004.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t3 a_42982_22004.t1 VDDH.t252 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X168 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t6 a_44255_3714.t0 GND.t863 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X169 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t4 GND.t510 GND.t509 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X170 a_35453_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t3 a_34856_8950.t0 GND.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X171 GND.t838 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t1 GND.t837 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X172 a_15374_19866.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.t0 VDDH.t499 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X173 VDDH.t225 VDDH.t223 VDDH.t224 VDDH.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X174 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t2 a_30608_7686.t4 GND.t771 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X175 VDDH.t285 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t0 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X176 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t26 VOUT.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 a_44062_18449.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t0 GND.t835 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X178 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t38 VDDH.t261 VDDH.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X179 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t5 GND.t381 GND.t380 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X180 GND.t482 DIN1.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t1 GND.t481 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X181 VDD.t35 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X182 GND.t40 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 a_44062_18093.t1 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X183 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t0 DIN5.t1 GND.t891 GND.t890 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X184 GND.t337 GND.t335 GND.t336 GND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X185 VDDH.t222 VDDH.t220 VDDH.t221 VDDH.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X186 VDDH.t546 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t6 VOUT.t38 VDDH.t545 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X187 a_15066_18696.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t3 a_16596_18696.t2 VDDH.t441 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X188 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t2 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X189 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t1 DIN8.t1 GND.t538 GND.t537 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X190 a_14615_14283.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t2 top_DAC_0/top_rseg_n_dcell_0.VH2.t1 GND.t457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X191 GND.t329 GND.t330 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 GND.t334 GND.t331 GND.t333 GND.t332 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X193 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t0 GND.t88 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X194 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t4 a_20823_20174.t3 GND.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X195 GND.t328 GND.t326 GND.t327 GND.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X196 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t30 VOUT.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 GND.t66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t30 GND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X198 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t3 a_14055_6250.t3 VDDH.t490 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X199 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t39 VDDH.t263 VDDH.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X200 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2.t0 GND.t368 sky130_fd_pr__res_xhigh_po_1p41 l=4.24
X201 GND.t428 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t10 GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X202 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t2 GND.t41 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X203 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t15 VDDH.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X204 a_43240_18130.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t3 a_42982_18130.t1 VDDH.t417 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X205 a_43240_19896.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t4 a_42982_19896.t1 VDDH.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X206 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t7 VDDH.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X207 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t2 GND.t88 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X208 GND.t68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t15 GND.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X209 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t4 GND.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X210 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t15 VDDH.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X211 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.t2 GND.t365 sky130_fd_pr__res_xhigh_po_1p41 l=3.58
X212 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58.t0 GND.t81 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X213 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t36 GND.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X214 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t6 a_24687_20174.t0 GND.t790 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X215 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15.t2 GND.t38 sky130_fd_pr__res_xhigh_po_1p41 l=5.32
X216 GND.t324 GND.t325 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 VDDH.t219 VDDH.t217 VDDH.t218 VDDH.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X218 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t23 VOUT.t52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t27 VDDH.t542 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X219 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t27 VDDH.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X220 a_8506_12595.t1 top_DAC_0/top_final_switch_0.VOUT[2].t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t1 GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X221 a_14672_18696.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4.t1 VDDH.t500 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X222 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t6 VDD.t36 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X223 a_35757_10031.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t5 a_33634_8950.t0 GND.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X224 a_43724_12342.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t8 VDDH.t473 VDDH.t472 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X225 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t19 top_DAC_0/top_final_switch_0.VOUT[4].t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t27 VDDH.t542 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X226 VDD.t107 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t2 VDD.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X227 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t5 top_DAC_0/top_final_switch_0.VOUT[1].t6 a_6778_12595.t2 GND.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X228 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t4 VDDH.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X229 VDDH.t264 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t16 VDDH.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X230 GND.t323 GND.t321 GND.t322 GND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X231 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t17 top_DAC_0/top_final_switch_0.VOUT[0].t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t3 VDDH.t559 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X232 VDD.t50 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t2 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X233 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.t0 GND.t368 sky130_fd_pr__res_xhigh_po_1p41 l=2.5
X234 a_8506_12595.t10 VOUT.t53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t6 GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X235 VDDH.t216 VDDH.t214 VDDH.t215 VDDH.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X236 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t2 GND.t669 GND.t668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X237 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t1 GND.t54 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X238 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50.t1 GND.t361 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X239 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t8 GND.t92 GND.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X240 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t11 VOUT.t54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t9 VDDH.t559 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X241 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t37 GND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X242 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t3 a_43240_18814.t1 VDDH.t425 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X243 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t15 VOUT.t55 a_6778_12595.t7 GND.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X244 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t5 a_21651_20174.t2 GND.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X245 a_42847_4906.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t1 VDD.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X246 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t3 VDD.t103 VDD.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X247 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t13 VDDH.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X248 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t3 a_30332_7686.t2 GND.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X249 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t1 GND.t387 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X250 GND.t639 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t4 a_44234_14916.t0 GND.t638 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X251 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t4 VDD.t79 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X252 a_45023_18840.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t5 GND.t641 GND.t640 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X253 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t1 GND.t540 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.087 ps=0.89 w=0.6 l=20
X254 a_44234_15906.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t1 GND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X255 VDDH.t381 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t0 VDDH.t380 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X256 a_28882_6250.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53.t0 GND.t929 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X257 GND.t21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 a_44062_21653.t1 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X258 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45.t2 GND.t80 sky130_fd_pr__res_xhigh_po_1p41 l=5.88
X259 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t2 a_39936_22083.t2 VDDH.t466 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=1
X260 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t41 VDDH.t265 VDDH.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X261 a_8051_10107.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t7 GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X262 a_43698_13726.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t10 a_44234_14282.t0 GND.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X263 a_29434_6250.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55.t0 GND.t930 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X264 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33.t1 GND.t22 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X265 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44.t2 GND.t13 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X266 GND.t320 GND.t318 GND.t319 GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X267 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t14 VDDH.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X268 a_19468_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t3 top_DAC_0/top_rseg_n_dcell_0.VS4.t1 VDDH.t530 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X269 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t27 VOUT.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 a_15863_13287.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t4 top_DAC_0/top_rseg_n_dcell_0.VH3.t1 VDDH.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X271 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t5 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X272 GND.t286 GND.t287 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 top_DAC_0/top_rseg_n_dcell_0.VS4.t3 top_DAC_0/top_rseg_n_dcell_0.SH[4].t2 top_DAC_0/top_final_switch_0.VOUT[0].t2 VDDH.t419 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X274 a_16872_18696.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1.t1 VDDH.t501 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X275 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t6 GND.t59 GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X276 GND.t442 GND.t443 GND.t361 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X277 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26.t0 GND.t9 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X278 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t7 a_30332_7686.t0 GND.t606 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X279 GND.t775 GND.t776 GND.t79 sky130_fd_pr__res_xhigh_po_1p41 l=3.94
X280 a_28882_6250.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37.t2 GND.t766 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X281 VDD.t19 DIN9.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t0 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X282 GND.t69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t29 GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X283 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t9 GND.t94 GND.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X284 top_DAC_0/top_final_switch_0.VOUT[4].t0 top_DAC_0/top_rseg_n_dcell_0.SH[1].t2 top_DAC_0/top_rseg_n_dcell_0.VS1.t6 GND.t454 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X285 a_39306_20477.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t11 GND.t146 GND.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=5.3
X286 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t6 VDDH.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X287 GND.t479 GND.t480 GND.t54 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X288 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t3 VDDH.t407 VDDH.t406 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X289 a_19946_8950.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t5 a_16891_7686.t0 VDDH.t448 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X290 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t11 a_6923_9707.t15 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X291 a_43724_12896.t1 a_43698_12736.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t1 VDDH.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X292 a_17732_18696.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t2 a_14514_18696.t1 VDDH.t395 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X293 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47.t2 GND.t693 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X294 a_28882_6250.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21.t2 GND.t607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X295 GND.t362 GND.t363 GND.t361 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X296 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t4 a_15353_7686.t3 VDDH.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X297 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t2 VDDH.t329 VDDH.t328 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X298 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t4 a_22203_20174.t3 GND.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X299 GND.t609 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t1 GND.t608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X300 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3.t2 GND.t365 sky130_fd_pr__res_xhigh_po_1p41 l=3.32
X301 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38.t2 GND.t364 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X302 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t5 VDD.t89 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X303 GND.t507 a_5111_10963.t0 a_5111_10963.t1 GND.t506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.232 ps=1.89 w=1.6 l=1
X304 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t12 a_6923_9707.t16 GND.t419 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X305 GND.t70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t28 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X306 a_33358_8950.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t6 a_27344_6250.t3 GND.t642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X307 VDD.t68 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 VDD.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X308 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t5 a_20823_20174.t4 GND.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X309 GND.t962 GND.t963 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X310 GND.t96 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t0 GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X311 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t5 VDDH.t273 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X312 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t5 VDD.t186 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X313 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t23 VOUT.t56 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t11 VDDH.t539 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X314 a_8473_23194.t2 ROUT1.t0 ROUT1.t1 VDDH.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X315 a_20076_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t4 a_19552_8950.t0 VDDH.t250 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X316 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t13 a_8051_10107.t10 GND.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X317 a_6923_9707.t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t26 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X318 GND.t664 GND.t665 GND.t57 sky130_fd_pr__res_xhigh_po_1p41 l=1.68
X319 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t6 VDDH.t272 VDDH.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X320 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t12 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t4 VDDH.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X321 a_44234_6996.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t0 GND.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X322 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t19 top_DAC_0/top_final_switch_0.VOUT[2].t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t7 VDDH.t539 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X323 a_8051_10107.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t5 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X324 a_44234_14282.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t4 GND.t897 GND.t896 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X325 a_34186_8950.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t7 a_28172_6250.t3 GND.t643 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X326 GND.t807 GND.t808 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X327 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t31 VOUT.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t15 VDDH.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X329 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t32 VOUT.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 VDDH.t346 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t3 VDDH.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X331 VDDH.t213 VDDH.t211 VDDH.t212 VDDH.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X332 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t6 a_23583_20174.t2 GND.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X333 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.t2 GND.t38 sky130_fd_pr__res_xhigh_po_1p41 l=5.73
X334 a_45343_4622.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t6 a_45343_4538.t1 GND.t938 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X335 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t2 a_43240_20238.t1 VDDH.t382 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X336 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t38 VDDH.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X337 VDDH.t210 VDDH.t208 VDDH.t209 VDDH.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X338 VDDH.t267 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t15 VDDH.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X339 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22.t1 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X340 a_45023_20264.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t6 GND.t824 GND.t823 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X341 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45.t1 GND.t80 sky130_fd_pr__res_xhigh_po_1p41 l=5.73
X342 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t6 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X343 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t11 GND.t97 GND.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X344 GND.t284 GND.t285 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 GND.t72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t27 GND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X346 a_43724_9926.t0 a_43698_9766.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t1 VDDH.t497 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X347 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t5 a_30332_7686.t4 GND.t767 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X348 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32.t1 GND.t364 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X349 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t28 VOUT.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 GND.t282 GND.t283 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 GND.t574 GND.t575 GND.t18 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X352 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t0 GND.t387 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X353 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t7 a_22203_20174.t2 GND.t165 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X354 GND.t921 GND.t922 GND.t60 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X355 a_23049_18133.t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t6 top_DAC_0/top_rseg_n_dcell_0.VL2.t8 GND.t768 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X356 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t6 a_21651_20174.t3 GND.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X357 a_43724_16302.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t9 VDDH.t427 VDDH.t426 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X358 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.t0 GND.t38 sky130_fd_pr__res_xhigh_po_1p41 l=6.14
X359 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t4 VDDH.t273 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X360 VDDH.t207 VDDH.t205 VDDH.t206 VDDH.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X361 VDDH.t204 VDDH.t202 VDDH.t203 VDDH.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X362 a_14615_13536.t0 top_DAC_0/top_rseg_n_dcell_0.SH[2].t3 top_DAC_0/top_final_switch_0.VOUT[1].t0 GND.t497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X363 GND.t923 GND.t924 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X364 VDDH.t201 VDDH.t199 VDDH.t200 VDDH.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X365 a_20656_10031.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t2 a_19468_10031.t2 VDDH.t522 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X366 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t7 a_45343_3530.t0 GND.t864 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X367 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t1 GND.t54 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X368 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t17 GND.t416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X369 top_DAC_0/top_rseg_n_dcell_0.VH3.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t8 a_18284_18696.t2 VDDH.t449 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X370 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t2 top_DAC_0/top_final_switch_0.VOUT[3].t4 a_8051_10107.t3 GND.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X371 GND.t280 GND.t281 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t6 VDD.t188 VDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X373 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t8 a_24411_20174.t2 GND.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X374 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t14 top_DAC_0/top_final_switch_0.VOUT[2].t7 a_8506_12595.t6 GND.t801 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X375 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t6 top_DAC_0/top_final_switch_0.VOUT[2].t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t20 VDDH.t540 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X376 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t10 VOUT.t57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t14 VDDH.t540 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X377 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t14 top_DAC_0/top_final_switch_0.VOUT[1].t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t2 VDDH.t336 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X378 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t43 VDDH.t269 VDDH.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X379 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t7 a_45343_4622.t0 GND.t825 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X380 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t11 VOUT.t58 a_8051_10107.t15 GND.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X381 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t34 GND.t74 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X382 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t12 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t0 GND.t501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X383 a_43240_21320.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t7 a_42982_21320.t0 VDDH.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X384 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t21 VOUT.t59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t7 VDDH.t336 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X385 a_38672_20477.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t4 GND.t367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X386 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t6 VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t29 VOUT.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t5 VOUT.t60 a_8506_12595.t9 GND.t801 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X389 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58.t2 GND.t81 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X390 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t9 a_23031_20174.t2 GND.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X391 top_DAC_0/top_rseg_n_dcell_0.SH[3].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t3 GND.t720 GND.t719 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X392 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t3 VDDH.t345 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X393 GND.t313 GND.t314 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t33 VOUT.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 GND.t886 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t2 GND.t885 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X396 top_DAC_0/top_rseg_n_dcell_0.VS4.t4 top_DAC_0/top_rseg_n_dcell_0.SH[4].t3 top_DAC_0/top_final_switch_0.VOUT[3].t3 VDDH.t419 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X397 a_34569_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t3 top_DAC_0/top_rseg_n_dcell_0.VS1.t0 GND.t415 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X398 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t2 VDDH.t1 VDDH.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X399 a_45023_19712.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t8 GND.t827 GND.t826 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X400 a_39306_20477.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t5 GND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X401 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26.t2 GND.t9 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X402 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t3 VDD.t56 VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X403 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t34 VOUT.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 top_DAC_0/top_rseg_n_dcell_0.SH[1].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t2 VDDH.t333 VDDH.t332 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X405 VDDH.t429 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t10 a_43724_12896.t0 VDDH.t428 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X406 a_28606_6250.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4.t1 GND.t828 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X407 GND.t11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t2 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X408 a_6778_12595.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t1 GND.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X409 GND.t311 GND.t312 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.t2 GND.t79 sky130_fd_pr__res_xhigh_po_1p41 l=4.09
X411 VDD.t181 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t2 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X412 GND.t947 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t26 GND.t468 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X413 a_44234_9332.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t4 GND.t959 GND.t958 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X414 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t44 VDDH.t270 VDDH.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X415 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t17 a_4415_23194.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t2 VDDH.t457 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X416 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t6 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X417 a_6923_9707.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t24 GND.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X418 a_28606_6250.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t7 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36.t2 GND.t769 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X419 a_29434_6250.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7.t2 GND.t570 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X420 VDD.t86 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t2 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X421 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t4 VDDH.t251 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X422 a_22469_18133.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t6 top_DAC_0/top_rseg_n_dcell_0.VL2.t4 GND.t931 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X423 VDDH.t564 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t11 VDDH.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X424 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34.t0 GND.t364 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X425 GND.t948 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t25 GND.t471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X426 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t8 a_20547_20174.t0 GND.t791 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X427 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.t1 GND.t60 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X428 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t3 a_45023_21136.t0 GND.t563 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X429 a_15374_19866.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15.t1 VDDH.t397 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X430 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.t0 GND.t167 sky130_fd_pr__res_xhigh_po_1p41 l=6.65
X431 VDDH.t565 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t14 VDDH.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X432 VDDH.t347 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t2 VDDH.t251 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X433 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t1 GND.t41 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X434 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t10 a_30056_7686.t1 GND.t610 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X435 a_28606_6250.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.t2 GND.t611 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X436 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t6 VDD.t166 VDD.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X437 a_36033_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t5 a_34304_8950.t0 GND.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X438 GND.t309 GND.t310 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1.t2 GND.t772 GND.t368 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X440 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t15 GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X441 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t11 VDDH.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X442 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t47 VDDH.t566 VDDH.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X443 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t6 a_43167_4634.t1 GND.t615 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X444 a_43698_8776.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t13 a_44234_9332.t1 GND.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X445 VDDH.t198 VDDH.t196 VDDH.t197 VDDH.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X446 VDDH.t195 VDDH.t193 VDDH.t194 VDDH.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X447 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t7 a_28172_6250.t1 GND.t625 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X448 a_14615_13785.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t3 top_DAC_0/top_rseg_n_dcell_0.VH2.t5 GND.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X449 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19.t1 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=4.96
X450 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t7 VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X451 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t37 GND.t949 GND.t473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X452 a_29434_6250.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t12 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23.t0 GND.t612 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X453 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t8 a_27344_6250.t4 GND.t770 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X454 a_45023_19988.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t7 GND.t577 GND.t576 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X455 top_DAC_0/top_rseg_n_dcell_0.VL2.t7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t5 a_14615_13536.t2 GND.t487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X456 a_15869_6250.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t3 a_20498_8950.t1 VDDH.t342 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X457 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t4 GND.t671 GND.t670 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t30 VOUT.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.t2 GND.t365 sky130_fd_pr__res_xhigh_po_1p41 l=3.68
X460 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t48 VDDH.t567 VDDH.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X461 a_29158_6250.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54.t0 GND.t626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X462 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.t1 GND.t9 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X463 VDDH.t431 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t11 a_43724_6956.t1 VDDH.t430 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X464 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t1 GND.t88 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X465 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2.t1 GND.t368 sky130_fd_pr__res_xhigh_po_1p41 l=3.73
X466 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6.t1 GND.t368 sky130_fd_pr__res_xhigh_po_1p41 l=2.86
X467 VDDH.t568 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t10 VDDH.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X468 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t11 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t10 a_5111_10963.t5 GND.t506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.232 ps=1.89 w=1.6 l=1
X469 VDDH.t192 VDDH.t190 VDDH.t191 VDDH.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X470 a_16615_7686.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t1 VDDH.t489 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X471 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t50 VDDH.t569 VDDH.t273 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X472 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t9 a_28172_6250.t4 GND.t634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X473 VDDH.t433 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t12 a_43724_9926.t1 VDDH.t432 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X474 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t10 a_24963_20174.t1 GND.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X475 VDD.t206 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X476 a_36888_19550.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t0 GND.t515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X477 GND.t545 GND.t546 GND.t38 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X478 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50.t2 GND.t361 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X479 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t7 VDD.t66 VDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X480 VDD.t11 DIN6.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t2 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X481 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t7 a_24411_20174.t3 GND.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X482 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t1 GND.t88 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X483 a_36033_10031.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t2 a_34873_10031.t1 GND.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X484 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t1 DIN4.t0 VDD.t215 VDD.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X485 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t13 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t1 GND.t501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X486 GND.t617 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t0 GND.t616 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X487 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t9 a_21375_20174.t0 GND.t792 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X488 a_43698_15706.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t3 a_43724_16302.t0 VDDH.t459 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X489 a_17443_7686.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t2 VDDH.t488 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X490 a_44062_20941.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t0 GND.t912 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X491 a_29158_6250.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38.t1 GND.t635 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X492 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t10 a_43240_22004.t0 VDDH.t538 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X493 VDDH.t570 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t9 VDDH.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X494 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t3 DIN7.t0 VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X495 a_35177_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t6 a_35132_8950.t0 GND.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X496 VDDH.t271 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t5 VDDH.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X497 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t7 a_45023_21412.t0 GND.t524 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X498 GND.t411 GND.t412 GND.t54 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X499 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t7 VDD.t31 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X500 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t1 DIN9.t1 GND.t512 GND.t511 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X501 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t36 VDDH.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X502 VDDH.t299 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t8 VDDH.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X503 GND.t966 GND.t967 GND.t364 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X504 a_20222_8950.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t9 a_17167_7686.t1 VDDH.t450 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X505 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t8 a_23031_20174.t3 GND.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X506 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t53 VDDH.t300 VDDH.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X507 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t3 GND.t724 GND.t723 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X508 a_24411_20174.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t4 a_22469_18133.t0 GND.t707 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X509 a_15224_18696.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t4 a_15066_18696.t1 VDDH.t495 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X510 a_45343_3530.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t7 GND.t957 GND.t956 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X511 a_17732_18696.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t4 a_15066_18696.t0 VDDH.t408 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X512 a_23629_18133.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t6 top_DAC_0/top_rseg_n_dcell_0.VH2.t4 GND.t914 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X513 top_DAC_0/top_rseg_n_dcell_0.VL3.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t7 a_15863_13785.t0 VDDH.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X514 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18.t1 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X515 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t17 top_DAC_0/top_final_switch_0.VOUT[4].t6 a_6923_9707.t12 GND.t814 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X516 a_42982_19156.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t7 a_42724_19156.t1 VDDH.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X517 GND.t701 a_36888_19786.t7 a_36888_19550.t2 GND.t493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X518 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t3 GND.t421 GND.t420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X519 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t1 GND.t19 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X520 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t3 top_DAC_0/top_final_switch_0.VOUT[3].t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t3 VDDH.t245 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X521 GND.t99 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t2 GND.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X522 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t9 a_43240_18130.t0 VDDH.t425 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X523 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t20 VDDH.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X524 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t3 VDD.t123 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X525 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t3 a_43240_19896.t0 VDDH.t382 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X526 top_DAC_0/top_rseg_n_dcell_0.SH[4].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t2 VDDH.t574 VDDH.t573 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X527 GND.t870 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t4 a_44234_11946.t0 GND.t869 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X528 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t18 VOUT.t61 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t15 VDDH.t245 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X529 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t21 top_DAC_0/top_final_switch_0.VOUT[2].t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t5 VDDH.t541 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X530 VDD.t85 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 VDD.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X531 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t18 VOUT.t62 a_6923_9707.t22 GND.t814 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X532 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t3 VDD.t202 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X533 a_44234_12936.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t0 GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X534 GND.t854 GND.t855 GND.t22 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X535 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t11 a_22203_20174.t0 GND.t782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X536 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t13 VOUT.t63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t9 VDDH.t541 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X537 GND.t317 GND.t315 GND.t316 GND.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X538 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t38 GND.t950 GND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X539 a_17148_18696.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t3 VDDH.t398 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X540 GND.t760 GND.t761 GND.t57 sky130_fd_pr__res_xhigh_po_1p41 l=2.35
X541 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t28 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t7 VDDH.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X542 GND.t951 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t13 GND.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X543 a_43698_10756.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t15 a_44234_11312.t1 GND.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X544 top_DAC_0/top_final_switch_0.VOUT[2].t1 top_DAC_0/top_rseg_n_dcell_0.SH[1].t3 top_DAC_0/top_rseg_n_dcell_0.VS1.t5 GND.t455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X545 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t2 GND.t54 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X546 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t54 VDDH.t302 VDDH.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X547 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t55 VDDH.t303 VDDH.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X548 GND.t308 GND.t306 GND.t307 GND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X549 a_5050_12595.t2 top_DAC_0/top_final_switch_0.VOUT[0].t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t21 GND.t872 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X550 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30.t2 GND.t9 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X551 GND.t278 GND.t279 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t11 a_29780_7686.t3 GND.t636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X553 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t9 GND.t866 GND.t865 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X554 VDD.t199 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t3 VDD.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X555 GND.t176 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t1 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X556 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.t0 GND.t79 sky130_fd_pr__res_xhigh_po_1p41 l=3.94
X557 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t8 VDD.t222 VDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X558 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t31 VOUT.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 VDD.t140 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t2 VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X560 VDDH.t435 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t13 a_43724_16856.t1 VDDH.t434 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X561 a_6923_9707.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t25 GND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X562 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t12 a_20823_20174.t0 GND.t783 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X563 VDDH.t304 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t56 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t12 VDDH.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X564 GND.t751 GND.t752 GND.t81 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X565 a_43724_10362.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t14 VDDH.t437 VDDH.t436 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X566 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t9 GND.t818 GND.t817 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X567 GND.t940 DIN4.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t2 GND.t939 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X568 VDD.t134 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t3 VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X569 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t10 GND.t645 GND.t644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X570 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t40 GND.t952 GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X571 a_14948_18696.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13.t2 VDDH.t399 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X572 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t1 GND.t387 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X573 VDD.t174 DIN0.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t0 VDD.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X574 GND.t716 DIN7.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t0 GND.t715 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X575 VDD.t96 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t2 VDD.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X576 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X577 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t8 VDDH.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X578 a_16891_7686.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t2 VDDH.t424 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X579 a_5050_12595.t8 VOUT.t64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t22 GND.t872 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X580 GND.t694 GND.t695 GND.t693 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X581 a_15593_6250.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t0 VDDH.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X582 VDD.t116 DIN3.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t0 VDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X583 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t32 VOUT.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t3 VDDH.t68 VDDH.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X585 a_17443_7686.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t2 VDDH.t531 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X586 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t57 VDDH.t305 VDDH.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X587 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t10 VDDH.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X588 a_43167_3162.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t8 GND.t143 GND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X589 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t21 a_8051_10107.t8 GND.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X590 a_14672_18696.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t5 a_14514_18696.t0 VDDH.t496 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X591 VDDH.t306 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t58 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t12 VDDH.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X592 GND.t709 GND.t710 GND.t19 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X593 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t15 VDDH.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X594 GND.t738 GND.t739 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X595 VDDH.t274 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t0 VDDH.t273 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X596 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t9 VDD.t22 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X597 a_35453_10031.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t4 a_34873_10031.t2 GND.t666 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X598 VDDH.t189 VDDH.t187 VDDH.t188 VDDH.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X599 GND.t953 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t23 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X600 a_42724_19156.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t7 VDDH.t369 VDDH.t368 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X601 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t42 GND.t467 GND.t429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X602 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t12 VDDH.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X603 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t6 VDDH.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X604 a_15869_6250.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t2 VDDH.t532 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X605 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t16 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X606 a_44479_4254.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t3 a_44479_4170.t1 GND.t410 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X607 GND.t946 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 a_44062_18805.t1 GND.t945 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X608 VOUT.t39 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t7 VDDH.t548 VDDH.t547 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X609 GND.t82 GND.t83 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X610 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t0 GND.t41 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X611 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t60 VDDH.t276 VDDH.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X612 top_DAC_0/top_final_switch_0.VOUT[4].t3 top_DAC_0/top_rseg_n_dcell_0.SH[3].t3 a_15863_13785.t2 VDDH.t563 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X613 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t29 VDDH.t273 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X614 GND.t903 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 a_44062_20229.t1 GND.t902 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X615 a_16596_18696.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.t1 VDDH.t400 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X616 a_43167_4634.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t10 GND.t174 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X617 a_15618_18696.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t4 a_14672_18696.t3 VDDH.t442 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X618 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t61 VDDH.t278 VDDH.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X619 a_44234_11312.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t4 GND.t774 GND.t773 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X620 a_29158_6250.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6.t2 GND.t749 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X621 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t10 VOUT.t65 a_8051_10107.t14 GND.t661 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X622 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t10 VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X623 a_23049_18133.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t13 top_DAC_0/top_rseg_n_dcell_0.VH2.t3 GND.t613 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X624 VDDH.t280 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t10 VDDH.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X625 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t25 VDDH.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X626 VDD.t64 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t3 VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X627 a_21651_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t3 a_22469_18133.t2 GND.t900 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X628 a_8506_12595.t8 VOUT.t66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t4 GND.t802 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X629 GND.t304 GND.t305 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 a_43724_7392.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t15 VDDH.t439 VDDH.t438 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X631 VDD.t98 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X632 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t14 a_29780_7686.t0 GND.t600 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X633 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t27 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X634 GND.t974 GND.t975 GND.t88 sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X635 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t7 VDD.t136 VDD.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X636 top_DAC_0/top_rseg_n_dcell_0.VL2.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t11 a_14615_14283.t2 GND.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X637 VDD.t99 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t3 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X638 a_43167_3438.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t9 GND.t560 GND.t559 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X639 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t9 top_DAC_0/top_final_switch_0.VOUT[3].t6 a_8051_10107.t2 GND.t661 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X640 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t1 DIN0.t1 VDD.t176 VDD.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X641 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t11 VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X642 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t10 a_27896_6250.t1 GND.t627 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X643 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t43 GND.t469 GND.t468 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X644 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35.t2 GND.t22 sky130_fd_pr__res_xhigh_po_1p41 l=4.81
X645 a_8506_12595.t7 top_DAC_0/top_final_switch_0.VOUT[2].t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t15 GND.t802 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X646 GND.t535 GND.t536 GND.t13 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X647 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t1 DIN3.t1 VDD.t118 VDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X648 GND.t688 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t1 GND.t687 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 a_43724_6956.t0 a_43698_6796.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t1 VDDH.t526 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X650 a_15041_6250.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t4 a_19670_8950.t1 VDDH.t343 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X651 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t15 a_30608_7686.t0 GND.t601 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X652 GND.t470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t20 GND.t432 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X653 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t23 a_6923_9707.t6 GND.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X654 GND.t302 GND.t303 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 GND.t100 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t6 GND.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X656 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t35 VOUT.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t9 a_27896_6250.t2 GND.t750 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X658 a_8473_23194.t3 ROUT1.t4 a_4415_23194.t1 VDDH.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X659 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t3 DIN6.t1 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X660 GND.t300 GND.t301 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 a_15317_6250.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t2 VDDH.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X662 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t2 DIN2.t2 GND.t857 GND.t856 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X663 a_43724_13332.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t16 VDDH.t3 VDDH.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X664 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t45 GND.t472 GND.t471 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X665 GND.t299 GND.t297 GND.t298 GND.t217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X666 a_44479_3254.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t9 GND.t830 GND.t829 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X667 a_29158_6250.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t16 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22.t0 GND.t602 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X668 GND.t726 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t4 a_44234_6996.t1 GND.t725 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X669 VDDH.t186 VDDH.t184 VDDH.t185 VDDH.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X670 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13.t0 GND.t79 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X671 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t13 a_22755_20174.t0 GND.t784 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X672 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t6 a_16181_7686.t2 VDDH.t487 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X673 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t12 a_27896_6250.t4 GND.t637 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X674 a_28882_6250.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5.t1 GND.t871 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X675 GND.t168 GND.t169 GND.t41 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X676 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42.t0 GND.t13 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X677 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t11 GND.t539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.087 pd=0.89 as=0.174 ps=1.78 w=0.6 l=20
X678 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t3 GND.t4 GND.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X679 a_42982_19554.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t5 a_42724_19554.t0 VDDH.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X680 VDD.t207 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t1 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X681 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t9 VDDH.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X682 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t12 a_43391_3878.t1 GND.t578 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X683 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t24 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t6 GND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X684 GND.t474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t6 GND.t473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X685 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t36 VOUT.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 a_17167_7686.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t2 VDDH.t486 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X687 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t30 VDDH.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X688 a_43391_3794.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t10 a_43391_3710.t1 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X689 GND.t881 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t7 a_44234_15906.t1 GND.t504 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X690 GND.t296 GND.t294 GND.t295 GND.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X691 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t7 GND.t419 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X692 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t1 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=1.94
X693 a_42982_20978.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t9 a_42724_20978.t1 VDDH.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X694 a_34580_8950.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t5 a_31318_7686.t3 GND.t458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X695 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t3 a_4415_23194.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t21 VDDH.t456 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X696 a_8051_10107.t1 top_DAC_0/top_final_switch_0.VOUT[3].t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t10 GND.t662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X697 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t14 a_24963_20174.t0 GND.t785 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X698 a_16615_7686.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t1 VDDH.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X699 VDDH.t281 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t10 VDDH.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X700 a_35132_8950.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t6 a_31870_7686.t1 GND.t459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X701 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t26 a_8051_10107.t7 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X702 a_43698_14716.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t16 a_44234_15272.t1 GND.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X703 VOUT.t44 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t6 GND.t876 GND.t875 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X704 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t10 VDD.t150 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X705 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t26 top_DAC_0/top_final_switch_0.VOUT[4].t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t18 VDDH.t543 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X706 a_15863_13536.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t4 top_DAC_0/top_rseg_n_dcell_0.VH3.t2 VDDH.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X707 a_44062_18449.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 GND.t86 GND.t85 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X708 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t6 GND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X709 a_20352_10031.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t6 a_20222_8950.t0 VDDH.t307 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X710 a_16320_18696.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3.t1 VDDH.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X711 top_DAC_0/top_rseg_n_dcell_0.VS4.t5 top_DAC_0/top_rseg_n_dcell_0.SH[4].t4 top_DAC_0/top_final_switch_0.VOUT[1].t2 VDDH.t419 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X712 VDDH.t183 VDDH.t181 VDDH.t182 VDDH.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X713 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t4 a_45023_19116.t0 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X714 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t26 VOUT.t67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t22 VDDH.t543 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X715 GND.t293 GND.t291 GND.t292 GND.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X716 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X717 a_8051_10107.t13 VOUT.t68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t9 GND.t662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X718 a_17443_7686.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t2 VDDH.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X719 a_31594_7686.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62.t0 GND.t628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X720 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t8 a_15905_7686.t2 VDDH.t485 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X721 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t7 GND.t690 GND.t689 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X722 GND.t7 GND.t8 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=5.22
X723 VDD.t204 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t4 a_42847_4906.t1 VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X724 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t15 a_23583_20174.t1 GND.t786 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X725 a_19772_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t4 top_DAC_0/top_rseg_n_dcell_0.VS4.t0 VDDH.t312 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X726 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t33 VOUT.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 VDDH.t180 VDDH.t178 VDDH.t179 VDDH.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X728 a_44255_3714.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t10 GND.t868 GND.t867 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X729 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t8 GND.t883 GND.t882 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X730 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t11 a_45023_20540.t0 GND.t936 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X731 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t0 GND.t41 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X732 a_43698_9766.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t3 a_43724_10362.t0 VDDH.t575 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X733 a_15098_19866.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t0 VDDH.t71 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X734 VDD.t209 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t1 VDD.t208 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X735 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t0 DIN1.t2 GND.t484 GND.t483 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X736 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t6 VDD.t201 VDD.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X737 VDDH.t282 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t9 VDDH.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X738 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t6 VDDH.t524 VDDH.t523 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X739 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18.t2 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X740 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t1 VDDH.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X741 VDD.t152 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t4 VDD.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X742 a_16891_7686.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t2 VDDH.t484 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X743 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t0 GND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X744 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t0 GND.t19 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X745 a_43724_13886.t1 a_43698_13726.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t1 VDDH.t339 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X746 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t2 VDDH.t349 VDDH.t348 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X747 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t2 top_DAC_0/top_final_switch_0.VOUT[0].t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t16 VDDH.t558 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X748 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t7 VDDH.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X749 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t9 a_45023_18288.t1 GND.t884 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X750 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t2 a_43240_21320.t1 VDDH.t382 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X751 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t0 GND.t88 sky130_fd_pr__res_xhigh_po_1p41 l=1.63
X752 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t65 VDDH.t283 VDDH.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X753 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t8 VOUT.t69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t10 VDDH.t558 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X754 GND.t290 GND.t288 GND.t289 GND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X755 a_6923_9707.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t0 GND.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X756 a_42847_3710.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t1 VDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X757 a_42724_19554.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t8 VDDH.t370 VDDH.t365 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X758 a_35453_10031.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t7 a_33910_8950.t0 GND.t391 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X759 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t5 a_13779_6250.t4 VDDH.t533 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X760 GND.t276 GND.t277 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 a_20656_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t8 a_19000_8950.t0 VDDH.t247 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X762 VDDH.t177 VDDH.t175 VDDH.t176 VDDH.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X763 a_23859_20174.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t6 a_24209_18133.t0 GND.t737 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X764 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.t0 GND.t60 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X765 a_16615_7686.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t2 VDDH.t534 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X766 a_24963_20174.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t5 a_22469_18133.t4 GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X767 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32.t0 GND.t9 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X768 a_42724_20978.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t9 VDDH.t410 VDDH.t365 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X769 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14.t1 GND.t57 sky130_fd_pr__res_xhigh_po_1p41 l=1.84
X770 a_42982_18472.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t11 a_42724_18472.t1 VDDH.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X771 a_15317_6250.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t0 VDDH.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X772 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t32 VDDH.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X773 GND.t275 GND.t272 GND.t274 GND.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X774 a_44234_7986.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t0 GND.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X775 VDDH.t358 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t7 VDDH.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X776 a_44234_15272.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t5 GND.t16 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X777 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t7 a_14607_6250.t4 VDDH.t420 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X778 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t47 GND.t476 GND.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X779 GND.t477 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t19 GND.t436 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X780 a_45023_19116.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t5 GND.t503 GND.t502 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X781 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t6 GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X782 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t37 VOUT.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 a_14948_18696.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.t0 VDDH.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X784 a_44062_22009.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 GND.t532 GND.t531 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X785 VDDH.t527 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t13 VDDH.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X786 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t7 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X787 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t5 VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X788 a_15593_6250.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t0 VDDH.t421 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X789 a_43698_6796.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t3 a_43724_7392.t1 VDDH.t334 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X790 GND.t478 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t18 GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X791 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t0 VDDH.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X792 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t6 a_45023_18564.t0 GND.t17 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X793 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.t1 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X794 GND.t270 GND.t271 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X795 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.t1 GND.t38 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X796 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t10 VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X797 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t17 VOUT.t70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t14 VDDH.t453 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X798 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X799 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t1 VDDH.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X800 a_17443_7686.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t6 VDDH.t64 VDDH.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X801 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t2 top_DAC_0/top_final_switch_0.VOUT[3].t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t2 VDDH.t453 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X802 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t8 VOUT.t71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t12 VDDH.t320 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X803 a_45023_18288.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t8 GND.t728 GND.t727 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X804 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.t0 GND.t60 sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X805 a_43724_17292.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t17 VDDH.t5 VDDH.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X806 GND.t646 GND.t647 GND.t22 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X807 a_23307_20174.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t6 a_24209_18133.t4 GND.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X808 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t4 top_DAC_0/top_final_switch_0.VOUT[2].t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t7 VDDH.t320 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X809 a_22203_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t4 a_22469_18133.t1 GND.t683 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X810 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t5 VDD.t130 VDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X811 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t31 a_6923_9707.t1 GND.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X812 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t34 VOUT.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X813 a_43698_12736.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t4 a_43724_13332.t0 VDDH.t451 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X814 GND.t430 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t10 GND.t429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X815 VDD.t183 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t2 VDD.t182 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X816 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t10 a_22479_20174.t3 GND.t401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X817 a_43724_16856.t0 a_43698_16696.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t1 VDDH.t503 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X818 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t11 a_44255_3162.t1 GND.t172 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X819 top_DAC_0/top_rseg_n_dcell_0.VL3.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t12 a_18008_18696.t2 VDDH.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X820 a_43698_6796.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t18 a_44234_7352.t1 GND.t904 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X821 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4.t2 GND.t368 sky130_fd_pr__res_xhigh_po_1p41 l=3.12
X822 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t13 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t5 VDDH.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X823 GND.t972 GND.t973 GND.t18 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X824 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t2 DIN9.t2 VDD.t72 VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X825 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52.t2 GND.t361 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X826 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t8 GND.t374 GND.t373 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X827 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t17 a_27896_6250.t0 GND.t603 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X828 a_42724_18472.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t10 VDDH.t411 VDDH.t368 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X829 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t67 VDDH.t359 VDDH.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X830 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.t0 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X831 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t12 a_27620_6250.t2 GND.t748 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X832 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t68 VDDH.t360 VDDH.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X833 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44.t0 GND.t13 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X834 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t12 a_27620_6250.t1 GND.t629 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X835 a_37410_19098.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t3 GND.t367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X836 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t0 GND.t19 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X837 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t11 VDD.t158 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X838 a_43240_19156.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t18 a_42982_19156.t0 VDDH.t417 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X839 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t11 a_21099_20174.t3 GND.t402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X840 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t6 a_43391_4174.t1 GND.t490 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X841 a_8506_12595.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t3 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X842 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t11 a_22479_20174.t2 GND.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X843 a_6923_9707.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t4 GND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X844 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t14 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t0 VDDH.t345 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X845 VDDH.t361 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t6 VDDH.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X846 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t2 GND.t384 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.087 ps=0.89 w=0.6 l=20
X847 VDD.t58 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X848 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X849 a_15317_6250.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t7 a_19946_8950.t0 VDDH.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X850 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.t0 GND.t57 sky130_fd_pr__res_xhigh_po_1p41 l=2.09
X851 a_28606_6250.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t13 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52.t0 GND.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X852 GND.t676 GND.t677 GND.t13 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X853 GND.t431 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t2 GND.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X854 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t0 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X855 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t13 VDDH.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X856 a_6923_9707.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t5 GND.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X857 a_22755_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t5 a_24209_18133.t1 GND.t630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X858 a_14790_18696.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t5 a_16872_18696.t2 VDDH.t443 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X859 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t6 a_15353_7686.t0 VDDH.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X860 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t13 a_27620_6250.t4 GND.t680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X861 VDDH.t174 VDDH.t172 VDDH.t173 VDDH.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X862 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t1 top_DAC_0/top_final_switch_0.VOUT[3].t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t1 VDDH.t454 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X863 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t9 VDDH.t580 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X864 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t70 VDDH.t362 VDDH.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X865 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t52 GND.t433 GND.t432 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X866 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t12 a_21099_20174.t2 GND.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X867 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t34 VDDH.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X868 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t71 VDDH.t363 VDDH.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X869 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t13 VOUT.t72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t16 VDDH.t454 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X870 a_39306_20477.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t3 GND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X871 a_15629_7686.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t13 a_19000_8950.t2 VDDH.t241 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X872 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t19 a_27620_6250.t0 GND.t604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X873 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t38 VOUT.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X874 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t7 a_16181_7686.t0 VDDH.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X875 a_36888_19786.t5 a_36888_19786.t4 GND.t699 GND.t698 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X876 top_DAC_0/top_rseg_n_dcell_0.SH[2].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t2 VDDH.t505 VDDH.t504 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X877 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t12 VDD.t185 VDD.t184 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X878 VDDH.t7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t18 a_43724_13886.t0 VDDH.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X879 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t39 VOUT.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X880 a_45023_20540.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t11 GND.t558 GND.t557 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X881 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.t1 GND.t81 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X882 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t6 GND.t756 GND.t755 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X883 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48.t2 GND.t361 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X884 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t1 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=2.04
X885 a_34873_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t7 top_DAC_0/top_rseg_n_dcell_0.VS1.t1 GND.t757 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X886 a_19670_8950.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t14 a_16615_7686.t1 VDDH.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X887 VDDH.t364 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t4 VDDH.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X888 a_15869_6250.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t2 VDDH.t483 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X889 a_39936_22083.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t5 VDDH.t467 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=1
X890 VDDH.t171 VDDH.t169 VDDH.t170 VDDH.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X891 a_17167_7686.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t1 VDDH.t340 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X892 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t0 GND.t54 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X893 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t11 a_15629_7686.t2 VDDH.t482 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X894 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t4 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X895 VDDH.t402 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t0 VDDH.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X896 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t15 VDDH.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X897 GND.t269 GND.t266 GND.t268 GND.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X898 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t3 GND.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X899 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30.t0 GND.t9 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X900 a_15593_6250.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t2 VDDH.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X901 top_DAC_0/top_rseg_n_dcell_0.VL3.t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t5 a_15863_13287.t1 VDDH.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X902 a_20498_8950.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t15 a_17443_7686.t1 VDDH.t243 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X903 GND.t257 GND.t258 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X904 GND.t944 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t2 a_44234_9966.t1 GND.t943 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X905 top_DAC_0/top_final_switch_0.VOUT[2].t2 top_DAC_0/top_rseg_n_dcell_0.SH[3].t4 a_15863_13287.t0 VDDH.t562 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X906 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t4 GND.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X907 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29.t1 GND.t60 sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X908 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.t0 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X909 VDDH.t168 VDDH.t166 VDDH.t167 VDDH.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X910 a_22469_18133.t5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t14 top_DAC_0/top_rseg_n_dcell_0.VH2.t6 GND.t681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X911 VDDH.t549 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t8 VOUT.t40 VDDH.t545 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X912 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52.t1 GND.t361 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X913 a_14615_14283.t0 top_DAC_0/top_rseg_n_dcell_0.SH[2].t4 top_DAC_0/top_final_switch_0.VOUT[4].t1 GND.t498 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X914 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t14 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t4 GND.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X915 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16.t2 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X916 GND.t255 GND.t256 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X917 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t53 GND.t434 GND.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X918 top_DAC_0/top_rseg_n_dcell_0.VL3.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t8 a_17732_18696.t1 VDDH.t375 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X919 VDDH.t165 VDDH.t162 VDDH.t164 VDDH.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X920 GND.t713 GND.t714 GND.t368 sky130_fd_pr__res_xhigh_po_1p41 l=2.5
X921 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t3 VDD.t180 VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X922 top_DAC_0/top_rseg_n_dcell_0.VL2.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t5 a_14615_13785.t1 GND.t487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X923 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.t0 GND.t22 sky130_fd_pr__res_xhigh_po_1p41 l=5.01
X924 top_DAC_0/top_final_switch_0.VOUT[0].t0 top_DAC_0/top_rseg_n_dcell_0.SH[1].t4 top_DAC_0/top_rseg_n_dcell_0.VS1.t4 GND.t455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X925 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t5 GND.t416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X926 a_20547_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t6 a_23049_18133.t2 GND.t631 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X927 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16.t0 GND.t57 sky130_fd_pr__res_xhigh_po_1p41 l=1.68
X928 a_34856_8950.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t9 a_31594_7686.t2 GND.t513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X929 VDDH.t452 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t0 VDDH.t380 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X930 GND.t388 GND.t389 GND.t387 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X931 VDDH.t9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t19 a_43724_7946.t1 VDDH.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X932 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t1 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X933 a_31042_7686.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60.t1 GND.t915 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X934 a_17148_18696.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.t1 VDDH.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X935 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t1 GND.t41 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X936 a_44062_21653.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t0 GND.t911 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X937 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42.t1 GND.t13 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X938 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t35 VOUT.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X939 VDDH.t551 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t5 VDDH.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X940 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.t2 GND.t22 sky130_fd_pr__res_xhigh_po_1p41 l=4.91
X941 a_45343_3978.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t3 a_45343_3894.t1 GND.t466 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X942 VDDH.t161 VDDH.t159 VDDH.t160 VDDH.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X943 a_31870_7686.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63.t1 GND.t916 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X944 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t24 VDDH.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X945 a_43698_16696.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t4 a_43724_17292.t0 VDDH.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X946 GND.t265 GND.t263 GND.t264 GND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X947 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t1 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X948 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17.t1 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X949 a_4415_23194.t0 ROUT1.t5 a_8473_23194.t0 VDDH.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X950 a_42982_21662.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t13 a_42724_21662.t1 VDDH.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X951 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t74 VDDH.t552 VDDH.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X952 GND.t500 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 a_44062_19517.t1 GND.t499 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X953 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6.t0 GND.t368 sky130_fd_pr__res_xhigh_po_1p41 l=2.66
X954 a_15317_6250.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t2 VDDH.t422 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X955 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t38 a_8506_12595.t4 GND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X956 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15.t2 GND.t79 sky130_fd_pr__res_xhigh_po_1p41 l=5.42
X957 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.t1 GND.t79 sky130_fd_pr__res_xhigh_po_1p41 l=4.19
X958 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.t0 GND.t80 sky130_fd_pr__res_xhigh_po_1p41 l=5.58
X959 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t40 VOUT.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X960 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t2 GND.t18 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X961 VDDH.t553 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t75 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t0 VDDH.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X962 a_15869_6250.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t2 VDDH.t341 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X963 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X964 GND.t435 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t14 GND.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X965 VDDH.t158 VDDH.t156 VDDH.t157 VDDH.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X966 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t13 a_43167_3438.t0 GND.t405 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X967 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t55 GND.t437 GND.t436 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X968 a_21099_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t4 a_23049_18133.t3 GND.t619 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X969 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t41 VOUT.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X970 a_43240_19554.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t7 a_42982_19554.t1 VDDH.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X971 VDDH.t155 VDDH.t153 VDDH.t154 VDDH.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X972 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t12 a_23859_20174.t3 GND.t403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X973 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t1 VDDH.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X974 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t0 GND.t387 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X975 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t3 VDD.t78 VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X976 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t3 GND.t461 GND.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X977 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t10 a_14607_6250.t0 VDDH.t518 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X978 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t8 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X979 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15.t0 GND.t38 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X980 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t47 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t28 VDDH.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X981 VDDH.t554 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t0 VDDH.t273 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X982 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t4 GND.t800 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X983 a_17167_7686.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t2 VDDH.t460 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X984 VDDH.t152 VDDH.t150 VDDH.t151 VDDH.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X985 a_8506_12595.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t1 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X986 GND.t692 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t8 a_44234_12936.t1 GND.t691 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X987 GND.t253 GND.t254 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X988 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t77 VDDH.t555 VDDH.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X989 VDDH.t149 VDDH.t147 VDDH.t148 VDDH.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X990 a_43240_20978.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t16 a_42982_20978.t0 VDDH.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X991 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t0 GND.t54 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X992 a_44234_13926.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t0 GND.t905 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X993 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t14 VDDH.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X994 a_20932_10031.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t8 a_19670_8950.t0 VDDH.t308 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X995 VDDH.t34 a_5111_8388.t2 a_5111_8388.t3 VDDH.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=0.696 ps=5.09 w=4.8 l=1
X996 GND.t878 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t7 VOUT.t45 GND.t877 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X997 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t9 VDD.t178 VDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X998 a_43698_11746.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t20 a_44234_12302.t1 GND.t906 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X999 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t14 a_23859_20174.t2 GND.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1000 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X1001 a_29158_6250.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t16 a_34856_8950.t2 GND.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1002 a_22193_18133.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t16 top_DAC_0/top_rseg_n_dcell_0.VH2.t7 GND.t917 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1003 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t17 a_27344_6250.t1 GND.t918 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1004 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t17 a_23031_20174.t0 GND.t777 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1005 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.t1 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=5.22
X1006 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t56 GND.t439 GND.t438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1007 VDDH.t146 VDDH.t144 VDDH.t145 VDDH.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1008 GND.t262 GND.t259 GND.t261 GND.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1009 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t2 a_36888_19786.t1 GND.t516 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1010 GND.t252 GND.t250 GND.t251 GND.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0 ps=0 w=1.6 l=1
X1011 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54.t2 GND.t361 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1012 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t5 GND.t593 GND.t592 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1013 GND.t746 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t14 a_27344_6250.t2 GND.t745 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1014 a_42724_21662.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t11 VDDH.t412 VDDH.t365 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1015 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62.t1 GND.t81 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1016 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t13 a_24687_20174.t3 GND.t404 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1017 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t15 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t5 GND.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X1018 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t0 VDDH.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1019 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t9 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1020 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t9 VDDH.t310 VDDH.t309 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1021 VDD.t40 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t3 VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1022 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t10 VDDH.t581 VDDH.t251 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1023 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t36 VOUT.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1024 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t15 a_28172_6250.t2 GND.t747 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1025 a_43724_10916.t0 a_43698_10756.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t1 VDDH.t521 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1026 GND.t444 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t13 GND.t416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1027 a_20932_10031.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t5 a_19772_10031.t2 VDDH.t458 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1028 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t40 a_6778_12595.t9 GND.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1029 a_42982_20580.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t5 a_42724_20580.t1 VDDH.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1030 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t2 VDDH.t80 VDDH.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1031 a_6923_9707.t13 top_DAC_0/top_final_switch_0.VOUT[4].t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t18 GND.t815 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1032 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t5 GND.t961 GND.t960 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1033 VDD.t154 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t2 VDD.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1034 GND.t246 GND.t247 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1035 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.t1 GND.t22 sky130_fd_pr__res_xhigh_po_1p41 l=5.01
X1036 a_15353_7686.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t17 a_18724_8950.t0 VDDH.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1037 a_20076_10031.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t10 a_20498_8950.t0 VDDH.t311 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1038 a_5111_8388.t5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t10 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t11 VDDH.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.696 pd=5.09 as=1.392 ps=10.18 w=4.8 l=1
X1039 a_36888_19786.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t1 GND.t515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1040 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t20 a_27344_6250.t0 GND.t605 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1041 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t14 a_44479_3530.t1 GND.t406 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1042 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t39 GND.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1043 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t9 a_45023_21688.t1 GND.t375 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1044 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t6 GND.t722 GND.t721 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1045 a_6923_9707.t21 VOUT.t73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t17 GND.t815 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1046 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t0 GND.t88 sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X1047 a_31318_7686.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t16 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13.t1 GND.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1048 a_16181_7686.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t18 a_19552_8950.t2 VDDH.t259 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1049 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t12 a_44479_3898.t1 GND.t556 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1050 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t58 GND.t445 GND.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1051 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.t1 GND.t167 sky130_fd_pr__res_xhigh_po_1p41 l=7.01
X1052 a_19000_8950.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t10 a_14055_6250.t2 VDDH.t376 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1053 GND.t447 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t17 GND.t446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1054 VDDH.t143 VDDH.t140 VDDH.t142 VDDH.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1055 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t21 a_28172_6250.t0 GND.t598 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1056 a_16891_7686.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t0 VDDH.t519 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1057 a_43240_18472.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t15 a_42982_18472.t1 VDDH.t417 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1058 a_14672_18696.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.t0 VDDH.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1059 a_45023_21412.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t4 GND.t565 GND.t564 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1060 VDDH.t556 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t4 VDDH.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1061 GND.t249 GND.t248 GND.t249 GND.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0 ps=0 w=1.6 l=1
X1062 VDD.t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t3 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1063 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t1 GND.t18 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1064 a_44234_12302.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t4 GND.t2 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1065 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t12 a_45343_3254.t0 GND.t831 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1066 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t29 VDDH.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1067 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t7 VDDH.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1068 GND.t244 GND.t245 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1069 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t31 VDDH.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1070 VDD.t62 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t0 VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1071 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t12 a_15353_7686.t2 VDDH.t481 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1072 a_43724_8382.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t20 VDDH.t11 VDDH.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1073 a_15593_6250.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t11 a_20222_8950.t1 VDDH.t377 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1074 GND.t243 GND.t241 GND.t242 GND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1075 top_DAC_0/top_final_switch_0.VOUT[3].t1 top_DAC_0/top_rseg_n_dcell_0.SH[1].t5 top_DAC_0/top_rseg_n_dcell_0.VS1.t2 GND.t456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1076 a_44234_16896.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t0 GND.t797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1077 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t6 VDDH.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1078 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17.t0 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=5.06
X1079 GND.t240 GND.t238 GND.t239 GND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1080 a_30332_7686.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t12 a_33910_8950.t1 GND.t514 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1081 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t0 GND.t41 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X1082 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.t2 GND.t57 sky130_fd_pr__res_xhigh_po_1p41 l=1.89
X1083 a_44062_19161.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t0 GND.t399 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1084 a_20823_20174.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t6 a_24209_18133.t2 GND.t618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1085 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t12 a_15629_7686.t3 VDDH.t520 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1086 a_43724_7946.t0 a_43698_7786.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t1 VDDH.t514 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1087 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t79 VDDH.t557 VDDH.t273 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1088 VDDH.t139 VDDH.t136 VDDH.t138 VDDH.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1089 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t0 GND.t19 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X1090 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t13 VDD.t156 VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1091 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.t2 GND.t22 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X1092 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t1 GND.t387 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1093 GND.t658 GND.t659 GND.t365 sky130_fd_pr__res_xhigh_po_1p41 l=3.83
X1094 a_31042_7686.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t17 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.t1 GND.t811 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1095 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t55 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t18 VDDH.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1096 a_15905_7686.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t19 a_19276_8950.t2 VDDH.t260 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1097 a_42724_20580.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t12 VDDH.t413 VDDH.t365 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1098 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t56 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t3 VDDH.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1099 a_44062_20585.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t0 GND.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1100 a_6923_9707.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t31 GND.t416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1101 a_43724_14322.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t21 VDDH.t13 VDDH.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1102 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t43 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t3 GND.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1103 VDDH.t492 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t0 VDDH.t380 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1104 GND.t810 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t7 a_44234_7986.t1 GND.t809 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1105 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t4 GND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1106 a_8051_10107.t12 VOUT.t74 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t8 GND.t663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1107 a_31870_7686.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15.t2 GND.t812 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1108 a_45023_21688.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t5 GND.t595 GND.t594 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1109 VDD.t26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t1 VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X1110 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t12 GND.t171 GND.t170 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1111 GND.t76 DIN6.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t0 GND.t75 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1112 a_44479_3898.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t12 GND.t127 GND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1113 GND.t237 GND.t235 GND.t236 GND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1114 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t14 VDD.t157 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t13 VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1116 VDDH.t560 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t0 VDDH.t380 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1117 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t3 DIN4.t2 GND.t942 GND.t941 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1118 VDD.t213 DIN2.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t3 VDD.t212 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1119 VDDH.t135 VDDH.t133 VDDH.t134 VDDH.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1120 VOUT.t46 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t8 GND.t879 GND.t875 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1121 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t14 VDDH.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1122 GND.t448 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t16 GND.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1123 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t58 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t37 VDDH.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1124 GND.t234 GND.t231 GND.t233 GND.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0 ps=0 w=1.6 l=1
X1125 a_8051_10107.t0 top_DAC_0/top_final_switch_0.VOUT[3].t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t11 GND.t663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1126 GND.t793 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t15 a_44234_16896.t0 GND.t504 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1127 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t13 VDD.t160 VDD.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1128 VDDH.t383 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t80 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t8 VDDH.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1129 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t37 VOUT.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1130 a_44062_19161.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 GND.t426 GND.t425 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X1131 a_15224_18696.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14.t0 VDDH.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1132 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t1 DIN7.t2 GND.t718 GND.t717 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1133 VDD.t195 DIN5.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t1 VDD.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1134 a_35757_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t9 a_34580_8950.t0 GND.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1135 a_20352_10031.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t6 a_19772_10031.t1 VDDH.t350 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1136 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t30 VDDH.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1137 VDDH.t132 VDDH.t129 VDDH.t131 VDDH.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1138 a_38672_20477.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t12 GND.t397 GND.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1769 pd=1.8 as=0.1769 ps=1.8 w=0.61 l=9.7
X1139 a_6778_12595.t5 top_DAC_0/top_final_switch_0.VOUT[1].t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t4 GND.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1140 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13.t1 GND.t79 sky130_fd_pr__res_xhigh_po_1p41 l=4.6
X1141 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1.t2 GND.t365 sky130_fd_pr__res_xhigh_po_1p41 l=3.17
X1142 VDD.t74 DIN8.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t2 VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1143 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t11 VDDH.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1144 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t4 VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1145 a_43698_15706.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t22 a_44234_16262.t1 GND.t797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1146 a_43994_22522.t3 ROUT2.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t4 VDDH.t338 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X1147 VDD.t21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t0 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1148 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t9 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t8 a_5111_8388.t4 VDDH.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=0.696 ps=5.09 w=4.8 l=1
X1149 a_44062_20585.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 GND.t744 GND.t743 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X1150 a_15041_6250.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t2 VDDH.t423 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1151 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.t1 GND.t57 sky130_fd_pr__res_xhigh_po_1p41 l=2.19
X1152 GND.t682 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t1 GND.t608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1153 a_15342_18696.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t6 a_16320_18696.t2 VDDH.t444 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1154 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t61 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t7 VDDH.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1155 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t4 a_44479_4254.t1 GND.t839 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1156 a_6778_12595.t8 VOUT.t75 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t14 GND.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1157 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t2 GND.t54 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X1158 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t15 a_20547_20174.t2 GND.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1159 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t62 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t3 VDDH.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X1160 top_DAC_0/top_rseg_n_dcell_0.SH[1].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t4 GND.t845 GND.t844 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1161 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t1 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=2.4
X1162 a_44479_4170.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t4 GND.t765 GND.t764 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1163 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t61 GND.t449 GND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1164 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t81 VDDH.t384 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1165 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t15 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1166 a_16891_7686.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.t2 VDDH.t461 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1167 a_44255_4614.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t4 a_44255_4530.t0 GND.t858 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1168 a_43698_10756.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t3 a_43724_11352.t0 VDDH.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X1169 GND.t620 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t1 GND.t608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1170 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t11 a_15629_7686.t1 VDDH.t321 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1171 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t13 a_14331_6250.t0 VDDH.t253 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1172 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.t1 GND.t60 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X1173 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t10 GND.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1174 a_43724_14876.t1 a_43698_14716.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t1 VDDH.t561 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1175 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t18 a_24411_20174.t1 GND.t778 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1176 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t62 GND.t450 GND.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1177 GND.t230 GND.t228 GND.t230 GND.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0 ps=0 w=1.6 l=1
X1178 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t3 VDDH.t353 VDDH.t352 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1179 GND.t932 GND.t933 GND.t9 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X1180 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t13 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1181 a_43391_3326.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t14 a_43391_3242.t0 GND.t832 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1182 GND.t226 GND.t227 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1183 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t18 a_43240_19156.t1 VDDH.t425 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1184 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.t0 GND.t81 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X1185 VDDH.t15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t22 a_43724_10916.t1 VDDH.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1186 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t6 VDD.t170 VDD.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1187 VDD.t193 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t3 VDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1188 a_28882_6250.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t20 a_34580_8950.t2 GND.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1189 a_36033_10031.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t11 a_33358_8950.t0 GND.t392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1190 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t8 a_45023_21964.t0 GND.t798 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1191 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t16 VDD.t142 VDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1192 a_17167_7686.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t2 VDDH.t322 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1193 a_44234_7352.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t2 GND.t582 GND.t581 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1194 GND.t893 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t1 GND.t892 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1195 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t7 VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1196 VDD.t54 DIN1.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t2 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1197 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14.t0 GND.t57 sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X1198 a_5111_8388.t1 a_5111_8388.t0 VDDH.t32 VDDH.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.696 pd=5.09 as=1.392 ps=10.18 w=4.8 l=1
X1199 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t0 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=1.78
X1200 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28.t1 GND.t9 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X1201 a_23583_20174.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t7 a_23049_18133.t0 GND.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1202 a_15374_19866.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t7 a_15342_18696.t1 VDDH.t525 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1203 a_14615_13785.t0 top_DAC_0/top_rseg_n_dcell_0.SH[2].t5 top_DAC_0/top_final_switch_0.VOUT[2].t0 GND.t497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X1204 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t2 DIN5.t3 VDD.t197 VDD.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1205 GND.t851 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t1 GND.t850 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1206 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t42 VOUT.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1207 GND.t225 GND.t222 GND.t224 GND.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1208 GND.t847 DIN0.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t2 GND.t846 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1209 a_18008_18696.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t6 a_15342_18696.t0 VDDH.t409 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1210 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t3 DIN8.t3 VDD.t76 VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1211 GND.t24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t0 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1212 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29.t0 GND.t60 sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X1213 a_8051_10107.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t2 GND.t419 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1214 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13.t1 GND.t38 sky130_fd_pr__res_xhigh_po_1p41 l=5.47
X1215 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t17 top_DAC_0/top_final_switch_0.VOUT[4].t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t25 VDDH.t544 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1216 a_44479_3530.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t15 GND.t121 GND.t120 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1217 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t4 VDDH.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1218 a_44234_8976.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t1 GND.t907 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1219 GND.t673 DIN3.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t2 GND.t672 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1220 a_44234_16262.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t7 GND.t505 GND.t504 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1221 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t47 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t0 GND.t501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X1222 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t82 VDDH.t385 VDDH.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1223 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54.t1 GND.t361 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1224 VDDH.t17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t23 a_39936_22083.t0 VDDH.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9.2
X1225 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t21 VOUT.t76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t25 VDDH.t544 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1226 a_5050_12595.t7 VOUT.t77 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t21 GND.t919 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1227 a_44062_18805.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t0 GND.t395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1228 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t48 a_8506_12595.t2 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1229 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3.t0 GND.t365 sky130_fd_pr__res_xhigh_po_1p41 l=3.37
X1230 VDD.t172 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t4 a_42847_3710.t1 VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1231 VDD.t94 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 VDD.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1232 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t83 VDDH.t386 VDDH.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1233 GND.t451 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t12 GND.t438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1234 a_31870_7686.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47.t2 GND.t684 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1235 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t4 GND.t542 GND.t541 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1236 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t64 GND.t453 GND.t452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1237 GND.t583 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t15 GND.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1238 a_43698_7786.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t3 a_43724_8382.t1 VDDH.t506 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X1239 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t0 GND.t18 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X1240 a_5050_12595.t1 top_DAC_0/top_final_switch_0.VOUT[0].t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t22 GND.t919 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1241 a_42982_18814.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t19 a_42724_18814.t1 VDDH.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1242 VDDH.t128 VDDH.t126 VDDH.t127 VDDH.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1243 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t1 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X1244 a_16596_18696.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2.t1 VDDH.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1245 VDDH.t387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t84 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t2 VDDH.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1246 a_35177_10031.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t12 a_34186_8950.t0 GND.t393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1247 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t85 VDDH.t388 VDDH.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1248 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.t2 GND.t361 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1249 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t43 VOUT.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1250 a_18724_8950.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t13 a_13779_6250.t1 VDDH.t414 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1251 a_43391_3710.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t16 GND.t123 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1252 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t15 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1253 GND.t220 GND.t221 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1254 GND.t585 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t13 GND.t584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1255 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t67 GND.t586 GND.t416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1256 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t10 a_14055_6250.t4 VDDH.t462 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1257 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t0 GND.t88 sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X1258 GND.t656 GND.t657 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X1259 a_15317_6250.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t2 VDDH.t480 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1260 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t0 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=2.14
X1261 a_19552_8950.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t14 a_14607_6250.t1 VDDH.t415 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1262 VDD.t128 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t3 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1263 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t2 GND.t19 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1264 VDDH.t125 VDDH.t123 VDDH.t124 VDDH.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1265 GND.t566 GND.t567 GND.t79 sky130_fd_pr__res_xhigh_po_1p41 l=5.42
X1266 GND.t841 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t0 GND.t840 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1267 a_43240_21662.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t14 a_42982_21662.t1 VDDH.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1268 a_43698_13726.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t4 a_43724_14322.t1 VDDH.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X1269 top_DAC_0/top_rseg_n_dcell_0.VS4.t6 top_DAC_0/top_rseg_n_dcell_0.SH[4].t5 top_DAC_0/top_final_switch_0.VOUT[4].t2 VDDH.t502 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X1270 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t86 VDDH.t389 VDDH.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1271 a_44062_18093.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t0 GND.t394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1272 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t3 VDDH.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1273 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t11 GND.t853 GND.t852 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1274 VDDH.t43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t87 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t1 VDDH.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1275 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t38 VOUT.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1276 a_15041_6250.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t2 VDDH.t463 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1277 GND.t219 GND.t216 GND.t218 GND.t217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1278 a_43994_22522.t1 ROUT2.t2 ROUT2.t3 VDDH.t338 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X1279 GND.t214 GND.t215 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1280 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t3 DIN0.t3 GND.t849 GND.t848 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1281 top_DAC_0/top_final_switch_0.VOUT[0].t3 top_DAC_0/top_rseg_n_dcell_0.SH[3].t5 top_DAC_0/top_rseg_n_dcell_0.VL3.t3 VDDH.t562 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1282 VDDH.t45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t88 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t2 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1283 a_43698_7786.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t24 a_44234_8342.t0 GND.t908 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1284 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t16 GND.t26 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1285 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t68 GND.t587 GND.t446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1286 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t3 DIN3.t3 GND.t675 GND.t674 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1287 VDD.t148 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 VDD.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1288 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t15 a_20547_20174.t3 GND.t703 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1289 a_15869_6250.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t2 VDDH.t464 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1290 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t20 a_30608_7686.t3 GND.t485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1291 a_30056_7686.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t15 a_33634_8950.t1 GND.t596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1292 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t1 DIN6.t3 GND.t78 GND.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1293 GND.t652 GND.t653 GND.t38 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X1294 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.t0 GND.t41 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X1295 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t7 GND.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1296 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t20 VOUT.t78 a_5050_12595.t6 GND.t920 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1297 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t12 VOUT.t79 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t15 VDDH.t455 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1298 a_20352_10031.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t10 a_19276_8950.t0 VDDH.t248 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1299 top_DAC_0/top_rseg_n_dcell_0.SH[4].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t4 GND.t580 GND.t579 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1300 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t4 GND.t697 GND.t696 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1301 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t0 top_DAC_0/top_final_switch_0.VOUT[3].t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t0 VDDH.t455 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1302 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t89 VDDH.t47 VDDH.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1303 a_31594_7686.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14.t2 GND.t486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1304 a_34304_8950.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t16 a_31042_7686.t1 GND.t597 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1305 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t20 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1306 a_15041_6250.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t1 VDDH.t479 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1307 a_16872_18696.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.t1 VDDH.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1308 ROUT1.t3 ROUT1.t2 a_8473_23194.t1 VDDH.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X1309 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t23 top_DAC_0/top_final_switch_0.VOUT[0].t9 a_5050_12595.t0 GND.t920 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1310 a_42724_18814.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t13 VDDH.t390 VDDH.t368 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1311 GND.t212 GND.t213 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1312 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.t2 GND.t167 sky130_fd_pr__res_xhigh_po_1p41 l=8.5
X1313 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t16 a_23307_20174.t2 GND.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1314 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t20 a_30332_7686.t1 GND.t621 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1315 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t8 GND.t419 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1316 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46.t0 GND.t13 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1317 a_44234_10956.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t25 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t0 GND.t909 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1318 a_18284_18696.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t3 a_15066_18696.t2 VDDH.t396 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1319 GND.t210 GND.t211 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1320 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t8 VDDH.t403 VDDH.t345 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X1321 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t1 top_DAC_0/top_final_switch_0.VOUT[1].t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t12 VDDH.t335 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1322 a_14615_14034.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t11 top_DAC_0/top_rseg_n_dcell_0.VH2.t0 GND.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1323 a_37410_19098.t3 a_37410_19098.t2 GND.t969 GND.t968 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1856 pd=1.86 as=0.1856 ps=1.86 w=0.64 l=12
X1324 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.t2 GND.t80 sky130_fd_pr__res_xhigh_po_1p41 l=5.32
X1325 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t6 VOUT.t80 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t20 VDDH.t335 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1326 a_44062_20229.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t0 GND.t400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1327 VDDH.t49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t90 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t2 VDDH.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1328 a_44255_4162.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t17 a_44255_4078.t1 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1329 a_31318_7686.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61.t0 GND.t622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1330 a_22755_20174.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t8 a_22193_18133.t0 GND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1331 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t9 GND.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1332 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t0 a_37410_19098.t0 GND.t799 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1333 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t17 a_21927_20174.t0 GND.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1334 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t52 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t0 GND.t501 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X1335 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.t0 GND.t38 sky130_fd_pr__res_xhigh_po_1p41 l=5.94
X1336 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62.t2 GND.t81 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1337 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t7 a_43240_19554.t0 VDDH.t382 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1338 VDDH.t122 VDDH.t120 VDDH.t121 VDDH.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1339 top_DAC_0/top_rseg_n_dcell_0.SH[3].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t4 VDDH.t517 VDDH.t516 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1340 VDDH.t19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t24 a_43724_14876.t0 VDDH.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1341 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t16 a_21375_20174.t3 GND.t704 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1342 a_44255_4530.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t4 a_44255_4446.t1 GND.t508 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1343 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t7 GND.t489 GND.t488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1344 a_42982_20238.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t7 a_42724_20238.t1 VDDH.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1345 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22.t2 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X1346 VDDH.t51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t91 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t5 VDDH.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1347 a_4415_23194.t5 a_4415_23194.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t1 VDDH.t457 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X1348 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1.t0 GND.t365 sky130_fd_pr__res_xhigh_po_1p41 l=3.27
X1349 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t1 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1350 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t3 a_43240_20978.t1 VDDH.t382 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1351 a_43391_3242.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t17 a_43391_3158.t1 GND.t794 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1352 top_DAC_0/top_rseg_n_dcell_0.VL3.t6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t6 a_15863_13536.t2 VDDH.t246 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X1353 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t20 VDDH.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1354 a_45023_18564.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t11 GND.t836 GND.t835 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1355 a_43240_20580.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t8 a_42982_20580.t0 VDDH.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1356 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t92 VDDH.t53 VDDH.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1357 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t16 VOUT.t81 a_6923_9707.t20 GND.t417 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1358 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t13 a_15353_7686.t4 VDDH.t323 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1359 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t15 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t1 VDDH.t345 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X1360 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t14 a_14055_6250.t0 VDDH.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1361 GND.t843 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t8 a_44234_10956.t1 GND.t842 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1362 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t8 GND.t895 GND.t894 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1363 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t39 VOUT.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1364 GND.t494 a_36888_19786.t2 a_36888_19786.t3 GND.t493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1365 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t40 VOUT.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1366 VDDH.t55 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t93 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t1 VDDH.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1367 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t19 top_DAC_0/top_final_switch_0.VOUT[4].t10 a_6923_9707.t14 GND.t417 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1368 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t0 GND.t19 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1369 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t14 a_16181_7686.t4 VDDH.t324 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1370 a_15041_6250.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t0 VDDH.t255 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1371 GND.t102 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t3 GND.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X1372 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t94 VDDH.t290 VDDH.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1373 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t0 GND.t18 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1374 top_DAC_0/top_final_switch_0.VOUT[1].t1 top_DAC_0/top_rseg_n_dcell_0.SH[1].t6 top_DAC_0/top_rseg_n_dcell_0.VS1.t3 GND.t455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1375 a_43994_22522.t2 ROUT2.t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t5 VDDH.t338 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X1376 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t15 a_14331_6250.t2 VDDH.t445 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1377 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t18 a_22755_20174.t3 GND.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1378 VDDH.t292 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t95 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t3 VDDH.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1379 a_18008_18696.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t4 a_14790_18696.t1 VDDH.t284 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1380 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t18 a_44255_4162.t0 GND.t795 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1381 VDDH.t119 VDDH.t117 VDDH.t118 VDDH.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1382 a_44255_3162.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t17 GND.t125 GND.t124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1383 a_6778_12595.t0 VOUT.t82 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t13 GND.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1384 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t16 a_45023_19988.t0 GND.t407 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1385 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t1 VDDH.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1386 a_44255_4078.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t15 GND.t874 GND.t873 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t7 VOUT.t83 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t9 VDDH.t325 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1388 VDDH.t116 VDDH.t113 VDDH.t115 VDDH.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1389 GND.t648 GND.t649 GND.t364 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X1390 VDDH.t112 VDDH.t110 VDDH.t111 VDDH.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1391 VDD.t189 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t1 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1392 VDDH.t582 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t2 VDDH.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1393 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t13 a_16181_7686.t3 VDDH.t465 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1394 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t1 top_DAC_0/top_final_switch_0.VOUT[0].t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t15 VDDH.t325 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1395 GND.t208 GND.t209 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1396 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t0 VDDH.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1397 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.t2 GND.t167 sky130_fd_pr__res_xhigh_po_1p41 l=11.57
X1398 a_44255_4446.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t5 GND.t651 GND.t650 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1399 a_6778_12595.t4 top_DAC_0/top_final_switch_0.VOUT[1].t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t3 GND.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1400 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t1 VDDH.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1401 VDDH.t293 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t96 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t1 VDDH.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1402 a_43391_4174.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t6 GND.t414 GND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1403 GND.t408 GND.t409 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X1404 a_42724_20238.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t14 VDDH.t391 VDDH.t365 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1405 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t12 VDDH.t583 VDDH.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1406 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t15 GND.t804 GND.t803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X1407 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t1 GND.t387 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1408 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.t1 GND.t167 sky130_fd_pr__res_xhigh_po_1p41 l=7.88
X1409 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.t1 GND.t365 sky130_fd_pr__res_xhigh_po_1p41 l=3.83
X1410 a_31594_7686.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46.t2 GND.t685 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1411 a_43391_3158.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t14 GND.t555 GND.t554 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1412 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t22 a_43240_18472.t0 VDDH.t425 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1413 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t69 GND.t588 GND.t419 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1414 VDD.t9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t1 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1415 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.t2 GND.t80 sky130_fd_pr__res_xhigh_po_1p41 l=5.47
X1416 a_43724_11352.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t25 VDDH.t21 VDDH.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1417 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t8 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t9 VDDH.t404 VDDH.t345 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X1418 GND.t207 GND.t205 GND.t206 GND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1419 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t21 VDDH.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1420 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19.t0 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X1421 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t6 VDDH.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1422 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t17 a_23307_20174.t4 GND.t705 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1423 a_6923_9707.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t2 GND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1424 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t44 VOUT.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1425 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t45 VOUT.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1426 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t14 a_13779_6250.t3 VDDH.t576 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1427 a_44255_3438.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t15 GND.t553 GND.t552 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1428 top_DAC_0/top_final_switch_0.VOUT[3].t2 top_DAC_0/top_rseg_n_dcell_0.SH[3].t6 a_15863_13536.t0 VDDH.t562 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1429 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t16 a_45023_20264.t0 GND.t551 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1430 a_44234_10322.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t5 GND.t544 GND.t543 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1431 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t70 GND.t589 GND.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1432 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t4 GND.t492 GND.t491 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1433 GND.t632 GND.t633 GND.t88 sky130_fd_pr__res_xhigh_po_1p41 l=1.63
X1434 a_19276_8950.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t17 a_14331_6250.t1 VDDH.t416 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1435 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t2 VDDH.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1436 GND.t880 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t9 VOUT.t47 GND.t877 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1437 a_24209_18133.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t22 top_DAC_0/top_rseg_n_dcell_0.VL2.t6 GND.t519 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1438 VDDH.t109 VDDH.t106 VDDH.t108 VDDH.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1439 a_23031_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t9 a_23049_18133.t4 GND.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1440 VDD.t191 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t2 VDD.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1441 VDDH.t584 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t3 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1442 GND.t590 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t10 GND.t452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1443 GND.t758 GND.t759 GND.t365 sky130_fd_pr__res_xhigh_po_1p41 l=3.17
X1444 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t55 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t1 GND.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1445 GND.t383 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t8 a_44234_13926.t0 GND.t382 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1446 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t15 a_14607_6250.t3 VDDH.t577 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1447 a_44234_14916.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t0 GND.t910 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1448 a_44062_19873.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t0 GND.t576 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1449 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t18 a_21927_20174.t2 GND.t706 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1450 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t0 a_4415_23194.t2 a_4415_23194.t3 VDDH.t456 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X1451 GND.t203 GND.t204 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1452 GND.t976 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t8 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1453 a_31318_7686.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45.t1 GND.t686 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1454 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t56 a_6923_9707.t3 GND.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1455 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t12 VDDH.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1456 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t23 a_29780_7686.t4 GND.t711 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1457 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t8 VOUT.t84 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t6 VDDH.t286 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1458 a_43698_12736.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t27 a_44234_13292.t1 GND.t796 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1459 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t5 VDDH.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1460 a_29780_7686.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t18 a_33358_8950.t1 GND.t525 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t73 GND.t977 GND.t584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t18 top_DAC_0/top_final_switch_0.VOUT[0].t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t0 VDDH.t286 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1463 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t15 a_13779_6250.t2 VDDH.t478 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1464 GND.t201 GND.t202 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1465 GND.t712 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t1 GND.t608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1466 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48.t0 GND.t13 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X1467 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t0 GND.t54 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X1468 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t19 a_24687_20174.t2 GND.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1469 GND.t199 GND.t200 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t97 VDDH.t294 VDDH.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1471 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t8 GND.t736 GND.t735 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1472 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t5 VDDH.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1473 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.t0 GND.t364 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X1474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t2 GND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1475 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t19 a_24135_20174.t3 GND.t707 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1476 VDD.t217 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t2 VDD.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X1477 VDD.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1478 a_30608_7686.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t19 a_34186_8950.t1 GND.t526 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1479 a_35757_10031.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t8 a_34569_10031.t1 GND.t422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1480 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t16 a_14607_6250.t2 VDDH.t477 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1481 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t74 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t5 VDDH.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1482 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t19 a_21099_20174.t0 GND.t779 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1483 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t16 a_15905_7686.t0 VDDH.t356 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1484 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.t1 GND.t365 sky130_fd_pr__res_xhigh_po_1p41 l=3.53
X1485 GND.t805 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t22 GND.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X1486 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t23 a_30056_7686.t2 GND.t623 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1487 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t58 a_8051_10107.t5 GND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1488 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t19 VDD.t144 VDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1489 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t21 VDDH.t355 VDDH.t354 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1490 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t75 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t2 VDDH.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1491 VDDH.t105 VDDH.t102 VDDH.t104 VDDH.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1492 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t4 VDDH.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1493 a_44062_19873.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 GND.t926 GND.t925 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X1494 a_43724_11906.t0 a_43698_11746.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t0 VDDH.t244 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1495 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t3 VDDH.t536 VDDH.t535 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1496 VDD.t46 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1497 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t16 a_14331_6250.t4 VDDH.t578 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1498 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t77 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t16 VDDH.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1499 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t1 GND.t18 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1500 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t41 VOUT.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1501 a_15593_6250.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t2 VDDH.t476 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1502 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t20 a_22755_20174.t4 GND.t708 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1503 GND.t369 GND.t370 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X1504 VDDH.t101 VDDH.t98 VDDH.t100 VDDH.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1505 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t59 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t0 GND.t416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1506 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t28 VDDH.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1507 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31.t1 GND.t60 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X1508 a_45343_3894.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t4 GND.t562 GND.t561 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1509 GND.t741 GND.t742 GND.t368 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X1510 VDD.t162 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 VDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1511 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t79 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t35 VDDH.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1512 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t4 VDDH.t251 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1513 a_42982_22004.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t20 a_42724_22004.t1 VDDH.t257 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1514 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.t2 GND.t57 sky130_fd_pr__res_xhigh_po_1p41 l=2.35
X1515 VDDH.t97 VDDH.t95 VDDH.t96 VDDH.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1516 VDD.t168 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t1 VDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1517 a_8051_10107.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t0 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1518 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t61 a_6923_9707.t17 GND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1519 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t23 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t17 GND.t806 GND.t803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X1520 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t24 VOUT.t85 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t20 VDDH.t326 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1521 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t62 a_6923_9707.t18 GND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1522 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t19 a_45023_19712.t1 GND.t376 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1523 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36.t1 GND.t364 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X1524 a_44234_13292.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t4 GND.t569 GND.t568 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1525 a_31318_7686.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t22 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29.t1 GND.t599 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1526 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t24 top_DAC_0/top_final_switch_0.VOUT[4].t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t16 VDDH.t326 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1527 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t2 GND.t19 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X1528 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t46 VOUT.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1529 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t74 GND.t978 GND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1530 VOUT.t41 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t9 VDDH.t550 VDDH.t547 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1531 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t80 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t1 VDDH.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1532 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t1 GND.t548 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1533 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t17 a_13779_6250.t0 VDDH.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1534 GND.t197 GND.t198 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1535 a_43724_9372.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t26 VDDH.t23 VDDH.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1536 GND.t196 GND.t193 GND.t195 GND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1537 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t81 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t0 VDDH.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1538 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t82 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t3 VDDH.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X1539 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.t0 GND.t167 sky130_fd_pr__res_xhigh_po_1p41 l=9.22
X1540 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t8 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1541 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t21 a_24135_20174.t2 GND.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1542 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t0 GND.t88 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X1543 a_43240_18814.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t23 a_42982_18814.t0 VDDH.t417 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1544 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t83 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t27 VDDH.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1545 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t16 a_15905_7686.t4 VDDH.t446 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1546 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t21 a_23583_20174.t3 GND.t702 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1547 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t24 a_30608_7686.t1 GND.t624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1548 a_15863_13785.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t13 top_DAC_0/top_rseg_n_dcell_0.VH3.t0 VDDH.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1549 a_44062_21297.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t0 GND.t564 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1550 a_42982_18130.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t24 a_42724_18130.t1 VDDH.t418 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1551 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t9 VOUT.t86 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t19 VDDH.t327 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1552 a_42982_19896.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t8 a_42724_19896.t1 VDDH.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1553 top_DAC_0/top_rseg_n_dcell_0.VS4.t2 top_DAC_0/top_rseg_n_dcell_0.SH[4].t6 top_DAC_0/top_final_switch_0.VOUT[2].t3 VDDH.t419 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X1554 a_43724_8936.t0 a_43698_8776.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t0 VDDH.t331 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1555 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t0 GND.t19 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X1556 GND.t104 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 a_44062_20941.t1 GND.t103 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X1557 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t17 a_14055_6250.t1 VDDH.t447 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1558 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.t2 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X1559 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t0 top_DAC_0/top_final_switch_0.VOUT[1].t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t11 VDDH.t327 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1560 a_29434_6250.t4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t22 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39.t2 GND.t859 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1561 GND.t192 GND.t189 GND.t191 GND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1562 VDD.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1563 a_20823_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t8 a_22193_18133.t3 GND.t533 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1564 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t84 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t12 VDDH.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1565 GND.t187 GND.t188 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1566 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t5 VDD.t131 VDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1567 a_43724_15312.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t27 VDDH.t25 VDDH.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1568 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t63 a_5050_12595.t4 GND.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1569 GND.t521 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t2 a_44234_8976.t1 GND.t520 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1570 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t2 GND.t18 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X1571 a_5050_12595.t5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t0 GND.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1572 VDD.t125 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t1 VDD.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1573 top_DAC_0/top_rseg_n_dcell_0.VL2.t5 top_DAC_0/top_rseg_n_dcell_0.SH[2].t6 top_DAC_0/top_final_switch_0.VOUT[0].t1 GND.t497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X1574 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t12 VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1575 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t17 a_15905_7686.t3 VDDH.t579 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1576 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t12 VDDH.t475 VDDH.t474 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1577 a_35177_10031.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t7 a_34569_10031.t2 GND.t667 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1578 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t0 VDDH.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1579 GND.t729 GND.t730 GND.t81 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1580 GND.t185 GND.t186 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1581 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t7 a_36888_19550.t1 GND.t516 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1582 a_42724_22004.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t15 VDDH.t393 VDDH.t392 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1583 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t5 a_45343_3978.t0 GND.t614 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1584 a_44062_22009.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t1 GND.t816 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1585 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t42 VOUT.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1586 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t85 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t19 VDDH.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1587 GND.t979 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t75 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t4 GND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1588 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t13 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1589 a_44062_21297.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 GND.t834 GND.t833 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X1590 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t2 VDDH.t57 VDDH.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1591 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35.t1 GND.t22 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X1592 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t43 VOUT.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1593 a_20076_10031.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t9 a_19468_10031.t1 VDDH.t330 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1594 VDD.t33 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t2 VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1595 GND.t980 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t12 GND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1596 a_43698_16696.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t28 a_44234_17252.t1 GND.t797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1597 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t20 a_21651_20174.t0 GND.t780 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1598 a_16320_18696.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.t0 VDDH.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1599 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t20 VDD.t146 VDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1600 VDD.t17 DIN4.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t0 VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1601 top_DAC_0/top_rseg_n_dcell_0.VH3.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t20 a_18008_18696.t1 VDDH.t379 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1602 a_5111_10963.t4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t8 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t9 GND.t462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.464 ps=3.78 w=1.6 l=1
X1603 a_33910_8950.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t22 a_27896_6250.t3 GND.t495 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1604 a_22479_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t9 a_23629_18133.t2 GND.t534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1605 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46.t1 GND.t13 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1606 VDD.t127 DIN7.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t2 VDD.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1607 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t4 a_43240_21662.t0 VDDH.t382 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1608 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t98 VDDH.t295 VDDH.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1609 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.t1 GND.t13 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X1610 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t86 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t26 VDDH.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1611 a_21375_20174.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t9 a_22193_18133.t2 GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1612 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36.t0 GND.t364 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X1613 GND.t655 DIN9.t3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t3 GND.t654 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1614 top_DAC_0/top_rseg_n_dcell_0.SH[2].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t4 GND.t679 GND.t678 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1615 GND.t184 GND.t181 GND.t183 GND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1616 a_42724_18130.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t16 VDDH.t394 VDDH.t368 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1617 GND.t179 GND.t180 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1618 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t23 a_30056_7686.t4 GND.t860 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1619 a_42724_19896.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t17 VDDH.t366 VDDH.t365 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1620 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.t1 GND.t12 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X1621 GND.t731 GND.t732 GND.t387 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1622 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t87 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t39 VDDH.t273 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1623 VDDH.t94 VDDH.t92 VDDH.t93 VDDH.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1624 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t47 VOUT.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1625 VDDH.t296 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t99 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t0 VDDH.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1626 a_43698_11746.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t4 a_43724_12342.t0 VDDH.t537 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X1627 a_15098_19866.t2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.t2 VDDH.t289 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1628 a_43994_22522.t0 ROUT2.t0 ROUT2.t1 VDDH.t338 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X1629 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60.t2 GND.t81 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1630 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t77 GND.t981 GND.t332 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1631 GND.t982 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t10 GND.t419 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1632 a_43724_15866.t0 a_43698_15706.t2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t0 VDDH.t373 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1633 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t4 VDDH.t372 VDDH.t371 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1634 VDDH.t91 VDDH.t88 VDDH.t90 VDDH.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1635 a_31042_7686.t3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44.t1 GND.t861 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1636 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t79 GND.t983 GND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1637 a_45343_3254.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t17 GND.t550 GND.t549 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1638 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t12 VOUT.t87 a_6778_12595.t1 GND.t418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1639 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t100 VDDH.t298 VDDH.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1640 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.t1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.t0 GND.t167 sky130_fd_pr__res_xhigh_po_1p41 l=7.42
X1641 VDDH.t239 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t101 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t0 VDDH.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1642 VDDH.t27 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t28 a_43724_11906.t1 VDDH.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1643 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t66 a_6923_9707.t7 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1644 a_43240_20238.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t9 a_42982_20238.t0 VDDH.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1645 GND.t42 GND.t43 GND.t41 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X1646 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t12 GND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1647 VDDH.t87 VDDH.t84 VDDH.t86 VDDH.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1648 a_44234_8342.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t2 GND.t754 GND.t753 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1649 GND.t133 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t80 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t9 GND.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1650 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t81 GND.t134 GND.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1651 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t21 a_22479_20174.t0 GND.t781 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1652 VDD.t132 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t1 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
R0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t10 231.017
R1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t8 230.155
R2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t7 230.155
R3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t4 229.369
R4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t6 229.369
R5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t13 229.369
R6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t5 229.369
R7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n0 203.923
R8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t14 158.716
R9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n2 157.927
R10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t16 157.856
R11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t12 157.856
R12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t11 157.07
R13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t9 157.07
R14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t15 157.07
R15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t17 157.07
R16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n6 152.475
R17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n12 152.475
R18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n18 152.238
R19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n3 152
R20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n15 152
R21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n9 152
R22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n23 101.49
R23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t2 26.5955
R24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t3 26.5955
R25 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 25.0963
R26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t0 24.9236
R27 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t1 24.9236
R28 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n20 23.8264
R29 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n21 21.9086
R30 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n16 19.8154
R31 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n10 18.9229
R32 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n7 17.1938
R33 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n13 16.9661
R34 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n19 15.7596
R35 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n5 14.4113
R36 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n22 13.0565
R37 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n4 12.5635
R38 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n1 10.7525
R39 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 7.11161
R40 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 6.6565
R41 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 5.68939
R42 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 5.45235
R43 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 5.45235
R44 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 5.04292
R45 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 4.3525
R46 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 2.5605
R47 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 2.47068
R48 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 2.13383
R49 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 2.10199
R50 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n24 1.93989
R51 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n17 1.38917
R52 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n8 1.30714
R53 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n14 0.920422
R54 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n11 0.900891
R55 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.229016
R56 VDD.n343 VDD.t203 674.802
R57 VDD.n173 VDD.n111 674.766
R58 VDD.n172 VDD.n112 674.766
R59 VDD.t63 VDD.n193 633.369
R60 VDD.t77 VDD.n381 553.428
R61 VDD.n85 VDD.t67 465.683
R62 VDD.n382 VDD 432.123
R63 VDD.n418 VDD.t129 420.43
R64 VDD.n194 VDD.t198 420.25
R65 VDD.t119 VDD.n217 420.25
R66 VDD.n218 VDD.t39 420.25
R67 VDD.t133 VDD.n241 420.25
R68 VDD.n242 VDD.t192 420.25
R69 VDD.t153 VDD.n265 420.25
R70 VDD.n266 VDD.t95 420.25
R71 VDD.t32 VDD.n289 420.25
R72 VDD.n290 VDD.t182 420.25
R73 VDD.n173 VDD.t45 414.33
R74 VDD.t0 VDD.n112 414.33
R75 VDD.t171 VDD 411.372
R76 VDD.n144 VDD 401.233
R77 VDD.t173 VDD 369.938
R78 VDD VDD.t53 369.938
R79 VDD.t212 VDD 369.938
R80 VDD VDD.t115 369.938
R81 VDD.t16 VDD 369.938
R82 VDD VDD.t194 369.938
R83 VDD.t10 VDD 369.938
R84 VDD VDD.t126 369.938
R85 VDD.t73 VDD 369.938
R86 VDD VDD.t18 369.938
R87 VDD VDD.t106 366.978
R88 VDD.t208 VDD 366.978
R89 VDD VDD.t34 361.06
R90 VDD VDD.t147 361.06
R91 VDD VDD.t93 361.06
R92 VDD VDD.t84 361.06
R93 VDD VDD.t205 361.06
R94 VDD VDD.t97 361.06
R95 VDD.t57 VDD 361.06
R96 VDD.t2 VDD 361.06
R97 VDD.t161 VDD 361.06
R98 VDD VDD.t8 361.06
R99 VDD.t190 VDD 361.06
R100 VDD.n323 VDD.t26 340.301
R101 VDD.n403 VDD.t211 340.301
R102 VDD.n306 VDD.t217 336.416
R103 VDD.n412 VDD.n313 327.377
R104 VDD.n333 VDD.n332 320.976
R105 VDD.n328 VDD.n326 320.976
R106 VDD.n430 VDD.n429 318.305
R107 VDD.n405 VDD.n317 318.305
R108 VDD.n41 VDD.n40 318.303
R109 VDD VDD.t77 313.707
R110 VDD.n33 VDD.n10 313.575
R111 VDD.n4 VDD.n3 278.858
R112 VDD.n5 VDD.n3 278.858
R113 VDD.n437 VDD.n3 278.858
R114 VDD.n435 VDD.n3 278.858
R115 VDD.n14 VDD.n13 278.858
R116 VDD.n13 VDD.n12 278.858
R117 VDD.n13 VDD.n2 278.858
R118 VDD.n85 VDD 270.827
R119 VDD.n110 VDD 270.827
R120 VDD.n174 VDD 270.827
R121 VDD.n171 VDD 270.827
R122 VDD.n163 VDD 270.827
R123 VDD.n11 VDD.n2 269.485
R124 VDD.n437 VDD.n436 269.485
R125 VDD.n12 VDD.n11 269.485
R126 VDD.n436 VDD.n5 269.485
R127 VDD.n14 VDD.n11 269.485
R128 VDD.n436 VDD.n4 269.485
R129 VDD.n436 VDD.n435 269.485
R130 VDD.n86 VDD.n85 267.296
R131 VDD.n110 VDD.n109 267.296
R132 VDD.n175 VDD.n174 267.296
R133 VDD.n171 VDD.n170 267.296
R134 VDD.n164 VDD.n163 267.296
R135 VDD.n297 VDD.t19 255.905
R136 VDD.n51 VDD.t183 255.905
R137 VDD.n282 VDD.t74 255.905
R138 VDD.n53 VDD.t33 255.905
R139 VDD.n273 VDD.t127 255.905
R140 VDD.n57 VDD.t96 255.905
R141 VDD.n258 VDD.t11 255.905
R142 VDD.n59 VDD.t154 255.905
R143 VDD.n249 VDD.t195 255.905
R144 VDD.n63 VDD.t193 255.905
R145 VDD.n234 VDD.t17 255.905
R146 VDD.n65 VDD.t134 255.905
R147 VDD.n225 VDD.t116 255.905
R148 VDD.n69 VDD.t40 255.905
R149 VDD.n210 VDD.t213 255.905
R150 VDD.n71 VDD.t120 255.905
R151 VDD.n201 VDD.t54 255.905
R152 VDD.n75 VDD.t199 255.905
R153 VDD.n187 VDD.t174 255.905
R154 VDD.n77 VDD.t64 255.905
R155 VDD.n39 VDD.t70 255.905
R156 VDD.n375 VDD.t78 255.905
R157 VDD.n308 VDD.t130 255.905
R158 VDD.n45 VDD.t36 255.904
R159 VDD.n308 VDD.t131 255.904
R160 VDD.n299 VDD.t72 252.95
R161 VDD.n296 VDD.t185 252.95
R162 VDD.n52 VDD.t76 252.95
R163 VDD.n283 VDD.t66 252.95
R164 VDD.n54 VDD.t224 252.95
R165 VDD.n272 VDD.t101 252.95
R166 VDD.n58 VDD.t13 252.95
R167 VDD.n259 VDD.t146 252.95
R168 VDD.n60 VDD.t197 252.95
R169 VDD.n248 VDD.t164 252.95
R170 VDD.n64 VDD.t215 252.95
R171 VDD.n235 VDD.t136 252.95
R172 VDD.n66 VDD.t118 252.95
R173 VDD.n224 VDD.t42 252.95
R174 VDD.n70 VDD.t138 252.95
R175 VDD.n211 VDD.t122 252.95
R176 VDD.n72 VDD.t52 252.95
R177 VDD.n200 VDD.t201 252.95
R178 VDD.n76 VDD.t176 252.95
R179 VDD.n188 VDD.t170 252.95
R180 VDD.n315 VDD.t56 250.722
R181 VDD.n37 VDD.t202 249.901
R182 VDD.n31 VDD.t92 249.52
R183 VDD.n403 VDD.t160 249.52
R184 VDD.n434 VDD.t186 249.387
R185 VDD.n17 VDD.t189 249.363
R186 VDD.n27 VDD.t207 249.363
R187 VDD.n363 VDD.t191 249.363
R188 VDD.n368 VDD.t209 249.363
R189 VDD.n352 VDD.t9 249.363
R190 VDD.n340 VDD.t107 249.363
R191 VDD.n88 VDD.t68 249.362
R192 VDD.n93 VDD.t35 249.362
R193 VDD.n98 VDD.t148 249.362
R194 VDD.n103 VDD.t94 249.362
R195 VDD.n79 VDD.t46 249.362
R196 VDD.n122 VDD.t85 249.362
R197 VDD.n127 VDD.t206 249.362
R198 VDD.n132 VDD.t98 249.362
R199 VDD.n162 VDD.t1 249.362
R200 VDD.n157 VDD.t58 249.362
R201 VDD.n154 VDD.t3 249.362
R202 VDD.n149 VDD.t162 249.362
R203 VDD.n17 VDD.t21 249.362
R204 VDD.n27 VDD.t181 249.362
R205 VDD.n406 VDD.t50 249.362
R206 VDD.n388 VDD.t83 249.062
R207 VDD.n324 VDD.t24 249.062
R208 VDD.n399 VDD.t168 248.929
R209 VDD.t67 VDD.t37 248.599
R210 VDD.t34 VDD.t102 248.599
R211 VDD.t147 VDD.t14 248.599
R212 VDD.t93 VDD.t104 248.599
R213 VDD.t45 VDD.t90 248.599
R214 VDD.t84 VDD.t155 248.599
R215 VDD.t205 VDD.t6 248.599
R216 VDD.t97 VDD.t141 248.599
R217 VDD.t59 VDD.t0 248.599
R218 VDD.t177 VDD.t57 248.599
R219 VDD.t165 VDD.t2 248.599
R220 VDD.t113 VDD.t161 248.599
R221 VDD.t169 VDD.t63 248.599
R222 VDD.t175 VDD.t173 248.599
R223 VDD.t198 VDD.t200 248.599
R224 VDD.t53 VDD.t51 248.599
R225 VDD.t121 VDD.t119 248.599
R226 VDD.t137 VDD.t212 248.599
R227 VDD.t39 VDD.t41 248.599
R228 VDD.t115 VDD.t117 248.599
R229 VDD.t135 VDD.t133 248.599
R230 VDD.t214 VDD.t16 248.599
R231 VDD.t192 VDD.t163 248.599
R232 VDD.t194 VDD.t196 248.599
R233 VDD.t145 VDD.t153 248.599
R234 VDD.t12 VDD.t10 248.599
R235 VDD.t95 VDD.t100 248.599
R236 VDD.t126 VDD.t223 248.599
R237 VDD.t65 VDD.t32 248.599
R238 VDD.t75 VDD.t73 248.599
R239 VDD.t182 VDD.t184 248.599
R240 VDD.t18 VDD.t71 248.599
R241 VDD.t106 VDD.t187 248.599
R242 VDD.t8 VDD.t143 248.599
R243 VDD.t87 VDD.t208 248.599
R244 VDD.t29 VDD.t190 248.599
R245 VDD.n20 VDD.t89 247.394
R246 VDD.n25 VDD.t158 247.394
R247 VDD.n335 VDD.t30 247.394
R248 VDD.n364 VDD.t88 247.394
R249 VDD.n337 VDD.t144 247.394
R250 VDD.n351 VDD.t188 247.394
R251 VDD.n388 VDD.t28 247.394
R252 VDD.n324 VDD.t109 247.394
R253 VDD.n92 VDD.t38 247.394
R254 VDD.n97 VDD.t103 247.394
R255 VDD.n102 VDD.t15 247.394
R256 VDD.n80 VDD.t105 247.394
R257 VDD.n121 VDD.t91 247.394
R258 VDD.n126 VDD.t156 247.394
R259 VDD.n131 VDD.t7 247.394
R260 VDD.n113 VDD.t142 247.394
R261 VDD.n137 VDD.t60 247.394
R262 VDD.n155 VDD.t178 247.394
R263 VDD.n141 VDD.t166 247.394
R264 VDD.n147 VDD.t114 247.394
R265 VDD.n20 VDD.t218 247.394
R266 VDD.n25 VDD.t22 247.394
R267 VDD.n31 VDD.t31 247.394
R268 VDD.n404 VDD.t48 247.394
R269 VDD.n393 VDD.t140 245.178
R270 VDD.n322 VDD.t125 245.178
R271 VDD.n407 VDD.t112 245.178
R272 VDD.n8 VDD.t86 245.178
R273 VDD.n373 VDD.t172 243.512
R274 VDD.n344 VDD.t204 243.512
R275 VDD.n394 VDD.t81 243.508
R276 VDD.n387 VDD 230.766
R277 VDD.n194 VDD 221.964
R278 VDD.n217 VDD 221.964
R279 VDD.n218 VDD 221.964
R280 VDD.n241 VDD 221.964
R281 VDD.n242 VDD 221.964
R282 VDD.n265 VDD 221.964
R283 VDD.n266 VDD 221.964
R284 VDD.n289 VDD 221.964
R285 VDD.n290 VDD 221.964
R286 VDD.n111 VDD 219.004
R287 VDD VDD.n172 219.004
R288 VDD.n381 VDD 219.004
R289 VDD.n400 VDD.n399 213.119
R290 VDD.n413 VDD.n312 213.119
R291 VDD.n195 VDD.n194 213.119
R292 VDD.n217 VDD.n216 213.119
R293 VDD.n219 VDD.n218 213.119
R294 VDD.n241 VDD.n240 213.119
R295 VDD.n243 VDD.n242 213.119
R296 VDD.n265 VDD.n264 213.119
R297 VDD.n267 VDD.n266 213.119
R298 VDD.n289 VDD.n288 213.119
R299 VDD.n291 VDD.n290 213.119
R300 VDD.n381 VDD.n380 213.119
R301 VDD.t203 VDD.t110 213.084
R302 VDD.t149 VDD.t171 213.084
R303 VDD.n402 VDD.n401 209.368
R304 VDD.n417 VDD.n416 209.368
R305 VDD.t37 VDD 207.166
R306 VDD.t102 VDD 207.166
R307 VDD.t14 VDD 207.166
R308 VDD.t104 VDD 207.166
R309 VDD.t90 VDD 207.166
R310 VDD.t155 VDD 207.166
R311 VDD.t6 VDD 207.166
R312 VDD.t141 VDD 207.166
R313 VDD VDD.t59 207.166
R314 VDD VDD.t177 207.166
R315 VDD VDD.t165 207.166
R316 VDD VDD.t113 207.166
R317 VDD.t187 VDD 207.166
R318 VDD.t143 VDD 207.166
R319 VDD VDD.t87 207.166
R320 VDD VDD.t29 207.166
R321 VDD.t49 VDD 206.45
R322 VDD VDD.t169 198.287
R323 VDD VDD.t175 198.287
R324 VDD.t200 VDD 198.287
R325 VDD.t51 VDD 198.287
R326 VDD VDD.t121 198.287
R327 VDD VDD.t137 198.287
R328 VDD.t41 VDD 198.287
R329 VDD.t117 VDD 198.287
R330 VDD VDD.t135 198.287
R331 VDD VDD.t214 198.287
R332 VDD.t163 VDD 198.287
R333 VDD.t196 VDD 198.287
R334 VDD VDD.t145 198.287
R335 VDD VDD.t12 198.287
R336 VDD.t100 VDD 198.287
R337 VDD.t223 VDD 198.287
R338 VDD VDD.t65 198.287
R339 VDD VDD.t75 198.287
R340 VDD.t184 VDD 198.287
R341 VDD.t71 VDD 198.287
R342 VDD.t110 VDD 189.409
R343 VDD VDD.t149 189.409
R344 VDD.t129 VDD 177.916
R345 VDD.t61 VDD.t179 140.989
R346 VDD.t47 VDD.t49 140.989
R347 VDD.t80 VDD.t167 140.989
R348 VDD.t43 VDD.t124 134.276
R349 VDD.t219 VDD.t108 134.276
R350 VDD.t139 VDD.t221 134.276
R351 VDD.t27 VDD.t151 134.276
R352 VDD VDD.n417 125.883
R353 VDD VDD.n400 124.206
R354 VDD VDD.t111 107.421
R355 VDD VDD.t159 107.421
R356 VDD.t23 VDD 107.421
R357 VDD VDD.t82 107.421
R358 VDD.t179 VDD.n312 100.707
R359 VDD.n401 VDD.t43 100.707
R360 VDD VDD.t4 97.3503
R361 VDD.n417 VDD.t216 93.9934
R362 VDD VDD.t25 90.6365
R363 VDD.n400 VDD.t167 80.5659
R364 VDD.n15 VDD.n4 76.0729
R365 VDD.n5 VDD.n1 76.0729
R366 VDD.n438 VDD.n437 76.0729
R367 VDD.n435 VDD.n434 76.0729
R368 VDD.n15 VDD.n14 76.0728
R369 VDD.n12 VDD.n1 76.0728
R370 VDD.n438 VDD.n2 76.0728
R371 VDD.t55 VDD.t61 72.1736
R372 VDD.t221 VDD 70.4952
R373 VDD.t111 VDD.t55 68.8168
R374 VDD.t210 VDD 67.1383
R375 VDD.n312 VDD.t216 60.4245
R376 VDD.n401 VDD.t210 60.4245
R377 VDD.n163 VDD.n112 51.3536
R378 VDD.n172 VDD.n171 51.3536
R379 VDD.n174 VDD.n173 51.3536
R380 VDD.n111 VDD.n110 51.3536
R381 VDD.n11 VDD 48.6651
R382 VDD.n423 VDD.n422 43.9358
R383 VDD.t159 VDD 43.6401
R384 VDD.n10 VDD.t79 38.4155
R385 VDD.n40 VDD.t123 38.4155
R386 VDD.n429 VDD.t150 38.4155
R387 VDD.n317 VDD.t157 38.4155
R388 VDD.n436 VDD 36.603
R389 VDD.n423 VDD.n47 34.6358
R390 VDD.n427 VDD.n47 34.6358
R391 VDD.n428 VDD.n427 34.6358
R392 VDD.n369 VDD.n357 34.6358
R393 VDD.n376 VDD.n336 34.6358
R394 VDD.n346 VDD.n345 34.6358
R395 VDD.n309 VDD.n304 34.6358
R396 VDD.n416 VDD.n305 34.6358
R397 VDD.n402 VDD.n322 33.5064
R398 VDD.n33 VDD.n32 33.1299
R399 VDD.n394 VDD.n393 33.1299
R400 VDD.n146 VDD.n144 32.4116
R401 VDD.n389 VDD.n333 30.8711
R402 VDD.n329 VDD.n328 30.8711
R403 VDD.n41 VDD.n6 27.4829
R404 VDD.n430 VDD.n428 27.4829
R405 VDD.t25 VDD.t80 26.8556
R406 VDD.n10 VDD.t128 26.5955
R407 VDD.n40 VDD.t132 26.5955
R408 VDD.n429 VDD.t99 26.5955
R409 VDD.n332 VDD.t222 26.5955
R410 VDD.n332 VDD.t152 26.5955
R411 VDD.n326 VDD.t44 26.5955
R412 VDD.n326 VDD.t220 26.5955
R413 VDD.n313 VDD.t180 26.5955
R414 VDD.n313 VDD.t62 26.5955
R415 VDD.n317 VDD.t5 26.5955
R416 VDD.n88 VDD.n84 25.977
R417 VDD.n93 VDD.n83 25.977
R418 VDD.n98 VDD.n82 25.977
R419 VDD.n104 VDD.n103 25.977
R420 VDD.n117 VDD.n79 25.977
R421 VDD.n122 VDD.n116 25.977
R422 VDD.n127 VDD.n115 25.977
R423 VDD.n133 VDD.n132 25.977
R424 VDD.n162 VDD.n161 25.977
R425 VDD.n157 VDD.n156 25.977
R426 VDD.n154 VDD.n153 25.977
R427 VDD.n149 VDD.n148 25.977
R428 VDD.n21 VDD.n17 25.977
R429 VDD.n27 VDD.n26 25.977
R430 VDD.n38 VDD.n37 25.977
R431 VDD.n363 VDD.n359 25.977
R432 VDD.n368 VDD.n358 25.977
R433 VDD.n353 VDD.n352 25.977
R434 VDD.n350 VDD.n340 25.977
R435 VDD.n298 VDD.n297 25.224
R436 VDD.n299 VDD.n298 25.224
R437 VDD.n295 VDD.n51 25.224
R438 VDD.n296 VDD.n295 25.224
R439 VDD.n282 VDD.n278 25.224
R440 VDD.n278 VDD.n52 25.224
R441 VDD.n284 VDD.n53 25.224
R442 VDD.n284 VDD.n283 25.224
R443 VDD.n274 VDD.n273 25.224
R444 VDD.n274 VDD.n54 25.224
R445 VDD.n271 VDD.n57 25.224
R446 VDD.n272 VDD.n271 25.224
R447 VDD.n258 VDD.n254 25.224
R448 VDD.n254 VDD.n58 25.224
R449 VDD.n260 VDD.n59 25.224
R450 VDD.n260 VDD.n259 25.224
R451 VDD.n250 VDD.n249 25.224
R452 VDD.n250 VDD.n60 25.224
R453 VDD.n247 VDD.n63 25.224
R454 VDD.n248 VDD.n247 25.224
R455 VDD.n234 VDD.n230 25.224
R456 VDD.n230 VDD.n64 25.224
R457 VDD.n236 VDD.n65 25.224
R458 VDD.n236 VDD.n235 25.224
R459 VDD.n226 VDD.n225 25.224
R460 VDD.n226 VDD.n66 25.224
R461 VDD.n223 VDD.n69 25.224
R462 VDD.n224 VDD.n223 25.224
R463 VDD.n210 VDD.n206 25.224
R464 VDD.n206 VDD.n70 25.224
R465 VDD.n212 VDD.n71 25.224
R466 VDD.n212 VDD.n211 25.224
R467 VDD.n202 VDD.n201 25.224
R468 VDD.n202 VDD.n72 25.224
R469 VDD.n199 VDD.n75 25.224
R470 VDD.n200 VDD.n199 25.224
R471 VDD.n187 VDD.n183 25.224
R472 VDD.n183 VDD.n76 25.224
R473 VDD.n189 VDD.n77 25.224
R474 VDD.n189 VDD.n188 25.224
R475 VDD.n87 VDD.n86 25.1591
R476 VDD.n109 VDD.n108 25.1591
R477 VDD.n176 VDD.n175 25.1591
R478 VDD.n170 VDD.n169 25.1591
R479 VDD.n165 VDD.n164 25.1591
R480 VDD.n92 VDD.n84 24.4711
R481 VDD.n97 VDD.n83 24.4711
R482 VDD.n102 VDD.n82 24.4711
R483 VDD.n104 VDD.n80 24.4711
R484 VDD.n121 VDD.n117 24.4711
R485 VDD.n126 VDD.n116 24.4711
R486 VDD.n131 VDD.n115 24.4711
R487 VDD.n133 VDD.n113 24.4711
R488 VDD.n161 VDD.n137 24.4711
R489 VDD.n156 VDD.n155 24.4711
R490 VDD.n153 VDD.n141 24.4711
R491 VDD.n148 VDD.n147 24.4711
R492 VDD.n21 VDD.n20 24.4711
R493 VDD.n26 VDD.n25 24.4711
R494 VDD.n32 VDD.n31 24.4711
R495 VDD.n359 VDD.n335 24.4711
R496 VDD.n364 VDD.n358 24.4711
R497 VDD.n374 VDD.n373 24.4711
R498 VDD.n353 VDD.n337 24.4711
R499 VDD.n351 VDD.n350 24.4711
R500 VDD.n389 VDD.n388 24.4711
R501 VDD.n412 VDD.n411 24.4711
R502 VDD.n329 VDD.n324 24.4711
R503 VDD.n434 VDD.n6 23.7181
R504 VDD.n434 VDD.n433 23.7181
R505 VDD.n369 VDD.n368 23.7181
R506 VDD.n380 VDD.n336 23.7181
R507 VDD.n346 VDD.n340 23.7181
R508 VDD.n418 VDD.n304 23.7181
R509 VDD.n37 VDD.n8 22.9652
R510 VDD.n395 VDD.n323 22.9652
R511 VDD.n403 VDD.n402 22.9652
R512 VDD.n413 VDD.n306 22.5887
R513 VDD.n407 VDD.n406 22.5887
R514 VDD.n13 VDD.t69 21.2133
R515 VDD.t20 VDD.n3 21.2133
R516 VDD.n413 VDD.n412 21.0829
R517 VDD.n297 VDD.n296 20.3299
R518 VDD.n283 VDD.n282 20.3299
R519 VDD.n273 VDD.n272 20.3299
R520 VDD.n259 VDD.n258 20.3299
R521 VDD.n249 VDD.n248 20.3299
R522 VDD.n235 VDD.n234 20.3299
R523 VDD.n225 VDD.n224 20.3299
R524 VDD.n211 VDD.n210 20.3299
R525 VDD.n201 VDD.n200 20.3299
R526 VDD.n188 VDD.n187 20.3299
R527 VDD.t4 VDD.t47 20.1418
R528 VDD.n373 VDD.n357 19.9534
R529 VDD.n345 VDD.n344 19.9534
R530 VDD.n406 VDD.n405 18.824
R531 VDD.n411 VDD.n315 18.4476
R532 VDD.t69 VDD.n11 17.4699
R533 VDD.n436 VDD.t20 17.4699
R534 VDD.n291 VDD.n51 17.3181
R535 VDD.n288 VDD.n53 17.3181
R536 VDD.n267 VDD.n57 17.3181
R537 VDD.n264 VDD.n59 17.3181
R538 VDD.n243 VDD.n63 17.3181
R539 VDD.n240 VDD.n65 17.3181
R540 VDD.n219 VDD.n69 17.3181
R541 VDD.n216 VDD.n71 17.3181
R542 VDD.n195 VDD.n75 17.3181
R543 VDD.n193 VDD.n77 17.3181
R544 VDD.n408 VDD.n315 16.1887
R545 VDD.n291 VDD.n52 15.8123
R546 VDD.n288 VDD.n54 15.8123
R547 VDD.n267 VDD.n58 15.8123
R548 VDD.n264 VDD.n60 15.8123
R549 VDD.n243 VDD.n64 15.8123
R550 VDD.n240 VDD.n66 15.8123
R551 VDD.n219 VDD.n70 15.8123
R552 VDD.n216 VDD.n72 15.8123
R553 VDD.n195 VDD.n76 15.8123
R554 VDD.n86 VDD 15.0074
R555 VDD.n109 VDD 15.0074
R556 VDD.n175 VDD 15.0074
R557 VDD.n170 VDD 15.0074
R558 VDD.n164 VDD 15.0074
R559 VDD.n399 VDD.n323 14.3064
R560 VDD.n405 VDD.n404 14.3064
R561 VDD.n404 VDD.n403 14.3064
R562 VDD.n344 VDD.n343 13.5534
R563 VDD.n88 VDD.n87 12.8005
R564 VDD.n93 VDD.n92 12.8005
R565 VDD.n98 VDD.n97 12.8005
R566 VDD.n103 VDD.n102 12.8005
R567 VDD.n108 VDD.n80 12.8005
R568 VDD.n176 VDD.n79 12.8005
R569 VDD.n122 VDD.n121 12.8005
R570 VDD.n127 VDD.n126 12.8005
R571 VDD.n132 VDD.n131 12.8005
R572 VDD.n169 VDD.n113 12.8005
R573 VDD.n165 VDD.n162 12.8005
R574 VDD.n157 VDD.n137 12.8005
R575 VDD.n155 VDD.n154 12.8005
R576 VDD.n149 VDD.n141 12.8005
R577 VDD.n147 VDD.n146 12.8005
R578 VDD.n438 VDD.n1 12.8005
R579 VDD.n20 VDD.n1 12.8005
R580 VDD.n25 VDD.n17 12.8005
R581 VDD.n27 VDD.n15 12.8005
R582 VDD.n31 VDD.n15 12.8005
R583 VDD.n382 VDD.n335 12.8005
R584 VDD.n364 VDD.n363 12.8005
R585 VDD.n380 VDD.n337 12.8005
R586 VDD.n352 VDD.n351 12.8005
R587 VDD.n388 VDD.n387 12.8005
R588 VDD.n399 VDD.n324 12.8005
R589 VDD.n179 VDD.n178 11.6828
R590 VDD.n167 VDD.n78 11.6828
R591 VDD.n376 VDD.n375 10.5417
R592 VDD.n309 VDD.n308 10.5417
R593 VDD VDD.n442 9.39425
R594 VDD.n87 VDD 9.32654
R595 VDD.n146 VDD.n145 9.3005
R596 VDD.n147 VDD.n143 9.3005
R597 VDD.n148 VDD.n142 9.3005
R598 VDD.n150 VDD.n149 9.3005
R599 VDD.n151 VDD.n141 9.3005
R600 VDD.n153 VDD.n152 9.3005
R601 VDD.n154 VDD.n140 9.3005
R602 VDD.n155 VDD.n139 9.3005
R603 VDD.n156 VDD.n138 9.3005
R604 VDD.n158 VDD.n157 9.3005
R605 VDD.n159 VDD.n137 9.3005
R606 VDD.n161 VDD.n160 9.3005
R607 VDD.n162 VDD.n136 9.3005
R608 VDD.n166 VDD.n165 9.3005
R609 VDD.n169 VDD.n168 9.3005
R610 VDD.n135 VDD.n113 9.3005
R611 VDD.n134 VDD.n133 9.3005
R612 VDD.n132 VDD.n114 9.3005
R613 VDD.n131 VDD.n130 9.3005
R614 VDD.n129 VDD.n115 9.3005
R615 VDD.n128 VDD.n127 9.3005
R616 VDD.n126 VDD.n125 9.3005
R617 VDD.n124 VDD.n116 9.3005
R618 VDD.n123 VDD.n122 9.3005
R619 VDD.n121 VDD.n120 9.3005
R620 VDD.n119 VDD.n117 9.3005
R621 VDD.n118 VDD.n79 9.3005
R622 VDD.n177 VDD.n176 9.3005
R623 VDD.n108 VDD.n107 9.3005
R624 VDD.n106 VDD.n80 9.3005
R625 VDD.n105 VDD.n104 9.3005
R626 VDD.n103 VDD.n81 9.3005
R627 VDD.n102 VDD.n101 9.3005
R628 VDD.n100 VDD.n82 9.3005
R629 VDD.n99 VDD.n98 9.3005
R630 VDD.n97 VDD.n96 9.3005
R631 VDD.n95 VDD.n83 9.3005
R632 VDD.n94 VDD.n93 9.3005
R633 VDD.n92 VDD.n91 9.3005
R634 VDD.n90 VDD.n84 9.3005
R635 VDD.n89 VDD.n88 9.3005
R636 VDD.n343 VDD.n303 9.3005
R637 VDD.n344 VDD.n342 9.3005
R638 VDD.n348 VDD.n340 9.3005
R639 VDD.n351 VDD.n339 9.3005
R640 VDD.n352 VDD.n338 9.3005
R641 VDD.n355 VDD.n337 9.3005
R642 VDD.n380 VDD.n379 9.3005
R643 VDD.n373 VDD.n372 9.3005
R644 VDD.n368 VDD.n367 9.3005
R645 VDD.n365 VDD.n364 9.3005
R646 VDD.n363 VDD.n362 9.3005
R647 VDD.n360 VDD.n335 9.3005
R648 VDD.n383 VDD.n382 9.3005
R649 VDD.n361 VDD.n359 9.3005
R650 VDD.n366 VDD.n358 9.3005
R651 VDD.n370 VDD.n369 9.3005
R652 VDD.n371 VDD.n357 9.3005
R653 VDD.n374 VDD.n356 9.3005
R654 VDD.n377 VDD.n376 9.3005
R655 VDD.n378 VDD.n336 9.3005
R656 VDD.n354 VDD.n353 9.3005
R657 VDD.n350 VDD.n349 9.3005
R658 VDD.n347 VDD.n346 9.3005
R659 VDD.n345 VDD.n341 9.3005
R660 VDD.n419 VDD.n418 9.3005
R661 VDD.n416 VDD.n415 9.3005
R662 VDD.n409 VDD.n408 9.3005
R663 VDD.n405 VDD.n318 9.3005
R664 VDD.n403 VDD.n320 9.3005
R665 VDD.n402 VDD.n321 9.3005
R666 VDD.n327 VDD.n325 9.3005
R667 VDD.n331 VDD.n324 9.3005
R668 VDD.n399 VDD.n398 9.3005
R669 VDD.n396 VDD.n395 9.3005
R670 VDD.n392 VDD.n391 9.3005
R671 VDD.n388 VDD.n334 9.3005
R672 VDD.n387 VDD.n386 9.3005
R673 VDD.n390 VDD.n389 9.3005
R674 VDD.n397 VDD.n323 9.3005
R675 VDD.n330 VDD.n329 9.3005
R676 VDD.n404 VDD.n319 9.3005
R677 VDD.n406 VDD.n316 9.3005
R678 VDD.n411 VDD.n410 9.3005
R679 VDD.n412 VDD.n314 9.3005
R680 VDD.n414 VDD.n413 9.3005
R681 VDD.n311 VDD.n305 9.3005
R682 VDD.n310 VDD.n309 9.3005
R683 VDD.n307 VDD.n304 9.3005
R684 VDD.n431 VDD.n430 9.3005
R685 VDD.n434 VDD.n44 9.3005
R686 VDD.n35 VDD.n34 9.3005
R687 VDD.n31 VDD.n30 9.3005
R688 VDD.n29 VDD.n15 9.3005
R689 VDD.n28 VDD.n27 9.3005
R690 VDD.n25 VDD.n24 9.3005
R691 VDD.n23 VDD.n17 9.3005
R692 VDD.n20 VDD.n19 9.3005
R693 VDD.n18 VDD.n1 9.3005
R694 VDD.n439 VDD.n438 9.3005
R695 VDD.n22 VDD.n21 9.3005
R696 VDD.n26 VDD.n16 9.3005
R697 VDD.n32 VDD.n9 9.3005
R698 VDD.n37 VDD.n36 9.3005
R699 VDD.n38 VDD.n7 9.3005
R700 VDD.n42 VDD.n41 9.3005
R701 VDD.n43 VDD.n6 9.3005
R702 VDD.n433 VDD.n432 9.3005
R703 VDD.n428 VDD.n46 9.3005
R704 VDD.n427 VDD.n426 9.3005
R705 VDD.n425 VDD.n47 9.3005
R706 VDD.n424 VDD.n423 9.3005
R707 VDD.n193 VDD.n192 9.3005
R708 VDD.n188 VDD.n182 9.3005
R709 VDD.n184 VDD.n76 9.3005
R710 VDD.n196 VDD.n195 9.3005
R711 VDD.n200 VDD.n74 9.3005
R712 VDD.n204 VDD.n72 9.3005
R713 VDD.n216 VDD.n215 9.3005
R714 VDD.n211 VDD.n205 9.3005
R715 VDD.n207 VDD.n70 9.3005
R716 VDD.n220 VDD.n219 9.3005
R717 VDD.n224 VDD.n68 9.3005
R718 VDD.n228 VDD.n66 9.3005
R719 VDD.n240 VDD.n239 9.3005
R720 VDD.n235 VDD.n229 9.3005
R721 VDD.n231 VDD.n64 9.3005
R722 VDD.n244 VDD.n243 9.3005
R723 VDD.n248 VDD.n62 9.3005
R724 VDD.n252 VDD.n60 9.3005
R725 VDD.n264 VDD.n263 9.3005
R726 VDD.n259 VDD.n253 9.3005
R727 VDD.n255 VDD.n58 9.3005
R728 VDD.n268 VDD.n267 9.3005
R729 VDD.n272 VDD.n56 9.3005
R730 VDD.n276 VDD.n54 9.3005
R731 VDD.n288 VDD.n287 9.3005
R732 VDD.n283 VDD.n277 9.3005
R733 VDD.n279 VDD.n52 9.3005
R734 VDD.n292 VDD.n291 9.3005
R735 VDD.n296 VDD.n50 9.3005
R736 VDD.n300 VDD.n299 9.3005
R737 VDD.n298 VDD.n48 9.3005
R738 VDD.n297 VDD.n49 9.3005
R739 VDD.n295 VDD.n294 9.3005
R740 VDD.n293 VDD.n51 9.3005
R741 VDD.n280 VDD.n278 9.3005
R742 VDD.n282 VDD.n281 9.3005
R743 VDD.n285 VDD.n284 9.3005
R744 VDD.n286 VDD.n53 9.3005
R745 VDD.n275 VDD.n274 9.3005
R746 VDD.n273 VDD.n55 9.3005
R747 VDD.n271 VDD.n270 9.3005
R748 VDD.n269 VDD.n57 9.3005
R749 VDD.n256 VDD.n254 9.3005
R750 VDD.n258 VDD.n257 9.3005
R751 VDD.n261 VDD.n260 9.3005
R752 VDD.n262 VDD.n59 9.3005
R753 VDD.n251 VDD.n250 9.3005
R754 VDD.n249 VDD.n61 9.3005
R755 VDD.n247 VDD.n246 9.3005
R756 VDD.n245 VDD.n63 9.3005
R757 VDD.n232 VDD.n230 9.3005
R758 VDD.n234 VDD.n233 9.3005
R759 VDD.n237 VDD.n236 9.3005
R760 VDD.n238 VDD.n65 9.3005
R761 VDD.n227 VDD.n226 9.3005
R762 VDD.n225 VDD.n67 9.3005
R763 VDD.n223 VDD.n222 9.3005
R764 VDD.n221 VDD.n69 9.3005
R765 VDD.n208 VDD.n206 9.3005
R766 VDD.n210 VDD.n209 9.3005
R767 VDD.n213 VDD.n212 9.3005
R768 VDD.n214 VDD.n71 9.3005
R769 VDD.n203 VDD.n202 9.3005
R770 VDD.n201 VDD.n73 9.3005
R771 VDD.n199 VDD.n198 9.3005
R772 VDD.n197 VDD.n75 9.3005
R773 VDD.n185 VDD.n183 9.3005
R774 VDD.n187 VDD.n186 9.3005
R775 VDD.n190 VDD.n189 9.3005
R776 VDD.n191 VDD.n77 9.3005
R777 VDD.n39 VDD.n38 8.28285
R778 VDD.n433 VDD.n45 8.28285
R779 VDD.n375 VDD.n374 8.28285
R780 VDD.n308 VDD.n305 8.28285
R781 VDD.n144 VDD 7.34877
R782 VDD.t124 VDD.t219 6.71428
R783 VDD.t108 VDD.t23 6.71428
R784 VDD.t151 VDD.t139 6.71428
R785 VDD.t82 VDD.t27 6.71428
R786 VDD.n180 VDD.n179 6.09998
R787 VDD.n441 VDD.n440 4.33704
R788 VDD VDD.n302 4.10787
R789 VDD.n420 VDD.n303 3.76683
R790 VDD.n392 VDD.n333 3.76521
R791 VDD.n328 VDD.n327 3.76521
R792 VDD.n384 VDD 3.09034
R793 VDD VDD.n385 3.09034
R794 VDD.n440 VDD 3.09034
R795 VDD.n420 VDD.n419 2.89503
R796 VDD.n422 VDD.n421 2.89503
R797 VDD.n181 VDD.n180 2.34946
R798 VDD.n301 VDD.n0 2.34946
R799 VDD.n302 VDD 2.27784
R800 VDD.n442 VDD.n0 2.24112
R801 VDD.n302 VDD.n301 2.16789
R802 VDD.n181 VDD.n78 1.91476
R803 VDD.n442 VDD.n441 1.82316
R804 VDD.n180 VDD.n0 1.73404
R805 VDD.n34 VDD.n33 1.50638
R806 VDD.n34 VDD.n8 1.12991
R807 VDD.n393 VDD.n392 1.12991
R808 VDD.n416 VDD.n306 1.12991
R809 VDD.n408 VDD.n407 1.12991
R810 VDD.n327 VDD.n322 1.12991
R811 VDD.n179 VDD.n78 1.12238
R812 VDD.n421 VDD.n420 0.872295
R813 VDD.n385 VDD.n384 0.872295
R814 VDD.n301 VDD 0.647576
R815 VDD.n192 VDD.n181 0.643669
R816 VDD.n440 VDD 0.462038
R817 VDD.n385 VDD 0.410756
R818 VDD.n41 VDD.n39 0.376971
R819 VDD.n430 VDD.n45 0.376971
R820 VDD.n395 VDD.n394 0.376971
R821 VDD.n441 VDD 0.302844
R822 VDD.n421 VDD 0.229667
R823 VDD.n90 VDD.n89 0.120292
R824 VDD.n91 VDD.n90 0.120292
R825 VDD.n95 VDD.n94 0.120292
R826 VDD.n96 VDD.n95 0.120292
R827 VDD.n100 VDD.n99 0.120292
R828 VDD.n101 VDD.n100 0.120292
R829 VDD.n105 VDD.n81 0.120292
R830 VDD.n106 VDD.n105 0.120292
R831 VDD.n119 VDD.n118 0.120292
R832 VDD.n120 VDD.n119 0.120292
R833 VDD.n124 VDD.n123 0.120292
R834 VDD.n125 VDD.n124 0.120292
R835 VDD.n129 VDD.n128 0.120292
R836 VDD.n130 VDD.n129 0.120292
R837 VDD.n134 VDD.n114 0.120292
R838 VDD.n135 VDD.n134 0.120292
R839 VDD.n160 VDD.n136 0.120292
R840 VDD.n160 VDD.n159 0.120292
R841 VDD.n158 VDD.n138 0.120292
R842 VDD.n139 VDD.n138 0.120292
R843 VDD.n152 VDD.n140 0.120292
R844 VDD.n152 VDD.n151 0.120292
R845 VDD.n150 VDD.n142 0.120292
R846 VDD.n143 VDD.n142 0.120292
R847 VDD.n342 VDD.n341 0.120292
R848 VDD.n347 VDD.n341 0.120292
R849 VDD.n349 VDD.n348 0.120292
R850 VDD.n349 VDD.n339 0.120292
R851 VDD.n354 VDD.n338 0.120292
R852 VDD.n355 VDD.n354 0.120292
R853 VDD.n378 VDD.n377 0.120292
R854 VDD.n377 VDD.n356 0.120292
R855 VDD.n372 VDD.n371 0.120292
R856 VDD.n371 VDD.n370 0.120292
R857 VDD.n367 VDD.n366 0.120292
R858 VDD.n366 VDD.n365 0.120292
R859 VDD.n362 VDD.n361 0.120292
R860 VDD.n361 VDD.n360 0.120292
R861 VDD.n310 VDD.n307 0.120292
R862 VDD.n311 VDD.n310 0.120292
R863 VDD.n410 VDD.n314 0.120292
R864 VDD.n410 VDD.n409 0.120292
R865 VDD.n318 VDD.n316 0.120292
R866 VDD.n319 VDD.n318 0.120292
R867 VDD.n330 VDD.n325 0.120292
R868 VDD.n331 VDD.n330 0.120292
R869 VDD.n397 VDD.n396 0.120292
R870 VDD.n391 VDD.n390 0.120292
R871 VDD.n390 VDD.n334 0.120292
R872 VDD.n425 VDD.n424 0.120292
R873 VDD.n426 VDD.n425 0.120292
R874 VDD.n431 VDD.n46 0.120292
R875 VDD.n432 VDD.n431 0.120292
R876 VDD.n43 VDD.n42 0.120292
R877 VDD.n42 VDD.n7 0.120292
R878 VDD.n35 VDD.n9 0.120292
R879 VDD.n30 VDD.n9 0.120292
R880 VDD.n28 VDD.n16 0.120292
R881 VDD.n24 VDD.n16 0.120292
R882 VDD.n23 VDD.n22 0.120292
R883 VDD.n22 VDD.n19 0.120292
R884 VDD VDD.n177 0.11899
R885 VDD VDD.n166 0.11899
R886 VDD.n424 VDD 0.109875
R887 VDD VDD.n46 0.104667
R888 VDD VDD.n167 0.09425
R889 VDD.n178 VDD 0.078625
R890 VDD.n191 VDD.n190 0.072375
R891 VDD.n190 VDD.n182 0.072375
R892 VDD.n186 VDD.n185 0.072375
R893 VDD.n185 VDD.n184 0.072375
R894 VDD.n198 VDD.n197 0.072375
R895 VDD.n198 VDD.n74 0.072375
R896 VDD.n203 VDD.n73 0.072375
R897 VDD.n204 VDD.n203 0.072375
R898 VDD.n214 VDD.n213 0.072375
R899 VDD.n213 VDD.n205 0.072375
R900 VDD.n209 VDD.n208 0.072375
R901 VDD.n208 VDD.n207 0.072375
R902 VDD.n222 VDD.n221 0.072375
R903 VDD.n222 VDD.n68 0.072375
R904 VDD.n227 VDD.n67 0.072375
R905 VDD.n228 VDD.n227 0.072375
R906 VDD.n238 VDD.n237 0.072375
R907 VDD.n237 VDD.n229 0.072375
R908 VDD.n233 VDD.n232 0.072375
R909 VDD.n232 VDD.n231 0.072375
R910 VDD.n246 VDD.n245 0.072375
R911 VDD.n246 VDD.n62 0.072375
R912 VDD.n251 VDD.n61 0.072375
R913 VDD.n252 VDD.n251 0.072375
R914 VDD.n262 VDD.n261 0.072375
R915 VDD.n261 VDD.n253 0.072375
R916 VDD.n257 VDD.n256 0.072375
R917 VDD.n256 VDD.n255 0.072375
R918 VDD.n270 VDD.n269 0.072375
R919 VDD.n270 VDD.n56 0.072375
R920 VDD.n275 VDD.n55 0.072375
R921 VDD.n276 VDD.n275 0.072375
R922 VDD.n286 VDD.n285 0.072375
R923 VDD.n285 VDD.n277 0.072375
R924 VDD.n281 VDD.n280 0.072375
R925 VDD.n280 VDD.n279 0.072375
R926 VDD.n294 VDD.n293 0.072375
R927 VDD.n294 VDD.n50 0.072375
R928 VDD.n49 VDD.n48 0.072375
R929 VDD.n300 VDD.n48 0.072375
R930 VDD.n89 VDD 0.0603958
R931 VDD.n94 VDD 0.0603958
R932 VDD.n99 VDD 0.0603958
R933 VDD VDD.n81 0.0603958
R934 VDD.n107 VDD 0.0603958
R935 VDD.n118 VDD 0.0603958
R936 VDD.n123 VDD 0.0603958
R937 VDD.n128 VDD 0.0603958
R938 VDD VDD.n114 0.0603958
R939 VDD.n168 VDD 0.0603958
R940 VDD.n136 VDD 0.0603958
R941 VDD VDD.n158 0.0603958
R942 VDD.n140 VDD 0.0603958
R943 VDD VDD.n150 0.0603958
R944 VDD.n145 VDD 0.0603958
R945 VDD.n342 VDD 0.0603958
R946 VDD.n348 VDD 0.0603958
R947 VDD VDD.n338 0.0603958
R948 VDD.n379 VDD 0.0603958
R949 VDD VDD.n378 0.0603958
R950 VDD.n372 VDD 0.0603958
R951 VDD.n367 VDD 0.0603958
R952 VDD.n362 VDD 0.0603958
R953 VDD.n383 VDD 0.0603958
R954 VDD.n307 VDD 0.0603958
R955 VDD.n415 VDD 0.0603958
R956 VDD VDD.n414 0.0603958
R957 VDD.n314 VDD 0.0603958
R958 VDD.n316 VDD 0.0603958
R959 VDD.n320 VDD 0.0603958
R960 VDD.n321 VDD 0.0603958
R961 VDD.n325 VDD 0.0603958
R962 VDD.n398 VDD 0.0603958
R963 VDD VDD.n397 0.0603958
R964 VDD.n391 VDD 0.0603958
R965 VDD.n386 VDD 0.0603958
R966 VDD VDD.n44 0.0603958
R967 VDD VDD.n43 0.0603958
R968 VDD.n36 VDD 0.0603958
R969 VDD VDD.n35 0.0603958
R970 VDD VDD.n29 0.0603958
R971 VDD VDD.n28 0.0603958
R972 VDD VDD.n23 0.0603958
R973 VDD VDD.n18 0.0603958
R974 VDD.n439 VDD 0.0603958
R975 VDD.n178 VDD 0.0408646
R976 VDD.n379 VDD 0.0382604
R977 VDD.n384 VDD 0.0365577
R978 VDD VDD.n191 0.0364375
R979 VDD.n186 VDD 0.0364375
R980 VDD.n196 VDD 0.0364375
R981 VDD.n197 VDD 0.0364375
R982 VDD VDD.n73 0.0364375
R983 VDD.n215 VDD 0.0364375
R984 VDD VDD.n214 0.0364375
R985 VDD.n209 VDD 0.0364375
R986 VDD.n220 VDD 0.0364375
R987 VDD.n221 VDD 0.0364375
R988 VDD VDD.n67 0.0364375
R989 VDD.n239 VDD 0.0364375
R990 VDD VDD.n238 0.0364375
R991 VDD.n233 VDD 0.0364375
R992 VDD.n244 VDD 0.0364375
R993 VDD.n245 VDD 0.0364375
R994 VDD VDD.n61 0.0364375
R995 VDD.n263 VDD 0.0364375
R996 VDD VDD.n262 0.0364375
R997 VDD.n257 VDD 0.0364375
R998 VDD.n268 VDD 0.0364375
R999 VDD.n269 VDD 0.0364375
R1000 VDD VDD.n55 0.0364375
R1001 VDD.n287 VDD 0.0364375
R1002 VDD VDD.n286 0.0364375
R1003 VDD.n281 VDD 0.0364375
R1004 VDD.n292 VDD 0.0364375
R1005 VDD.n293 VDD 0.0364375
R1006 VDD VDD.n49 0.0364375
R1007 VDD VDD.n303 0.03175
R1008 VDD VDD.n383 0.03175
R1009 VDD.n419 VDD 0.03175
R1010 VDD.n415 VDD 0.03175
R1011 VDD.n414 VDD 0.03175
R1012 VDD VDD.n321 0.03175
R1013 VDD.n398 VDD 0.03175
R1014 VDD.n386 VDD 0.03175
R1015 VDD.n29 VDD 0.03175
R1016 VDD.n18 VDD 0.03175
R1017 VDD VDD.n439 0.03175
R1018 VDD.n107 VDD 0.0265417
R1019 VDD.n177 VDD 0.0265417
R1020 VDD.n168 VDD 0.0265417
R1021 VDD.n166 VDD 0.0265417
R1022 VDD.n145 VDD 0.0265417
R1023 VDD.n167 VDD 0.0252396
R1024 VDD.n91 VDD 0.0239375
R1025 VDD.n96 VDD 0.0239375
R1026 VDD.n101 VDD 0.0239375
R1027 VDD VDD.n106 0.0239375
R1028 VDD.n120 VDD 0.0239375
R1029 VDD.n125 VDD 0.0239375
R1030 VDD.n130 VDD 0.0239375
R1031 VDD VDD.n135 0.0239375
R1032 VDD.n159 VDD 0.0239375
R1033 VDD VDD.n139 0.0239375
R1034 VDD.n151 VDD 0.0239375
R1035 VDD VDD.n143 0.0239375
R1036 VDD.n339 VDD 0.0239375
R1037 VDD VDD.n355 0.0239375
R1038 VDD.n365 VDD 0.0239375
R1039 VDD.n360 VDD 0.0239375
R1040 VDD VDD.n319 0.0239375
R1041 VDD.n396 VDD 0.0239375
R1042 VDD.n24 VDD 0.0239375
R1043 VDD.n19 VDD 0.0239375
R1044 VDD VDD.n356 0.0226354
R1045 VDD VDD.n311 0.0226354
R1046 VDD.n432 VDD 0.0226354
R1047 VDD VDD.n7 0.0226354
R1048 VDD VDD.n347 0.0213333
R1049 VDD.n370 VDD 0.0213333
R1050 VDD.n409 VDD 0.0213333
R1051 VDD VDD.n320 0.0213333
R1052 VDD VDD.n331 0.0213333
R1053 VDD VDD.n334 0.0213333
R1054 VDD.n44 VDD 0.0213333
R1055 VDD.n36 VDD 0.0213333
R1056 VDD.n30 VDD 0.0213333
R1057 VDD.n192 VDD 0.01925
R1058 VDD VDD.n196 0.01925
R1059 VDD.n215 VDD 0.01925
R1060 VDD VDD.n220 0.01925
R1061 VDD.n239 VDD 0.01925
R1062 VDD VDD.n244 0.01925
R1063 VDD.n263 VDD 0.01925
R1064 VDD VDD.n268 0.01925
R1065 VDD.n287 VDD 0.01925
R1066 VDD VDD.n292 0.01925
R1067 VDD.n426 VDD 0.016125
R1068 VDD VDD.n182 0.0137813
R1069 VDD.n184 VDD 0.0137813
R1070 VDD.n74 VDD 0.0137813
R1071 VDD VDD.n204 0.0137813
R1072 VDD VDD.n205 0.0137813
R1073 VDD.n207 VDD 0.0137813
R1074 VDD.n68 VDD 0.0137813
R1075 VDD VDD.n228 0.0137813
R1076 VDD VDD.n229 0.0137813
R1077 VDD.n231 VDD 0.0137813
R1078 VDD.n62 VDD 0.0137813
R1079 VDD VDD.n252 0.0137813
R1080 VDD VDD.n253 0.0137813
R1081 VDD.n255 VDD 0.0137813
R1082 VDD.n56 VDD 0.0137813
R1083 VDD VDD.n276 0.0137813
R1084 VDD VDD.n277 0.0137813
R1085 VDD.n279 VDD 0.0137813
R1086 VDD.n50 VDD 0.0137813
R1087 VDD VDD.n300 0.0137813
R1088 VDD.n422 VDD 0.0109167
R1089 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 593.154
R1090 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 231.554
R1091 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 140.53
R1092 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 26.5955
R1093 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 26.5955
R1094 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 16.5652
R1095 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 9.03579
R1096 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 6.02403
R1097 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 1.72748
R1098 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t5 230.363
R1099 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t9 230.155
R1100 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t6 229.369
R1101 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t7 212.081
R1102 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t13 212.081
R1103 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n0 203.923
R1104 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n3 186.001
R1105 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t4 158.064
R1106 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t11 157.856
R1107 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t10 157.07
R1108 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n8 155.058
R1109 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n11 154.91
R1110 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n5 152
R1111 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t12 139.78
R1112 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t8 139.78
R1113 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n16 101.49
R1114 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n2 61.346
R1115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n9 33.2524
R1116 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n13 29.6212
R1117 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t2 26.5955
R1118 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t3 26.5955
R1119 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t0 24.9236
R1120 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t1 24.9236
R1121 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n6 20.0252
R1122 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n12 18.1725
R1123 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n15 13.5685
R1124 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n1 10.7525
R1125 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n14 9.64425
R1126 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n4 9.30224
R1127 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 6.6565
R1128 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 5.92643
R1129 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 5.04292
R1130 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 3.8405
R1131 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 3.78232
R1132 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 3.0725
R1133 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 2.5605
R1134 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n7 2.17042
R1135 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n17 1.93989
R1136 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n10 1.93214
R1137 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 1.33781
R1138 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.490734
R1139 GND.n1582 GND.n1581 2.89982e+06
R1140 GND.n1581 GND.n1578 135084
R1141 GND.n1506 GND.n237 75097.7
R1142 GND.n669 GND.n668 74752.4
R1143 GND.n1581 GND.t875 54281.4
R1144 GND.n1583 GND.n194 53707.2
R1145 GND.n1316 GND.n369 52236.1
R1146 GND.n1505 GND.n239 40814.8
R1147 GND.n1354 GND.n240 39303.2
R1148 GND.n1358 GND.n237 37209.3
R1149 GND.n194 GND.n193 35921.1
R1150 GND.n1564 GND.n199 32324.4
R1151 GND.n1517 GND.n200 32324.4
R1152 GND.n1517 GND.n199 32321.1
R1153 GND.n1564 GND.n200 32321.1
R1154 GND.n669 GND.n231 31697.7
R1155 GND.n1506 GND.n236 30691.4
R1156 GND.n335 GND.n334 28676.6
R1157 GND.n1331 GND.n335 28676.6
R1158 GND.n1393 GND.n334 28673.3
R1159 GND.n1393 GND.n1331 28673.3
R1160 GND.n1390 GND.n1332 27409.3
R1161 GND.n1390 GND.n1333 27409.3
R1162 GND.n1369 GND.n1332 27406
R1163 GND.n1369 GND.n1333 27406
R1164 GND.n1216 GND.t844 19674.4
R1165 GND.n1867 GND.n7 19095.8
R1166 GND.n1361 GND.n1360 19032.4
R1167 GND.t384 GND.t339 16471.1
R1168 GND.t719 GND.t579 15956
R1169 GND.t678 GND.t719 15956
R1170 GND.t844 GND.t678 15956
R1171 GND.t723 GND.t960 15812.5
R1172 GND.n1868 GND.n5 15808.4
R1173 GND.n1868 GND.n6 15808.4
R1174 GND.n1835 GND.n5 15805.2
R1175 GND.n1835 GND.n6 15805.2
R1176 GND.n665 GND.t58 15691
R1177 GND.n1090 GND.n416 15303.1
R1178 GND.n1216 GND.t723 15099.2
R1179 GND.t539 GND.n1848 14676.3
R1180 GND.n1355 GND.n239 14517.6
R1181 GND.n1505 GND.n238 14097.4
R1182 GND.t579 GND.t696 13619
R1183 GND.n1568 GND.n195 13432.1
R1184 GND.n1576 GND.n195 13432.1
R1185 GND.n1568 GND.n196 13432.1
R1186 GND.n1576 GND.n196 13432.1
R1187 GND.n1860 GND.n17 13405
R1188 GND.n1860 GND.n1859 13405
R1189 GND.t223 GND.t540 13246.6
R1190 GND.n1182 GND.n1147 12669.3
R1191 GND.n1853 GND.n1851 12564.6
R1192 GND.n1851 GND.n29 12564.6
R1193 GND.n1849 GND.t539 11803.2
R1194 GND.t3 GND.t735 11314.3
R1195 GND.t668 GND.t592 11314.3
R1196 GND.t491 GND.t644 11314.3
R1197 GND.t460 GND.t517 11314.3
R1198 GND.t420 GND.t488 11314.3
R1199 GND.n324 GND.n240 11217.1
R1200 GND.n1716 GND.n1715 11046.2
R1201 GND.n1716 GND.n18 11046.2
R1202 GND.n1673 GND.n181 11046.2
R1203 GND.n1673 GND.n23 11046.2
R1204 GND.n1601 GND.n1600 11046.2
R1205 GND.n1600 GND.n24 11046.2
R1206 GND.n1504 GND.n231 10105.7
R1207 GND.n1506 GND.n1505 10065.1
R1208 GND.n1550 GND.n213 10050.6
R1209 GND.n1548 GND.n213 10050.6
R1210 GND.n1316 GND.n1315 9941.15
R1211 GND.t122 GND.t140 9900
R1212 GND.n1363 GND.n1354 9777.78
R1213 GND.n1550 GND.n214 9474.26
R1214 GND.n1548 GND.n215 9474.26
R1215 GND.n1362 GND.n1353 9451.85
R1216 GND.n1356 GND.n7 9253.97
R1217 GND.n1363 GND.n1362 9201.59
R1218 GND.n1356 GND.n1353 8875.66
R1219 GND.n260 GND.n231 8850.66
R1220 GND.n1848 GND.n8 8814.47
R1221 GND.t496 GND.t457 8567.4
R1222 GND.n1514 GND.n233 8548.9
R1223 GND.n1514 GND.n1511 8548.9
R1224 GND.n1558 GND.n205 8548.9
R1225 GND.n1558 GND.n1557 8548.9
R1226 GND.n254 GND.n241 8242.76
R1227 GND.n1216 GND.n384 8095.54
R1228 GND.n233 GND.n220 7972.6
R1229 GND.n1539 GND.n220 7972.6
R1230 GND.n1539 GND.n226 7972.6
R1231 GND.n226 GND.n205 7972.6
R1232 GND.n1511 GND.n219 7972.6
R1233 GND.n1540 GND.n219 7972.6
R1234 GND.n1540 GND.n206 7972.6
R1235 GND.n1557 GND.n206 7972.6
R1236 GND.t960 GND.t490 7871.88
R1237 GND.n1317 GND.t554 7700
R1238 GND.n434 GND.n426 7416.07
R1239 GND.n430 GND.n426 7416.07
R1240 GND.n434 GND.n429 7416.07
R1241 GND.n430 GND.n429 7416.07
R1242 GND.n1194 GND.n411 7376.47
R1243 GND.n1170 GND.n1168 7376.47
R1244 GND.n1215 GND.t888 7333.33
R1245 GND.n1407 GND.n317 7323.68
R1246 GND.n1565 GND.n193 7195.46
R1247 GND.n1850 GND.n1849 6629.1
R1248 GND.n1124 GND.n1123 6513.16
R1249 GND.n1182 GND.n1181 6156.3
R1250 GND.t394 GND.n665 6141.67
R1251 GND.n1196 GND.n400 6036.13
R1252 GND.n1820 GND.n151 5956.02
R1253 GND.n1807 GND.n151 5956.02
R1254 GND.n671 GND.n670 5949.49
R1255 GND.n8 GND.t384 5876.32
R1256 GND.n1584 GND.n1583 5498.19
R1257 GND.t816 GND.t911 5438.89
R1258 GND.t911 GND.t564 5438.89
R1259 GND.t564 GND.t912 5438.89
R1260 GND.t398 GND.t912 5438.89
R1261 GND.t398 GND.t400 5438.89
R1262 GND.t913 GND.t576 5438.89
R1263 GND.t399 GND.t913 5438.89
R1264 GND.t395 GND.t399 5438.89
R1265 GND.t835 GND.t395 5438.89
R1266 GND.t394 GND.t835 5438.89
R1267 GND.n1361 GND.n1355 5191.76
R1268 GND.n670 GND.n669 5155.69
R1269 GND.n1463 GND.n278 5016.93
R1270 GND.n1367 GND.n7 5009.74
R1271 GND.n1503 GND.n240 4999.47
R1272 GND.n1103 GND.n295 4924.62
R1273 GND.n1443 GND.n295 4924.62
R1274 GND.n1360 GND.n1356 4726.5
R1275 GND.n159 GND.n152 4724.07
R1276 GND.n1810 GND.n159 4724.07
R1277 GND.n1030 GND.n1029 4714.29
R1278 GND.n1011 GND.n888 4714.29
R1279 GND.n1002 GND.n1001 4714.29
R1280 GND.n983 GND.n920 4714.29
R1281 GND.n974 GND.n973 4714.29
R1282 GND.t58 GND.t3 4641.76
R1283 GND.t735 GND.t668 4641.76
R1284 GND.t592 GND.t491 4641.76
R1285 GND.t644 GND.t460 4641.76
R1286 GND.t517 GND.t420 4641.76
R1287 GND.t488 GND.t888 4641.76
R1288 GND.t696 GND.t755 4641.76
R1289 GND.n1555 GND.n208 4597.17
R1290 GND.n1555 GND.n209 4597.17
R1291 GND.n1866 GND.n8 4580.42
R1292 GND.n696 GND.n611 4533.07
R1293 GND.n696 GND.n612 4533.07
R1294 GND.n1476 GND.n267 4458.86
R1295 GND.n268 GND.n267 4458.86
R1296 GND.n268 GND.n266 4458.86
R1297 GND.n1476 GND.n266 4458.86
R1298 GND.n1421 GND.n301 4458.86
R1299 GND.n1421 GND.n302 4458.86
R1300 GND.n1086 GND.n302 4458.86
R1301 GND.n1086 GND.n301 4458.86
R1302 GND.n1147 GND.n417 4458.86
R1303 GND.n1104 GND.n417 4458.86
R1304 GND.n1104 GND.n418 4458.86
R1305 GND.n1147 GND.n418 4458.86
R1306 GND.n1501 GND.n243 4458.86
R1307 GND.n1501 GND.n244 4458.86
R1308 GND.n244 GND.n242 4458.86
R1309 GND.n243 GND.n242 4458.86
R1310 GND.n1491 GND.n252 4458.86
R1311 GND.n1491 GND.n253 4458.86
R1312 GND.n1493 GND.n253 4458.86
R1313 GND.n1493 GND.n252 4458.86
R1314 GND.n1483 GND.n259 4458.86
R1315 GND.n1485 GND.n259 4458.86
R1316 GND.n1485 GND.n258 4458.86
R1317 GND.n1483 GND.n258 4458.86
R1318 GND.n328 GND.n323 4458.86
R1319 GND.n330 GND.n323 4458.86
R1320 GND.n330 GND.n322 4458.86
R1321 GND.n328 GND.n322 4458.86
R1322 GND.n1404 GND.n315 4458.86
R1323 GND.n1404 GND.n316 4458.86
R1324 GND.n1408 GND.n316 4458.86
R1325 GND.n1408 GND.n315 4458.86
R1326 GND.n1414 GND.n309 4458.86
R1327 GND.n1416 GND.n309 4458.86
R1328 GND.n1416 GND.n308 4458.86
R1329 GND.n1414 GND.n308 4458.86
R1330 GND.n1139 GND.n1121 4458.86
R1331 GND.n1139 GND.n1125 4458.86
R1332 GND.n1141 GND.n1121 4458.86
R1333 GND.n1141 GND.n1125 4458.86
R1334 GND.n1366 GND.n1353 4451.25
R1335 GND.n1774 GND.n162 4431.2
R1336 GND.n1774 GND.n163 4431.2
R1337 GND.n1712 GND.n1604 4431.2
R1338 GND.n1712 GND.n1603 4431.2
R1339 GND.n1362 GND.n1361 4206.29
R1340 GND.n1598 GND.n185 4099.91
R1341 GND.n214 GND.n209 4020.88
R1342 GND.n215 GND.n208 4020.88
R1343 GND.n1109 GND.n277 3998.27
R1344 GND.t755 GND.n1215 3980.95
R1345 GND.n1466 GND.n277 3956.88
R1346 GND.n1433 GND.n300 3883.67
R1347 GND.n1357 GND.n190 3871.62
R1348 GND.n1425 GND.n300 3842.28
R1349 GND.n1505 GND.n1504 3789.17
R1350 GND.n1364 GND.n1363 3752.03
R1351 GND.n1359 GND.n190 3679.31
R1352 GND.n1590 GND.n185 3661.93
R1353 GND.n1114 GND.n1112 3641.73
R1354 GND.n1820 GND.n150 3513.17
R1355 GND.n1807 GND.n1776 3513.17
R1356 GND.n1354 GND.n239 3386.33
R1357 GND.t140 GND.t832 3300
R1358 GND.n1215 GND.n392 3253.78
R1359 GND.n672 GND.n456 3250.5
R1360 GND.n854 GND.n456 3250.5
R1361 GND.n854 GND.n457 3250.5
R1362 GND.n850 GND.n457 3250.5
R1363 GND.n850 GND.n461 3250.5
R1364 GND.n846 GND.n461 3250.5
R1365 GND.n846 GND.n473 3250.5
R1366 GND.n841 GND.n473 3250.5
R1367 GND.n841 GND.n480 3250.5
R1368 GND.t400 GND.n697 3193.06
R1369 GND.n1360 GND.n1359 3175.99
R1370 GND.n1357 GND.n193 3165.9
R1371 GND.n860 GND.n451 3151.5
R1372 GND.n458 GND.n451 3151.5
R1373 GND.n459 GND.n458 3151.5
R1374 GND.n460 GND.n459 3151.5
R1375 GND.n476 GND.n460 3151.5
R1376 GND.n477 GND.n476 3151.5
R1377 GND.n478 GND.n477 3151.5
R1378 GND.n479 GND.n478 3151.5
R1379 GND.n485 GND.n479 3151.5
R1380 GND.n1368 GND.n8 3148.07
R1381 GND.n1598 GND.n184 3111.98
R1382 GND.t457 GND.t87 3062.55
R1383 GND.t456 GND.t496 3062.55
R1384 GND.n1425 GND.n287 3036.9
R1385 GND.n1736 GND.n1731 2982.78
R1386 GND.n1737 GND.n1736 2982.78
R1387 GND.n1737 GND.n1732 2982.78
R1388 GND.n1732 GND.n1731 2982.78
R1389 GND.t832 GND.t794 2887.5
R1390 GND.t794 GND.t554 2887.5
R1391 GND.n22 GND.n8 2813.2
R1392 GND.n436 GND.n286 2801.33
R1393 GND.n1590 GND.n1589 2772.79
R1394 GND.n1611 GND.n1604 2750.4
R1395 GND.n1611 GND.n1610 2750.4
R1396 GND.n1610 GND.n12 2750.4
R1397 GND.n1757 GND.n12 2750.4
R1398 GND.n1757 GND.n1751 2750.4
R1399 GND.n1768 GND.n1751 2750.4
R1400 GND.n1768 GND.n1752 2750.4
R1401 GND.n1752 GND.n163 2750.4
R1402 GND.n1609 GND.n1603 2750.4
R1403 GND.n1609 GND.n1608 2750.4
R1404 GND.n1608 GND.n11 2750.4
R1405 GND.n1761 GND.n11 2750.4
R1406 GND.n1761 GND.n1753 2750.4
R1407 GND.n1766 GND.n1753 2750.4
R1408 GND.n1766 GND.n1755 2750.4
R1409 GND.n1755 GND.n162 2750.4
R1410 GND.t267 GND.t30 2721.05
R1411 GND.t30 GND.t32 2721.05
R1412 GND.t32 GND.t432 2721.05
R1413 GND.t432 GND.t452 2721.05
R1414 GND.t452 GND.t584 2721.05
R1415 GND.t584 GND.t429 2721.05
R1416 GND.t34 GND.t436 2721.05
R1417 GND.t471 GND.t34 2721.05
R1418 GND.t473 GND.t471 2721.05
R1419 GND.t446 GND.t473 2721.05
R1420 GND.t67 GND.t446 2721.05
R1421 GND.t468 GND.t67 2721.05
R1422 GND.t438 GND.t468 2721.05
R1423 GND.t63 GND.t438 2721.05
R1424 GND.t332 GND.t63 2721.05
R1425 GND.t273 GND.t332 2721.05
R1426 GND.n670 GND.n578 2710.35
R1427 GND.t877 GND.n1578 2601.35
R1428 GND.n1583 GND.n1582 2554.93
R1429 GND.n1818 GND.n135 2533.93
R1430 GND.n1818 GND.n136 2533.93
R1431 GND.n1831 GND.n136 2533.93
R1432 GND.n1831 GND.n135 2533.93
R1433 GND.n1589 GND.n1588 2517.57
R1434 GND.n1584 GND.n193 2511.21
R1435 GND.n1435 GND.n294 2463.9
R1436 GND.n1812 GND.n1811 2384.32
R1437 GND.n1812 GND.n153 2384.32
R1438 GND.n1473 GND.n269 2381.13
R1439 GND.n1319 GND.n1318 2374.87
R1440 GND.n1811 GND.n156 2339.75
R1441 GND.n1776 GND.n156 2339.75
R1442 GND.n153 GND.n152 2339.75
R1443 GND.n1816 GND.n153 2339.75
R1444 GND.n1816 GND.n150 2339.75
R1445 GND.n1811 GND.n1810 2339.75
R1446 GND.n21 GND.n18 2317.47
R1447 GND.n23 GND.n21 2317.47
R1448 GND.n1715 GND.n1714 2317.47
R1449 GND.n1714 GND.n181 2317.47
R1450 GND.n1715 GND.n17 2276.08
R1451 GND.n1859 GND.n18 2276.08
R1452 GND.n1585 GND.n1584 2269.61
R1453 GND.n1463 GND.n279 2266.53
R1454 GND.n1852 GND.n22 2221.71
R1455 GND.t392 GND.t55 2200
R1456 GND.t422 GND.t666 2200
R1457 GND.t667 GND.t757 2200
R1458 GND.t757 GND.t415 2200
R1459 GND.n1866 GND.t436 2185.53
R1460 GND.n1473 GND.n270 2101
R1461 GND.n1446 GND.n293 2040.52
R1462 GND.n29 GND.t267 2024.68
R1463 GND.t635 GND.t766 1997.37
R1464 GND.t766 GND.t769 1997.37
R1465 GND.t637 GND.t634 1997.37
R1466 GND.t680 GND.t637 1997.37
R1467 GND.t770 GND.t680 1997.37
R1468 GND.t612 GND.t602 1997.37
R1469 GND.t602 GND.t607 1997.37
R1470 GND.t607 GND.t611 1997.37
R1471 GND.t598 GND.t603 1997.37
R1472 GND.t603 GND.t604 1997.37
R1473 GND.t604 GND.t605 1997.37
R1474 GND.t749 GND.t570 1997.37
R1475 GND.t871 GND.t749 1997.37
R1476 GND.t828 GND.t871 1997.37
R1477 GND.t747 GND.t750 1997.37
R1478 GND.t750 GND.t748 1997.37
R1479 GND.t748 GND.t745 1997.37
R1480 GND.t55 GND.t422 1997.37
R1481 GND.t666 GND.t667 1997.37
R1482 GND.t153 GND.t465 1997.37
R1483 GND.t154 GND.t153 1997.37
R1484 GND.t464 GND.t154 1997.37
R1485 GND.t643 GND.t495 1997.37
R1486 GND.t495 GND.t463 1997.37
R1487 GND.t463 GND.t642 1997.37
R1488 GND.t528 GND.t530 1997.37
R1489 GND.t530 GND.t599 1997.37
R1490 GND.t599 GND.t527 1997.37
R1491 GND.t601 GND.t606 1997.37
R1492 GND.t606 GND.t610 1997.37
R1493 GND.t610 GND.t600 1997.37
R1494 GND.t812 GND.t486 1997.37
R1495 GND.t486 GND.t366 1997.37
R1496 GND.t366 GND.t811 1997.37
R1497 GND.t131 GND.t485 1997.37
R1498 GND.t44 GND.t131 1997.37
R1499 GND.t711 GND.t44 1997.37
R1500 GND.n1852 GND.t273 1982.89
R1501 GND.n1466 GND.n270 1951.38
R1502 GND.t877 GND.n1579 1917.57
R1503 GND.t875 GND.n1579 1917.57
R1504 GND.n1869 GND.n4 1874.45
R1505 GND.n1869 GND.n3 1874.45
R1506 GND.n1836 GND.n3 1874.07
R1507 GND.n1405 GND.n240 1773.03
R1508 GND.n1867 GND.t223 1763.49
R1509 GND.n1359 GND.n1358 1739.72
R1510 GND.n133 GND.n4 1734.78
R1511 GND.t745 GND.n323 1687.7
R1512 GND.n244 GND.t711 1687.7
R1513 GND.n1594 GND.n189 1686.07
R1514 GND.n1614 GND.n1609 1680.8
R1515 GND.n1614 GND.n1611 1680.8
R1516 GND.n1864 GND.n11 1680.8
R1517 GND.n1864 GND.n12 1680.8
R1518 GND.n1758 GND.n1753 1680.8
R1519 GND.n1758 GND.n1751 1680.8
R1520 GND.n1755 GND.n1754 1680.8
R1521 GND.n1754 GND.n1752 1680.8
R1522 GND.n1433 GND.n293 1664.88
R1523 GND.t885 GND.n384 1608.12
R1524 GND.n1358 GND.n1357 1603.26
R1525 GND.n1269 GND.t721 1576.25
R1526 GND.t368 GND.t57 1548.86
R1527 GND.n317 GND.t770 1541.45
R1528 GND.n1407 GND.t612 1541.45
R1529 GND.t605 GND.n1405 1541.45
R1530 GND.t570 GND.n324 1541.45
R1531 GND.t415 GND.n236 1541.45
R1532 GND.t465 GND.n260 1541.45
R1533 GND.t642 GND.n238 1541.45
R1534 GND.n1124 GND.t636 1541.45
R1535 GND.n1123 GND.t528 1541.45
R1536 GND.t600 GND.n254 1541.45
R1537 GND.n1847 GND.n28 1485.93
R1538 GND.n1847 GND.n30 1485.93
R1539 GND.n1602 GND.n181 1477.07
R1540 GND.n1602 GND.n1601 1477.07
R1541 GND.n1857 GND.n23 1477.07
R1542 GND.n1857 GND.n24 1477.07
R1543 GND.n294 GND.n279 1464.33
R1544 GND.n1215 GND.n1214 1460.5
R1545 GND.n1109 GND.n269 1438.87
R1546 GND.n1853 GND.n24 1435.68
R1547 GND.n1601 GND.n29 1435.68
R1548 GND.n1587 GND.n184 1373.22
R1549 GND.t88 GND.t56 1346.78
R1550 GND.n1503 GND.t812 1346.05
R1551 GND.n1318 GND.n1317 1339.85
R1552 GND.n1717 GND.n178 1306.35
R1553 GND.n1717 GND.n180 1306.35
R1554 GND.n1700 GND.n1699 1306.35
R1555 GND.n1699 GND.n25 1306.35
R1556 GND.n1702 GND.n27 1306.35
R1557 GND.n1855 GND.n27 1306.35
R1558 GND.n428 GND.t390 1302.63
R1559 GND.t9 GND.t5 1261.42
R1560 GND.n390 GND.n377 1255.62
R1561 GND.n1355 GND.n237 1240.24
R1562 GND.n1588 GND.n1585 1222.22
R1563 GND.n1183 GND.n1182 1220.17
R1564 GND.n1038 GND.n1037 1219.11
R1565 GND.n391 GND.n380 1198.25
R1566 GND.n1283 GND.n381 1198.25
R1567 GND.n386 GND.n373 1198.25
R1568 GND.n1270 GND.n1269 1198.25
R1569 GND.n1268 GND.n1267 1198.25
R1570 GND.n1257 GND.n1256 1198.25
R1571 GND.n1255 GND.n1254 1198.25
R1572 GND.n515 GND.n501 1198.25
R1573 GND.n367 GND.n366 1198.25
R1574 GND.n726 GND.n578 1198.25
R1575 GND.n737 GND.n575 1198.25
R1576 GND.n748 GND.n571 1198.25
R1577 GND.n759 GND.n567 1198.25
R1578 GND.n770 GND.n563 1198.25
R1579 GND.n781 GND.n559 1198.25
R1580 GND.n792 GND.n555 1198.25
R1581 GND.n803 GND.n551 1198.25
R1582 GND.n814 GND.n547 1198.25
R1583 GND.n825 GND.n543 1198.25
R1584 GND.n1320 GND.n1319 1198.25
R1585 GND.n1243 GND.n1240 1198.01
R1586 GND.t0 GND.t88 1185.54
R1587 GND.n668 GND 1178.42
R1588 GND GND.n698 1177.5
R1589 GND.n609 GND 1177.5
R1590 GND GND.n620 1177.5
R1591 GND.n663 GND 1177.5
R1592 GND GND.n680 1177.5
R1593 GND.n1551 GND.n212 1153.51
R1594 GND.t5 GND.n240 1142.5
R1595 GND.t54 GND.n1364 1134.47
R1596 GND.t387 GND.n1366 1108.21
R1597 GND GND.t954 1104.21
R1598 GND.t19 GND.t548 1102.37
R1599 GND.t41 GND.n1367 1095.81
R1600 GND.n1552 GND.n1551 1083.11
R1601 GND.n1547 GND.n216 1083.11
R1602 GND.t504 GND.n678 1034.5
R1603 GND.n1504 GND.n1503 1020.1
R1604 GND.n1330 GND.t364 1011.91
R1605 GND.n183 GND.t456 1007.93
R1606 GND.n1415 GND.t769 998.684
R1607 GND.n1415 GND.t634 998.684
R1608 GND.t611 GND.n1406 998.684
R1609 GND.n1406 GND.t598 998.684
R1610 GND.n329 GND.t828 998.684
R1611 GND.n329 GND.t747 998.684
R1612 GND.n1484 GND.t464 998.684
R1613 GND.n1484 GND.t643 998.684
R1614 GND.n1492 GND.t527 998.684
R1615 GND.n1492 GND.t601 998.684
R1616 GND.t811 GND.n1502 998.684
R1617 GND.n1502 GND.t485 998.684
R1618 GND.n1480 GND.n1479 982.966
R1619 GND.n1513 GND.n1512 981.836
R1620 GND.n1392 GND.t368 938.22
R1621 GND.t405 GND.t559 938.072
R1622 GND.n679 GND.t504 935.114
R1623 GND.n1785 GND.n1776 922.962
R1624 GND.n1785 GND.n150 922.962
R1625 GND.n1512 GND.n218 911.436
R1626 GND.n1541 GND.n218 911.436
R1627 GND.n1542 GND.n1541 911.436
R1628 GND.n1435 GND.n293 904.067
R1629 GND.n1446 GND.n287 900.884
R1630 GND.t832 GND.t955 893.402
R1631 GND.t794 GND.t142 893.402
R1632 GND.n1039 GND.n1038 890.795
R1633 GND.t217 GND.n22 889.937
R1634 GND.n1589 GND.n189 889.139
R1635 GND.n1037 GND.n867 887.395
R1636 GND.n1031 GND.n867 887.395
R1637 GND.n1031 GND.n1030 887.395
R1638 GND.n1029 GND.n877 887.395
R1639 GND.n1023 GND.n877 887.395
R1640 GND.n1023 GND.n1022 887.395
R1641 GND.n1022 GND.n1021 887.395
R1642 GND.n1021 GND.n888 887.395
R1643 GND.n1011 GND.n1010 887.395
R1644 GND.n1010 GND.n1009 887.395
R1645 GND.n1009 GND.n899 887.395
R1646 GND.n1003 GND.n899 887.395
R1647 GND.n1003 GND.n1002 887.395
R1648 GND.n1001 GND.n909 887.395
R1649 GND.n995 GND.n909 887.395
R1650 GND.n995 GND.n994 887.395
R1651 GND.n994 GND.n993 887.395
R1652 GND.n993 GND.n920 887.395
R1653 GND.n983 GND.n982 887.395
R1654 GND.n982 GND.n981 887.395
R1655 GND.n981 GND.n931 887.395
R1656 GND.n975 GND.n931 887.395
R1657 GND.n975 GND.n974 887.395
R1658 GND.n973 GND.n941 887.395
R1659 GND.n967 GND.n941 887.395
R1660 GND.n967 GND.n966 887.395
R1661 GND.n966 GND.n965 887.395
R1662 GND.n965 GND.n392 887.395
R1663 GND.n1214 GND.n393 887.395
R1664 GND.n1208 GND.n393 887.395
R1665 GND.n1208 GND.n1207 887.395
R1666 GND.n1207 GND.n1206 887.395
R1667 GND.n1206 GND.n400 887.395
R1668 GND.n1196 GND.n1195 887.395
R1669 GND.n1195 GND.n1194 887.395
R1670 GND.n1184 GND.n411 887.395
R1671 GND.n1184 GND.n1183 887.395
R1672 GND.n1181 GND.n1148 887.395
R1673 GND.n1168 GND.n1148 887.395
R1674 GND.n1170 GND.n1169 887.395
R1675 GND.n1169 GND.n369 887.395
R1676 GND.t960 GND 859.899
R1677 GND.n432 GND.n431 852.33
R1678 GND.n433 GND.n432 852.33
R1679 GND GND.n386 848.731
R1680 GND.t721 GND 842.913
R1681 GND.n1114 GND.n436 840.4
R1682 GND GND.n391 837.563
R1683 GND.n1577 GND.t79 835.664
R1684 GND.n698 GND.n609 827.04
R1685 GND.n663 GND.n620 827.04
R1686 GND.n1315 GND 826.396
R1687 GND.t390 GND.n231 817.764
R1688 GND.n1713 GND.n1599 799.255
R1689 GND.t365 GND.n1566 790.207
R1690 GND.t18 GND.n1365 786.471
R1691 GND.n427 GND.n264 781.929
R1692 GND.n427 GND.n261 781.929
R1693 GND GND.t173 781.726
R1694 GND.t821 GND 781.726
R1695 GND.n1585 GND.t498 778.601
R1696 GND.t795 GND.t839 775.48
R1697 GND.n1059 GND.n1047 769.572
R1698 GND.n1068 GND.n1049 769.572
R1699 GND.n1077 GND.n1051 769.572
R1700 GND.n1084 GND.n1083 769.572
R1701 GND.n680 GND.n679 765.375
R1702 GND.n1391 GND.t56 758.747
R1703 GND.n1547 GND.n1546 739.765
R1704 GND.n1834 GND.n1833 735.025
R1705 GND.t498 GND.n192 715.226
R1706 GND.n192 GND.t454 715.226
R1707 GND.t670 GND 714.721
R1708 GND.t122 GND 714.721
R1709 GND GND.t554 714.721
R1710 GND.n1821 GND.n149 709.271
R1711 GND.n1806 GND.n149 709.271
R1712 GND.n1269 GND.n1217 708.047
R1713 GND.t764 GND.t410 708.047
R1714 GND.t120 GND.t406 708.047
R1715 GND.t829 GND.t141 708.047
R1716 GND.n1318 GND.n368 708.047
R1717 GND.t862 GND.t10 708.047
R1718 GND.t10 GND.t122 708.047
R1719 GND.n1567 GND.t365 701.784
R1720 GND.n665 GND.t797 700.206
R1721 GND.n428 GND.t392 694.737
R1722 GND.n1582 GND.n1577 684.348
R1723 GND.t937 GND 681.218
R1724 GND.n1559 GND.n204 675.013
R1725 GND.n1402 GND.n319 669.365
R1726 GND.n1566 GND.t79 656.327
R1727 GND.n1808 GND.n1775 655.385
R1728 GND.n389 GND.n388 649.043
R1729 GND.n318 GND.n246 646.4
R1730 GND.n678 GND.n671 634.702
R1731 GND.n1368 GND.t41 623.778
R1732 GND GND.n368 623.755
R1733 GND.t140 GND 603.047
R1734 GND.n218 GND.n216 601.977
R1735 GND.n1546 GND.n1542 601.977
R1736 GND.n1545 GND.n1544 601.977
R1737 GND.n1315 GND.n1314 599.125
R1738 GND.n1239 GND.n368 599.125
R1739 GND.n1274 GND.n384 599.125
R1740 GND.n1462 GND.n280 592.888
R1741 GND.n1216 GND.t147 590.955
R1742 GND.t413 GND.n389 590.039
R1743 GND.t126 GND 590.038
R1744 GND GND.t867 590.038
R1745 GND GND.t552 590.038
R1746 GND.n1076 GND.n1075 585
R1747 GND.n1074 GND.n1050 585
R1748 GND.n1091 GND.n1050 585
R1749 GND.n1067 GND.n1066 585
R1750 GND.n1065 GND.n1048 585
R1751 GND.n1091 GND.n1048 585
R1752 GND.n1058 GND.n1057 585
R1753 GND.n1056 GND.n1046 585
R1754 GND.n1091 GND.n1046 585
R1755 GND.n1093 GND.n1092 585
R1756 GND.n1092 GND.n1091 585
R1757 GND.n1044 GND.n1043 585
R1758 GND.n1166 GND.n1165 585
R1759 GND.n1166 GND.n369 585
R1760 GND.n1167 GND.n1160 585
R1761 GND.n1169 GND.n1167 585
R1762 GND.n1172 GND.n1171 585
R1763 GND.n1171 GND.n1170 585
R1764 GND.n1177 GND.n1157 585
R1765 GND.n1168 GND.n1157 585
R1766 GND.n1178 GND.n1149 585
R1767 GND.n1149 GND.n1148 585
R1768 GND.n1180 GND.n1179 585
R1769 GND.n1181 GND.n1180 585
R1770 GND.n1150 GND.n415 585
R1771 GND.n1183 GND.n415 585
R1772 GND.n1185 GND.n414 585
R1773 GND.n1185 GND.n1184 585
R1774 GND.n1187 GND.n1186 585
R1775 GND.n1186 GND.n411 585
R1776 GND.n1193 GND.n1192 585
R1777 GND.n1194 GND.n1193 585
R1778 GND.n410 GND.n409 585
R1779 GND.n1195 GND.n410 585
R1780 GND.n1198 GND.n1197 585
R1781 GND.n1197 GND.n1196 585
R1782 GND.n1203 GND.n401 585
R1783 GND.n401 GND.n400 585
R1784 GND.n1205 GND.n1204 585
R1785 GND.n1206 GND.n1205 585
R1786 GND.n399 GND.n398 585
R1787 GND.n1207 GND.n399 585
R1788 GND.n1210 GND.n1209 585
R1789 GND.n1209 GND.n1208 585
R1790 GND.n1211 GND.n394 585
R1791 GND.n394 GND.n393 585
R1792 GND.n1213 GND.n1212 585
R1793 GND.n1214 GND.n1213 585
R1794 GND.n962 GND.n952 585
R1795 GND.n952 GND.n392 585
R1796 GND.n964 GND.n963 585
R1797 GND.n965 GND.n964 585
R1798 GND.n951 GND.n950 585
R1799 GND.n966 GND.n951 585
R1800 GND.n969 GND.n968 585
R1801 GND.n968 GND.n967 585
R1802 GND.n970 GND.n942 585
R1803 GND.n942 GND.n941 585
R1804 GND.n972 GND.n971 585
R1805 GND.n973 GND.n972 585
R1806 GND.n940 GND.n939 585
R1807 GND.n974 GND.n940 585
R1808 GND.n977 GND.n976 585
R1809 GND.n976 GND.n975 585
R1810 GND.n978 GND.n932 585
R1811 GND.n932 GND.n931 585
R1812 GND.n980 GND.n979 585
R1813 GND.n981 GND.n980 585
R1814 GND.n930 GND.n929 585
R1815 GND.n982 GND.n930 585
R1816 GND.n985 GND.n984 585
R1817 GND.n984 GND.n983 585
R1818 GND.n990 GND.n921 585
R1819 GND.n921 GND.n920 585
R1820 GND.n992 GND.n991 585
R1821 GND.n993 GND.n992 585
R1822 GND.n919 GND.n918 585
R1823 GND.n994 GND.n919 585
R1824 GND.n997 GND.n996 585
R1825 GND.n996 GND.n995 585
R1826 GND.n998 GND.n910 585
R1827 GND.n910 GND.n909 585
R1828 GND.n1000 GND.n999 585
R1829 GND.n1001 GND.n1000 585
R1830 GND.n908 GND.n907 585
R1831 GND.n1002 GND.n908 585
R1832 GND.n1005 GND.n1004 585
R1833 GND.n1004 GND.n1003 585
R1834 GND.n1006 GND.n900 585
R1835 GND.n900 GND.n899 585
R1836 GND.n1008 GND.n1007 585
R1837 GND.n1009 GND.n1008 585
R1838 GND.n898 GND.n897 585
R1839 GND.n1010 GND.n898 585
R1840 GND.n1013 GND.n1012 585
R1841 GND.n1012 GND.n1011 585
R1842 GND.n1018 GND.n889 585
R1843 GND.n889 GND.n888 585
R1844 GND.n1020 GND.n1019 585
R1845 GND.n1021 GND.n1020 585
R1846 GND.n887 GND.n886 585
R1847 GND.n1022 GND.n887 585
R1848 GND.n1025 GND.n1024 585
R1849 GND.n1024 GND.n1023 585
R1850 GND.n1026 GND.n878 585
R1851 GND.n878 GND.n877 585
R1852 GND.n1028 GND.n1027 585
R1853 GND.n1029 GND.n1028 585
R1854 GND.n876 GND.n875 585
R1855 GND.n1030 GND.n876 585
R1856 GND.n1033 GND.n1032 585
R1857 GND.n1032 GND.n1031 585
R1858 GND.n1034 GND.n868 585
R1859 GND.n868 GND.n867 585
R1860 GND.n1036 GND.n1035 585
R1861 GND.n1037 GND.n1036 585
R1862 GND.n866 GND.n865 585
R1863 GND.n1127 GND 583.907
R1864 GND.n1441 GND.n297 582.4
R1865 GND.n222 GND.n215 576.293
R1866 GND.n222 GND.n214 576.293
R1867 GND.n1509 GND.n220 576.293
R1868 GND.n1509 GND.n219 576.293
R1869 GND.n226 GND.n225 576.293
R1870 GND.n225 GND.n206 576.293
R1871 GND.n1544 GND.n207 568.095
R1872 GND.n1518 GND.n230 566.203
R1873 GND.t797 GND.n450 562.423
R1874 GND.n1560 GND.n1559 542.871
R1875 GND GND.t650 539.465
R1876 GND GND.t873 539.465
R1877 GND.n1036 GND.n866 539.294
R1878 GND.n1036 GND.n868 539.294
R1879 GND.n1032 GND.n868 539.294
R1880 GND.n1032 GND.n876 539.294
R1881 GND.n1028 GND.n878 539.294
R1882 GND.n1024 GND.n878 539.294
R1883 GND.n1024 GND.n887 539.294
R1884 GND.n1020 GND.n887 539.294
R1885 GND.n1020 GND.n889 539.294
R1886 GND.n1012 GND.n898 539.294
R1887 GND.n1008 GND.n898 539.294
R1888 GND.n1008 GND.n900 539.294
R1889 GND.n1004 GND.n900 539.294
R1890 GND.n1004 GND.n908 539.294
R1891 GND.n1000 GND.n910 539.294
R1892 GND.n996 GND.n910 539.294
R1893 GND.n996 GND.n919 539.294
R1894 GND.n992 GND.n919 539.294
R1895 GND.n992 GND.n921 539.294
R1896 GND.n984 GND.n930 539.294
R1897 GND.n980 GND.n930 539.294
R1898 GND.n980 GND.n932 539.294
R1899 GND.n976 GND.n932 539.294
R1900 GND.n976 GND.n940 539.294
R1901 GND.n972 GND.n942 539.294
R1902 GND.n968 GND.n942 539.294
R1903 GND.n968 GND.n951 539.294
R1904 GND.n964 GND.n951 539.294
R1905 GND.n964 GND.n952 539.294
R1906 GND.n1213 GND.n394 539.294
R1907 GND.n1209 GND.n394 539.294
R1908 GND.n1209 GND.n399 539.294
R1909 GND.n1205 GND.n399 539.294
R1910 GND.n1205 GND.n401 539.294
R1911 GND.n1197 GND.n410 539.294
R1912 GND.n1193 GND.n410 539.294
R1913 GND.n1186 GND.n1185 539.294
R1914 GND.n1185 GND.n415 539.294
R1915 GND.n1180 GND.n1149 539.294
R1916 GND.n1157 GND.n1149 539.294
R1917 GND.n1171 GND.n1167 539.294
R1918 GND.n1167 GND.n1166 539.294
R1919 GND.n1057 GND.n1046 539.294
R1920 GND.n1066 GND.n1048 539.294
R1921 GND.n1075 GND.n1050 539.294
R1922 GND.n1092 GND.n1044 539.294
R1923 GND.n391 GND.t615 536.042
R1924 GND.n386 GND.t405 536.042
R1925 GND.n1866 GND.t429 535.527
R1926 GND.n1554 GND.n1553 530.072
R1927 GND.n1773 GND.n1772 528.942
R1928 GND.n1773 GND.n164 528.942
R1929 GND.n1711 GND.n1605 528.942
R1930 GND.n614 GND.n613 525.178
R1931 GND.n695 GND.n694 525.178
R1932 GND GND.t547 522.606
R1933 GND GND.t172 522.606
R1934 GND.n160 GND.n139 521.788
R1935 GND.n1182 GND.n416 517.648
R1936 GND.n447 GND.n297 516.841
R1937 GND.n1538 GND.n227 514.26
R1938 GND.n327 GND.n321 514.26
R1939 GND.n1085 GND.n304 514.26
R1940 GND.n1482 GND.n256 514.26
R1941 GND.n1477 GND.n265 514.26
R1942 GND.n1146 GND.n419 514.26
R1943 GND.n1500 GND.n1499 514.26
R1944 GND.n1146 GND.n1145 514.26
R1945 GND.n1394 GND.n333 511.591
R1946 GND.n1455 GND.n286 502.967
R1947 GND.n1112 GND.n441 502.967
R1948 GND.t960 GND.t937 502.538
R1949 GND.n1455 GND.n279 499.784
R1950 GND.n441 GND.n278 499.784
R1951 GND.n1111 GND.n269 499.784
R1952 GND.n1118 GND.n270 499.784
R1953 GND.n1112 GND.n1111 496.601
R1954 GND.n1118 GND.n436 496.601
R1955 GND.n1535 GND.n203 496.188
R1956 GND.n232 GND.n229 494.683
R1957 GND.n1575 GND.n197 492.817
R1958 GND.t615 GND.n381 491.372
R1959 GND.n1513 GND.n229 487.154
R1960 GND.n1563 GND.n201 483.003
R1961 GND.t373 GND.t858 480.461
R1962 GND.t723 GND.t885 480.204
R1963 GND.n1537 GND.n1536 475.86
R1964 GND.n1389 GND.n1388 475.536
R1965 GND.t364 GND.n231 473.488
R1966 GND.n1597 GND.n1596 473.224
R1967 GND.n1107 GND.n276 472.848
R1968 GND.n1467 GND.n276 472.848
R1969 GND.n1507 GND.n228 472.471
R1970 GND GND.t27 472.031
R1971 GND.n1103 GND.n278 471.134
R1972 GND.n1443 GND.n294 471.134
R1973 GND.t454 GND.n183 470.783
R1974 GND.t49 GND.t151 470.267
R1975 GND.t910 GND.t144 470.267
R1976 GND.t905 GND.t796 470.267
R1977 GND.t149 GND.t906 470.267
R1978 GND.t150 GND.t47 470.267
R1979 GND.t909 GND.t48 470.267
R1980 GND.t46 GND.t148 470.267
R1981 GND GND.t832 469.036
R1982 GND.n1370 GND.n1352 461.243
R1983 GND.n1575 GND.n1574 461.243
R1984 GND.n1563 GND.n1562 461.243
R1985 GND.n1519 GND.n1518 461.243
R1986 GND.n348 GND.n347 461.243
R1987 GND.n1371 GND.n1370 459.964
R1988 GND.n1850 GND.n8 459.788
R1989 GND.n1553 GND.n1552 459.671
R1990 GND.n1545 GND.n1543 459.671
R1991 GND.n1431 GND.n1427 459.295
R1992 GND.n1427 GND.n1426 459.295
R1993 GND.n349 GND.n348 459.111
R1994 GND.n1389 GND.n1335 458.043
R1995 GND.t723 GND.t670 457.868
R1996 GND.n1569 GND.n198 449.296
R1997 GND.n388 GND.t578 446.745
R1998 GND.t578 GND.n387 446.745
R1999 GND.t173 GND.n381 446.702
R2000 GND.n331 GND.n319 443.86
R2001 GND.n1419 GND.n304 443.86
R2002 GND.n1418 GND.n1417 443.86
R2003 GND.n1417 GND.n306 443.86
R2004 GND.n1401 GND.n313 443.86
R2005 GND.n327 GND.n326 443.86
R2006 GND.n1129 GND.n1128 443.86
R2007 GND.n1128 GND.n1127 443.86
R2008 GND.n1486 GND.n257 443.86
R2009 GND.n1487 GND.n1486 443.86
R2010 GND.n1138 GND.n1137 443.86
R2011 GND.n1490 GND.n1489 443.86
R2012 GND.n1500 GND.n245 443.86
R2013 GND.n1145 GND.n1144 443.86
R2014 GND.n1143 GND.n1142 443.86
R2015 GND.n1142 GND.n425 443.86
R2016 GND.n1494 GND.n251 443.86
R2017 GND.n1495 GND.n1494 443.86
R2018 GND.n1497 GND.n1496 443.86
R2019 GND.n1498 GND.n1497 443.86
R2020 GND GND.t375 442.539
R2021 GND GND.t551 442.539
R2022 GND.t155 GND 442.539
R2023 GND.n232 GND.n228 438.966
R2024 GND.n1560 GND.n203 438.966
R2025 GND.n1240 GND.t124 438.315
R2026 GND.n1217 GND.n1216 436.238
R2027 GND.n1538 GND.n1537 435.577
R2028 GND.n1481 GND.n1480 431.812
R2029 GND.n1115 GND.n437 430.252
R2030 GND.n1496 GND.n1495 428.8
R2031 GND.n1402 GND.n1401 427.671
R2032 GND.n1596 GND.n187 423.154
R2033 GND.n1821 GND.n148 422.582
R2034 GND.n1806 GND.n1778 422.582
R2035 GND.n1536 GND.n1535 415.248
R2036 GND.n1543 GND.n210 415.248
R2037 GND.n1490 GND.n255 414.872
R2038 GND.t858 GND 413.027
R2039 GND.n1488 GND.n245 399.812
R2040 GND.n1775 GND.n161 399.562
R2041 GND GND.n257 399.06
R2042 GND.n1507 GND.n227 397.176
R2043 GND.n1520 GND.n1519 390.416
R2044 GND.n313 GND.n306 380.988
R2045 GND.n1411 GND.n1410 380.988
R2046 GND.n1516 GND.n1515 380.676
R2047 GND.t490 GND.n390 370.882
R2048 GND.n1268 GND.t650 370.882
R2049 GND.n1256 GND.t556 370.882
R2050 GND.t863 GND.n1255 370.882
R2051 GND.n1426 GND.n288 364.048
R2052 GND.t920 GND.t872 363.033
R2053 GND GND.n1569 362.88
R2054 GND.n387 GND.t862 362.454
R2055 GND.n1395 GND.n1394 361.601
R2056 GND.n1597 GND.n186 360.283
R2057 GND.t506 GND.t887 358.81
R2058 GND.n1745 GND.n1730 357.647
R2059 GND.n1745 GND.n1744 357.647
R2060 GND.n1738 GND.n1730 357.647
R2061 GND.n1744 GND.n1738 357.647
R2062 GND.n1820 GND.t232 353.01
R2063 GND.n1144 GND.n420 350.872
R2064 GND.n1143 GND.n423 350.872
R2065 GND.n425 GND.n311 350.872
R2066 GND.n1412 GND.n251 350.872
R2067 GND.n1495 GND.n250 350.872
R2068 GND.n1496 GND.n248 350.872
R2069 GND.n1498 GND.n246 350.872
R2070 GND.n1453 GND.n287 350.168
R2071 GND.n1453 GND.n286 346.983
R2072 GND.n1085 GND.n420 345.976
R2073 GND.n1546 GND.n1545 343.341
R2074 GND.n1544 GND.n1542 343.341
R2075 GND.n1365 GND.t54 342.896
R2076 GND.n1137 GND.n1136 338.825
R2077 GND.n425 GND.n251 338.825
R2078 GND.n390 GND.t413 337.166
R2079 GND.t508 GND.n1268 337.166
R2080 GND.n1256 GND.t126 337.166
R2081 GND.n1255 GND.t867 337.166
R2082 GND GND.t490 335.026
R2083 GND.n1130 GND.n1129 332.8
R2084 GND.n1133 GND.n1127 332.8
R2085 GND.n257 GND.n255 332.8
R2086 GND.n1488 GND.n1487 332.8
R2087 GND.n1116 GND.n285 330.865
R2088 GND.t151 GND.t15 328.938
R2089 GND.t638 GND.t910 328.938
R2090 GND.t144 GND.t896 328.938
R2091 GND.t382 GND.t905 328.938
R2092 GND.t796 GND.t568 328.938
R2093 GND.t691 GND.t149 328.938
R2094 GND.t906 GND.t1 328.938
R2095 GND.t47 GND.t869 328.938
R2096 GND.t773 GND.t150 328.938
R2097 GND.t842 GND.t909 328.938
R2098 GND.t48 GND.t543 328.938
R2099 GND.t943 GND.t46 328.938
R2100 GND.t954 GND.t373 328.736
R2101 GND.n1606 GND.n1605 325.272
R2102 GND.n1607 GND.n1606 325.272
R2103 GND.n1607 GND.n13 325.272
R2104 GND.n1762 GND.n13 325.272
R2105 GND.n1763 GND.n1762 325.272
R2106 GND.n1765 GND.n1763 325.272
R2107 GND.n1765 GND.n1764 325.272
R2108 GND.n1764 GND.n164 325.272
R2109 GND.n191 GND.n187 321.507
R2110 GND.n1419 GND.n1418 317.365
R2111 GND.n310 GND.n303 317.365
R2112 GND.t229 GND.n1808 316.447
R2113 GND.n1131 GND.n1130 313.601
R2114 GND.n583 GND.n230 312.353
R2115 GND.n423 GND.n303 310.589
R2116 GND.n1772 GND.n1771 309.8
R2117 GND.n207 GND.n204 306.825
R2118 GND.t524 GND.t564 304.7
R2119 GND.t835 GND.t17 304.7
R2120 GND.n1830 GND.n137 304.565
R2121 GND.n1817 GND.n137 304.565
R2122 GND.n210 GND 303.06
R2123 GND.n1132 GND.n1131 301.553
R2124 GND.n1144 GND.n1143 301.553
R2125 GND.n1587 GND.n189 299.673
R2126 GND.n585 GND.n584 299.553
R2127 GND GND.n204 298.918
R2128 GND.t825 GND 296.161
R2129 GND.n332 GND.n331 295.906
R2130 GND GND.t508 295.019
R2131 GND.n1478 GND.n1477 294.776
R2132 GND.n1437 GND.n296 291.205
R2133 GND.t911 GND.t594 290.19
R2134 GND.t400 GND.t823 290.19
R2135 GND.t640 GND.t395 290.19
R2136 GND.n1412 GND.n1411 289.13
R2137 GND.n1813 GND.n155 281.976
R2138 GND.n1814 GND.n1813 281.976
R2139 GND.n158 GND.n157 281.976
R2140 GND.n1472 GND.n271 281.601
R2141 GND.n1777 GND.n155 281.601
R2142 GND.n1778 GND.n1777 281.601
R2143 GND.n157 GND.n154 281.601
R2144 GND.n1814 GND.n154 281.601
R2145 GND.n1815 GND.n1814 281.601
R2146 GND.n1815 GND.n148 281.601
R2147 GND.n160 GND.n155 281.601
R2148 GND.t475 GND.t138 280.075
R2149 GND.t377 GND.t419 280.075
R2150 GND.t539 GND.n22 279.555
R2151 GND.n1771 GND.n1748 278.966
R2152 GND.n1710 GND.n1709 278.966
R2153 GND.n182 GND.n178 278.966
R2154 GND.n1700 GND.n182 278.966
R2155 GND.n180 GND.n179 278.966
R2156 GND.n179 GND.n25 278.966
R2157 GND.t816 GND.t798 275.68
R2158 GND.t398 GND.t936 275.68
R2159 GND.t14 GND.t399 275.68
R2160 GND.n1233 GND.t874 274.812
R2161 GND.n1261 GND.t765 274.812
R2162 GND.n527 GND.t178 274.812
R2163 GND.n516 GND.t562 274.812
R2164 GND.n180 GND.n19 274.072
R2165 GND.n1618 GND.n178 274.072
R2166 GND.n1133 GND.n1132 272.565
R2167 GND.t839 GND 269.733
R2168 GND.t556 GND 269.733
R2169 GND.n1759 GND.t71 263.688
R2170 GND.n1574 GND.n1573 259.873
R2171 GND.n311 GND.n310 259.765
R2172 GND GND.t821 256.853
R2173 GND.n1461 GND.n281 256.753
R2174 GND.t594 GND 253.917
R2175 GND.t564 GND 253.917
R2176 GND.t385 GND 253.917
R2177 GND.t823 GND 253.917
R2178 GND GND.t576 253.917
R2179 GND GND.t826 253.917
R2180 GND GND.t640 253.917
R2181 GND GND.t835 253.917
R2182 GND GND.t727 253.917
R2183 GND.n584 GND.n583 253.26
R2184 GND GND.t863 252.875
R2185 GND.t406 GND 252.875
R2186 GND.t141 GND 252.875
R2187 GND.n588 GND.n201 251.339
R2188 GND.n590 GND.n589 249.207
R2189 GND.t576 GND.n610 246.237
R2190 GND.n1613 GND.t65 242.832
R2191 GND.n1325 GND.t746 242.202
R2192 GND.n1447 GND.n292 241.319
R2193 GND.n318 GND.n248 241.319
R2194 GND.n1478 GND.n264 240.565
R2195 GND.n1481 GND.n261 240.565
R2196 GND.n1471 GND.n272 237.177
R2197 GND.t873 GND 236.016
R2198 GND.n1397 GND.n1396 235.98
R2199 GND.n1467 GND.n272 235.672
R2200 GND GND.t833 232.153
R2201 GND.t912 GND.n609 232.153
R2202 GND.n698 GND.t398 232.153
R2203 GND.t925 GND 232.153
R2204 GND.n620 GND.t913 232.153
R2205 GND.t399 GND.n663 232.153
R2206 GND.t85 GND 232.153
R2207 GND.n680 GND.t394 232.153
R2208 GND.n668 GND.t816 230.849
R2209 GND.n592 GND.n591 229.579
R2210 GND.n1858 GND.n22 228.679
R2211 GND.n667 GND.t524 228.524
R2212 GND.t17 GND.n664 228.524
R2213 GND.t907 GND.t908 228.131
R2214 GND.t904 GND.t152 228.131
R2215 GND.n587 GND.n586 226.544
R2216 GND.n314 GND.n250 226.26
R2217 GND.t662 GND.t137 225.698
R2218 GND.t371 GND.t20 224.898
R2219 GND.t557 GND.t902 224.898
R2220 GND.t945 GND.t502 224.898
R2221 GND.n1665 GND.t268 222.456
R2222 GND.n174 GND.t359 222.456
R2223 GND.n170 GND.t236 222.456
R2224 GND.n1723 GND.t243 222.456
R2225 GND.n1719 GND.t308 222.456
R2226 GND.n1644 GND.t275 222.456
R2227 GND.n1639 GND.t196 222.456
R2228 GND.n1662 GND.t356 222.456
R2229 GND.n35 GND.t295 222.452
R2230 GND.n47 GND.t317 222.452
R2231 GND.n1674 GND.t322 222.452
R2232 GND.n173 GND.t293 222.452
R2233 GND.n169 GND.t328 222.452
R2234 GND.n1724 GND.t183 222.452
R2235 GND.n1720 GND.t239 222.452
R2236 GND.n1688 GND.t352 222.452
R2237 GND.n51 GND.t298 222.379
R2238 GND.n38 GND.t225 222.379
R2239 GND.n1838 GND.t299 222.355
R2240 GND.n39 GND.t224 222.355
R2241 GND.n53 GND.t341 222.297
R2242 GND.n55 GND.t218 222.297
R2243 GND.n1 GND.t340 222.263
R2244 GND.n57 GND.t219 222.263
R2245 GND.n1621 GND.t192 222.228
R2246 GND.n1621 GND.t191 222.228
R2247 GND.n1619 GND.t290 222.228
R2248 GND.n1619 GND.t289 222.228
R2249 GND.n165 GND.t337 222.228
R2250 GND.n165 GND.t336 222.228
R2251 GND.n1691 GND.t207 222.228
R2252 GND.n1691 GND.t206 222.228
R2253 GND.n439 GND.t146 222.188
R2254 GND.n298 GND.t699 222.023
R2255 GND.n298 GND.t701 221.905
R2256 GND.n290 GND.t494 221.851
R2257 GND.n290 GND.t700 221.851
R2258 GND.n31 GND.t948 221.851
R2259 GND.n31 GND.t978 221.851
R2260 GND.n1659 GND.t444 221.851
R2261 GND.n1659 GND.t262 221.851
R2262 GND.n1667 GND.t69 221.851
R2263 GND.n1667 GND.t320 221.851
R2264 GND.n1663 GND.t261 221.851
R2265 GND.n1663 GND.t357 221.851
R2266 GND.n1666 GND.t319 221.851
R2267 GND.n1666 GND.t269 221.851
R2268 GND.n36 GND.t31 221.851
R2269 GND.n36 GND.t296 221.851
R2270 GND.n34 GND.t470 221.851
R2271 GND.n34 GND.t33 221.851
R2272 GND.n33 GND.t585 221.851
R2273 GND.n33 GND.t453 221.851
R2274 GND.n32 GND.t477 221.851
R2275 GND.n32 GND.t467 221.851
R2276 GND.n44 GND.t447 221.851
R2277 GND.n44 GND.t949 221.851
R2278 GND.n45 GND.t947 221.851
R2279 GND.n45 GND.t134 221.851
R2280 GND.n46 GND.t980 221.851
R2281 GND.n46 GND.t439 221.851
R2282 GND.n48 GND.t316 221.851
R2283 GND.n48 GND.t981 221.851
R2284 GND.n1675 GND.t583 221.851
R2285 GND.n1675 GND.t323 221.851
R2286 GND.n1678 GND.t66 221.851
R2287 GND.n1678 GND.t586 221.851
R2288 GND.n1680 GND.t478 221.851
R2289 GND.n1680 GND.t476 221.851
R2290 GND.n1682 GND.t70 221.851
R2291 GND.n1682 GND.t62 221.851
R2292 GND.n171 GND.t327 221.851
R2293 GND.n171 GND.t237 221.851
R2294 GND.n175 GND.t292 221.851
R2295 GND.n175 GND.t360 221.851
R2296 GND.n1721 GND.t307 221.851
R2297 GND.n1721 GND.t240 221.851
R2298 GND.n1725 GND.t242 221.851
R2299 GND.n1725 GND.t184 221.851
R2300 GND.n1684 GND.t133 221.851
R2301 GND.n1684 GND.t445 221.851
R2302 GND.n1685 GND.t953 221.851
R2303 GND.n1685 GND.t29 221.851
R2304 GND.n1686 GND.t982 221.851
R2305 GND.n1686 GND.t450 221.851
R2306 GND.n1687 GND.t448 221.851
R2307 GND.n1687 GND.t950 221.851
R2308 GND.n1689 GND.t351 221.851
R2309 GND.n1689 GND.t449 221.851
R2310 GND.n1640 GND.t195 221.851
R2311 GND.n1640 GND.t265 221.851
R2312 GND.n1645 GND.t274 221.851
R2313 GND.n1645 GND.t334 221.851
R2314 GND.n1638 GND.t264 221.851
R2315 GND.n1638 GND.t434 221.851
R2316 GND.n1648 GND.t333 221.851
R2317 GND.n1648 GND.t64 221.851
R2318 GND.n1630 GND.t976 221.851
R2319 GND.n1630 GND.t589 221.851
R2320 GND.n1631 GND.t474 221.851
R2321 GND.n1631 GND.t472 221.851
R2322 GND.n1632 GND.t435 221.851
R2323 GND.n1632 GND.t74 221.851
R2324 GND.n1633 GND.t68 221.851
R2325 GND.n1633 GND.t587 221.851
R2326 GND.n1634 GND.t72 221.851
R2327 GND.n1634 GND.t588 221.851
R2328 GND.n1635 GND.t451 221.851
R2329 GND.n1635 GND.t469 221.851
R2330 GND.n1624 GND.t951 221.851
R2331 GND.n1624 GND.t983 221.851
R2332 GND.n1625 GND.t590 221.851
R2333 GND.n1625 GND.t433 221.851
R2334 GND.n1626 GND.t979 221.851
R2335 GND.n1626 GND.t952 221.851
R2336 GND.n1627 GND.t430 221.851
R2337 GND.n1627 GND.t977 221.851
R2338 GND.n1628 GND.t431 221.851
R2339 GND.n1628 GND.t37 221.851
R2340 GND.n1629 GND.t35 221.851
R2341 GND.n1629 GND.t437 221.851
R2342 GND.n1459 GND.t397 221.738
R2343 GND.n1410 GND.n250 217.601
R2344 GND GND.n667 214.016
R2345 GND GND.n697 214.016
R2346 GND.n664 GND 214.016
R2347 GND.t798 GND.t531 210.387
R2348 GND.t833 GND.t563 210.387
R2349 GND.t936 GND.t743 210.387
R2350 GND.t376 GND.t925 210.387
R2351 GND.t425 GND.t14 210.387
R2352 GND.t884 GND.t85 210.387
R2353 GND.n359 GND.n358 207.393
R2354 GND.n671 GND.t49 205.118
R2355 GND.t801 GND.t132 204.843
R2356 GND.n1713 GND.t190 204.097
R2357 GND.n1764 GND.n1749 203.672
R2358 GND.n1770 GND.n1749 203.672
R2359 GND.n1763 GND.n1756 203.672
R2360 GND.n1756 GND.n1750 203.672
R2361 GND.n1863 GND.n13 203.672
R2362 GND.n1863 GND.n1862 203.672
R2363 GND.n1615 GND.n1606 203.672
R2364 GND.n1616 GND.n1615 203.672
R2365 GND.n1711 GND.n1710 203.672
R2366 GND.n314 GND.n248 202.542
R2367 GND.n1432 GND.n292 201.788
R2368 GND.n1091 GND.n1051 200.215
R2369 GND.n1091 GND.n1049 200.215
R2370 GND.n1091 GND.n1047 200.215
R2371 GND.n1091 GND.n1084 200.215
R2372 GND.t98 GND.t93 200.107
R2373 GND.n1595 GND.n188 197.272
R2374 GND.n1596 GND.n1595 197.272
R2375 GND.n580 GND.n197 196.726
R2376 GND.n491 GND.n485 196.256
R2377 GND.t103 GND.t385 195.879
R2378 GND.t826 GND.t499 195.879
R2379 GND.t727 GND.t39 195.879
R2380 GND.n332 GND.n321 195.766
R2381 GND.n1503 GND.n241 195.395
R2382 GND.n1587 GND.n1586 195
R2383 GND.n1588 GND.n1587 195
R2384 GND.t105 GND.t663 192.179
R2385 GND.t89 GND.t90 192.179
R2386 GND.n579 GND.n198 192.034
R2387 GND.n1392 GND.n1391 189.688
R2388 GND.t128 GND.t139 188.454
R2389 GND.n589 GND.n588 188.194
R2390 GND.t552 GND 185.441
R2391 GND.t124 GND 185.441
R2392 GND.n697 GND.n610 184.678
R2393 GND.n1075 GND.n1051 184.572
R2394 GND.n1066 GND.n1049 184.572
R2395 GND.n1057 GND.n1047 184.572
R2396 GND.n1084 GND.n1044 184.572
R2397 GND.n1520 GND.n229 184.471
R2398 GND.n1523 GND.n228 184.471
R2399 GND.n1526 GND.n227 184.471
R2400 GND.n1537 GND.n1530 184.471
R2401 GND.n1535 GND.n1534 184.471
R2402 GND.n1561 GND.n1560 184.471
R2403 GND.n1413 GND.n311 184.095
R2404 GND.t194 GND.n20 183.24
R2405 GND.n578 GND.t840 183.065
R2406 GND.n575 GND.t892 183.065
R2407 GND.n571 GND.t687 183.065
R2408 GND.n567 GND.t378 183.065
R2409 GND.n563 GND.t850 183.065
R2410 GND.n559 GND.t837 183.065
R2411 GND.n555 GND.t819 183.065
R2412 GND.n551 GND.t23 183.065
R2413 GND.n547 GND.t175 183.065
R2414 GND.n543 GND.t616 183.065
R2415 GND.n1387 GND.n1386 180.087
R2416 GND.n1703 GND.n1700 179.577
R2417 GND.n1703 GND.n1702 179.577
R2418 GND.n1856 GND.n25 179.577
R2419 GND.n1856 GND.n1855 179.577
R2420 GND.n593 GND.n592 179.019
R2421 GND.n1562 GND.n1561 179.004
R2422 GND.t559 GND.t140 178.68
R2423 GND.n1735 GND.t919 177.296
R2424 GND.n1734 GND.t462 177.296
R2425 GND.n1108 GND.n271 175.06
R2426 GND.n1855 GND.n1854 174.683
R2427 GND.n1702 GND.n1701 174.683
R2428 GND.n1522 GND.n1521 173.474
R2429 GND.n296 GND.n281 172.746
R2430 GND.n363 GND.n362 172.619
R2431 GND.t129 GND.t194 172.067
R2432 GND.n355 GND.n354 171.554
R2433 GND.n1347 GND.n1346 171.339
R2434 GND.n1377 GND.n1376 171.339
R2435 GND.n1398 GND.n1397 171.339
R2436 GND.n351 GND.n350 171.339
R2437 GND.n346 GND.n345 171.339
R2438 GND.n342 GND.n341 171.339
R2439 GND.n1138 GND.n1133 171.294
R2440 GND.n1383 GND.n1382 171.126
R2441 GND.n1533 GND.n202 170.487
R2442 GND.n1351 GND.n1350 170.274
R2443 GND.n1342 GND.n1341 170.274
R2444 GND.n1338 GND.n1337 170.274
R2445 GND.n1529 GND.n1528 170.274
R2446 GND.n337 GND.n336 170.274
R2447 GND.n1373 GND.n1372 170.06
R2448 GND.n422 GND.n420 168.282
R2449 GND.t815 GND.t416 167.599
R2450 GND.t487 GND.n1591 164.619
R2451 GND.n1592 GND.t109 164.619
R2452 GND.n1592 GND.t497 164.619
R2453 GND.n1571 GND.n1570 163.874
R2454 GND.n727 GND.t841 162.471
R2455 GND.n732 GND.t847 162.471
R2456 GND.n738 GND.t893 162.471
R2457 GND.n743 GND.t482 162.471
R2458 GND.n749 GND.t688 162.471
R2459 GND.n754 GND.t734 162.471
R2460 GND.n760 GND.t379 162.471
R2461 GND.n765 GND.t673 162.471
R2462 GND.n771 GND.t851 162.471
R2463 GND.n776 GND.t940 162.471
R2464 GND.n782 GND.t838 162.471
R2465 GND.n787 GND.t935 162.471
R2466 GND.n793 GND.t820 162.471
R2467 GND.n798 GND.t76 162.471
R2468 GND.n804 GND.t24 162.471
R2469 GND.n809 GND.t716 162.471
R2470 GND.n815 GND.t176 162.471
R2471 GND.n820 GND.t441 162.471
R2472 GND.n826 GND.t617 162.471
R2473 GND.n831 GND.t655 162.471
R2474 GND.n1834 GND.t217 162.389
R2475 GND.n1567 GND.n1565 161.903
R2476 GND.n1829 GND.n1828 161.882
R2477 GND.n1828 GND.n140 161.882
R2478 GND.n1586 GND.n186 161.506
R2479 GND GND.t846 161.149
R2480 GND GND.t481 161.149
R2481 GND GND.t733 161.149
R2482 GND GND.t672 161.149
R2483 GND GND.t939 161.149
R2484 GND GND.t934 161.149
R2485 GND GND.t75 161.149
R2486 GND GND.t715 161.149
R2487 GND GND.t440 161.149
R2488 GND GND.t654 161.149
R2489 GND.n731 GND.t510 160.017
R2490 GND.n574 GND.t849 160.017
R2491 GND.n742 GND.t895 160.017
R2492 GND.n570 GND.t484 160.017
R2493 GND.n753 GND.t690 160.017
R2494 GND.n566 GND.t857 160.017
R2495 GND.n764 GND.t381 160.017
R2496 GND.n562 GND.t675 160.017
R2497 GND.n775 GND.t853 160.017
R2498 GND.n558 GND.t942 160.017
R2499 GND.n786 GND.t883 160.017
R2500 GND.n554 GND.t891 160.017
R2501 GND.n797 GND.t818 160.017
R2502 GND.n550 GND.t78 160.017
R2503 GND.n808 GND.t26 160.017
R2504 GND.n546 GND.t718 160.017
R2505 GND.n819 GND.t171 160.017
R2506 GND.n542 GND.t538 160.017
R2507 GND.n540 GND.t866 160.017
R2508 GND.n833 GND.t512 160.017
R2509 GND.t520 GND.t907 159.571
R2510 GND.t908 GND.t753 159.571
R2511 GND.t152 GND.t809 159.571
R2512 GND.t581 GND.t904 159.571
R2513 GND.t725 GND.t147 159.571
R2514 GND.n1221 GND.t722 158.361
R2515 GND.n1228 GND.t374 158.361
R2516 GND.n376 GND.t542 158.361
R2517 GND.n378 GND.t961 158.361
R2518 GND.n497 GND.t523 158.361
R2519 GND.n1300 GND.t800 155.63
R2520 GND.n1413 GND.n1412 154.73
R2521 GND.n1298 GND.t11 154.131
R2522 GND.n1275 GND.t886 154.131
R2523 GND.n1055 GND.t620 153.707
R2524 GND.n1277 GND.t724 153.631
R2525 GND.n863 GND.n862 153.276
R2526 GND.t875 GND.t803 152.794
R2527 GND.n1278 GND.t671 152.381
R2528 GND.n1532 GND.n1531 152.139
R2529 GND.n1527 GND.n1526 151.779
R2530 GND.n1240 GND 151.725
R2531 GND.n357 GND.n356 151.714
R2532 GND.n1349 GND.n1348 151.5
R2533 GND.n1340 GND.n1339 151.5
R2534 GND.n1375 GND.n1374 151.5
R2535 GND.n1525 GND.n1524 151.5
R2536 GND.n344 GND.n343 151.5
R2537 GND.n340 GND.n339 151.5
R2538 GND.n490 GND.n489 151.256
R2539 GND.n491 GND.n490 151.256
R2540 GND.n488 GND.n487 151.256
R2541 GND.n489 GND.n488 151.256
R2542 GND.n486 GND.n471 151.256
R2543 GND.n487 GND.n486 151.256
R2544 GND.n474 GND.n469 151.256
R2545 GND.n474 GND.n471 151.256
R2546 GND.n468 GND.n467 151.256
R2547 GND.n469 GND.n468 151.256
R2548 GND.n466 GND.n465 151.256
R2549 GND.n467 GND.n466 151.256
R2550 GND.n856 GND.n452 151.256
R2551 GND.n465 GND.n452 151.256
R2552 GND.n859 GND.n449 151.256
R2553 GND.n859 GND.n858 151.256
R2554 GND.n858 GND.n857 151.256
R2555 GND.n857 GND.n856 151.256
R2556 GND.n862 GND.n449 151.256
R2557 GND.t814 GND.t190 151.21
R2558 GND.n1244 GND.t830 150.922
R2559 GND.n1248 GND.t553 150.922
R2560 GND.n1249 GND.t121 150.922
R2561 GND.n1235 GND.t868 150.922
R2562 GND.n1234 GND.t127 150.922
R2563 GND.n1305 GND.t560 150.922
R2564 GND.n1293 GND.t414 150.922
R2565 GND.n1289 GND.t822 150.922
R2566 GND.n1284 GND.t174 150.922
R2567 GND.n1243 GND.t125 150.922
R2568 GND.n510 GND.t957 150.922
R2569 GND.n505 GND.t550 150.922
R2570 GND.n633 GND.t558 150.922
R2571 GND.n716 GND.t372 150.922
R2572 GND.n703 GND.t386 150.922
R2573 GND.n709 GND.t565 150.922
R2574 GND.n603 GND.t595 150.922
R2575 GND.n641 GND.t577 150.922
R2576 GND.n647 GND.t827 150.922
R2577 GND.n684 GND.t728 150.922
R2578 GND.n690 GND.t836 150.922
R2579 GND.n652 GND.t641 150.922
R2580 GND.n657 GND.t503 150.922
R2581 GND.n635 GND.t824 150.922
R2582 GND.n353 GND.n352 150.434
R2583 GND.n1300 GND.t123 149.493
R2584 GND.n1218 GND.t651 149.493
R2585 GND.n1400 GND.n320 149.367
R2586 GND.n1479 GND.n1478 149.083
R2587 GND.n1062 GND.t682 149.067
R2588 GND.n1071 GND.t609 149.067
R2589 GND.n1080 GND.t712 149.067
R2590 GND.n871 GND.t59 149.067
R2591 GND.n881 GND.t4 149.067
R2592 GND.n891 GND.t736 149.067
R2593 GND.n1015 GND.t669 149.067
R2594 GND.n903 GND.t593 149.067
R2595 GND.n913 GND.t492 149.067
R2596 GND.n923 GND.t645 149.067
R2597 GND.n987 GND.t461 149.067
R2598 GND.n935 GND.t518 149.067
R2599 GND.n945 GND.t421 149.067
R2600 GND.n954 GND.t489 149.067
R2601 GND.n959 GND.t889 149.067
R2602 GND.n403 GND.t756 149.067
R2603 GND.n1200 GND.t697 149.067
R2604 GND.n1189 GND.t580 149.067
R2605 GND.n1153 GND.t720 149.067
R2606 GND.n1174 GND.t679 149.067
R2607 GND.n1162 GND.t845 149.067
R2608 GND.n1385 GND.n1384 148.087
R2609 GND.n1307 GND.t143 147.411
R2610 GND.n1559 GND.n1558 146.25
R2611 GND.n1558 GND.n194 146.25
R2612 GND.n312 GND.n309 146.25
R2613 GND.n317 GND.n309 146.25
R2614 GND.n1409 GND.n1408 146.25
R2615 GND.n1408 GND.n1407 146.25
R2616 GND.n1404 GND.n1403 146.25
R2617 GND.n1405 GND.n1404 146.25
R2618 GND.n325 GND.n322 146.25
R2619 GND.n324 GND.n322 146.25
R2620 GND.n323 GND.n321 146.25
R2621 GND.n213 GND.n212 146.25
R2622 GND.n1510 GND.n213 146.25
R2623 GND.n222 GND.n211 146.25
R2624 GND.n223 GND.n222 146.25
R2625 GND.n1555 GND.n1554 146.25
R2626 GND.n1556 GND.n1555 146.25
R2627 GND.n1514 GND.n1513 146.25
R2628 GND.n1515 GND.n1514 146.25
R2629 GND.n1509 GND.n1508 146.25
R2630 GND.n1510 GND.n1509 146.25
R2631 GND.n225 GND.n217 146.25
R2632 GND.n225 GND.n224 146.25
R2633 GND.n431 GND.n430 146.25
R2634 GND.n430 GND.n236 146.25
R2635 GND.n262 GND.n258 146.25
R2636 GND.n260 GND.n258 146.25
R2637 GND.n259 GND.n256 146.25
R2638 GND.n259 GND.n238 146.25
R2639 GND.n1135 GND.n252 146.25
R2640 GND.n1123 GND.n252 146.25
R2641 GND.n253 GND.n249 146.25
R2642 GND.n254 GND.n253 146.25
R2643 GND.n247 GND.n243 146.25
R2644 GND.n243 GND.n241 146.25
R2645 GND.n1134 GND.n1125 146.25
R2646 GND.n1125 GND.n1124 146.25
R2647 GND.n1499 GND.n244 146.25
R2648 GND.n1147 GND.n1146 146.25
R2649 GND.n1086 GND.n1085 146.25
R2650 GND.n1087 GND.n1086 146.25
R2651 GND.n1421 GND.n1420 146.25
R2652 GND.n1422 GND.n1421 146.25
R2653 GND.n308 GND.n305 146.25
R2654 GND.n308 GND.n307 146.25
R2655 GND.n1104 GND.n421 146.25
R2656 GND.n1105 GND.n1104 146.25
R2657 GND.n1121 GND.n424 146.25
R2658 GND.n1121 GND.n1120 146.25
R2659 GND.n266 GND.n265 146.25
R2660 GND.n1088 GND.n266 146.25
R2661 GND.n267 GND.n263 146.25
R2662 GND.n1423 GND.n267 146.25
R2663 GND.n434 GND.n433 146.25
R2664 GND.n435 GND.n434 146.25
R2665 GND.n1453 GND.n1452 146.25
R2666 GND.n1454 GND.n1453 146.25
R2667 GND.n1308 GND.t555 146.245
R2668 GND.t540 GND.n1866 145.504
R2669 GND.n1330 GND.t9 144.454
R2670 GND.n591 GND.n590 143.393
R2671 GND.n361 GND.n360 142.754
R2672 GND.n1833 GND.t93 142.712
R2673 GND.n1830 GND.n1829 142.683
R2674 GND.n1817 GND.n140 142.683
R2675 GND.t132 GND.n10 140.037
R2676 GND.n1836 GND.n133 139.294
R2677 GND.n1524 GND.n1523 138.897
R2678 GND.t661 GND.t36 137.804
R2679 GND.n844 GND.t958 137.728
R2680 GND.n1345 GND.n1344 137.47
R2681 GND.n1337 GND.n1335 137.419
R2682 GND.n358 GND.n333 135.286
R2683 GND.n1733 GND.n22 135.083
R2684 GND.n586 GND.n585 135.073
R2685 GND.n423 GND.n422 133.272
R2686 GND.n1531 GND.n1530 133.137
R2687 GND.n1379 GND.n1378 132.907
R2688 GND.n1790 GND.t228 132.465
R2689 GND.n146 GND.t231 132.465
R2690 GND.n1796 GND.t250 132.465
R2691 GND.n1802 GND.t248 132.465
R2692 GND.n1572 GND.n1571 132.071
R2693 GND.n1521 GND.n1520 131.857
R2694 GND.n1130 GND.n419 130.26
R2695 GND.t137 GND.n1865 129.609
R2696 GND.n360 GND.n359 128.887
R2697 GND.t260 GND.t814 128.864
R2698 GND.n1097 GND.t969 127.977
R2699 GND.n1599 GND.n183 125.885
R2700 GND.n1534 GND.n1533 125.457
R2701 GND.t522 GND 125.046
R2702 GND.n1038 GND.n866 121.496
R2703 GND.n1561 GND.n202 120.55
R2704 GND.n1809 GND.t229 119.444
R2705 GND.t232 GND.n1819 119.444
R2706 GND.n581 GND.n579 117.99
R2707 GND.t109 GND.t487 117.692
R2708 GND.t497 GND.t455 117.692
R2709 GND.n1103 GND.n1102 117.001
R2710 GND.n1110 GND.n1103 117.001
R2711 GND.n442 GND.n441 117.001
R2712 GND.n1110 GND.n441 117.001
R2713 GND.n1443 GND.n1442 117.001
R2714 GND.n1444 GND.n1443 117.001
R2715 GND.n1456 GND.n1455 117.001
R2716 GND.n1455 GND.n1454 117.001
R2717 GND.n1111 GND.n446 117.001
R2718 GND.n1111 GND.n1110 117.001
R2719 GND.n1118 GND.n1117 117.001
R2720 GND.n1119 GND.n1118 117.001
R2721 GND.t802 GND.t28 116.947
R2722 GND.n1554 GND.n210 114.825
R2723 GND.t65 GND.t815 112.478
R2724 GND.n1436 GND.n292 111.812
R2725 GND.n1523 GND.n1522 110.311
R2726 GND.t563 GND.t103 108.822
R2727 GND.t499 GND.t376 108.822
R2728 GND.t39 GND.t884 108.822
R2729 GND.n1669 GND.t318 108.365
R2730 GND.n1665 GND.t266 108.365
R2731 GND.n52 GND.t338 108.365
R2732 GND.n56 GND.t216 108.365
R2733 GND.n51 GND.t297 108.365
R2734 GND.n38 GND.t222 108.365
R2735 GND.n35 GND.t294 108.365
R2736 GND.n47 GND.t315 108.365
R2737 GND.n1621 GND.t189 108.365
R2738 GND.n1674 GND.t321 108.365
R2739 GND.n1619 GND.t288 108.365
R2740 GND.n165 GND.t335 108.365
R2741 GND.n174 GND.t358 108.365
R2742 GND.n173 GND.t291 108.365
R2743 GND.n170 GND.t235 108.365
R2744 GND.n169 GND.t326 108.365
R2745 GND.n1724 GND.t181 108.365
R2746 GND.n1723 GND.t241 108.365
R2747 GND.n1720 GND.t238 108.365
R2748 GND.n1719 GND.t306 108.365
R2749 GND.n1688 GND.t350 108.365
R2750 GND.n1691 GND.t205 108.365
R2751 GND.n1644 GND.t272 108.365
R2752 GND.n1642 GND.t263 108.365
R2753 GND.n1647 GND.t331 108.365
R2754 GND.n1639 GND.t193 108.365
R2755 GND.n1662 GND.t355 108.365
R2756 GND.n1661 GND.t259 108.365
R2757 GND.t840 GND.t509 108.293
R2758 GND.t846 GND.t848 108.293
R2759 GND.t892 GND.t894 108.293
R2760 GND.t481 GND.t483 108.293
R2761 GND.t687 GND.t689 108.293
R2762 GND.t733 GND.t856 108.293
R2763 GND.t378 GND.t380 108.293
R2764 GND.t672 GND.t674 108.293
R2765 GND.t850 GND.t852 108.293
R2766 GND.t939 GND.t941 108.293
R2767 GND.t837 GND.t882 108.293
R2768 GND.t934 GND.t890 108.293
R2769 GND.t819 GND.t817 108.293
R2770 GND.t75 GND.t77 108.293
R2771 GND.t23 GND.t25 108.293
R2772 GND.t715 GND.t717 108.293
R2773 GND.t175 GND.t170 108.293
R2774 GND.t440 GND.t537 108.293
R2775 GND.t616 GND.t865 108.293
R2776 GND.t654 GND.t511 108.293
R2777 GND.t182 GND.t129 108.007
R2778 GND.n1534 GND.n1532 106.257
R2779 GND.n679 GND.n450 106.16
R2780 GND.n1388 GND.n1387 102.433
R2781 GND.n501 GND.t864 102.377
R2782 GND.n191 GND.n188 101.647
R2783 GND.n1570 GND 100.496
R2784 GND.n1399 GND.n1398 100.299
R2785 GND.n1580 GND.t877 100.053
R2786 GND.n1396 GND.n1395 99.6436
R2787 GND.n1116 GND.n1115 99.3887
R2788 GND.t57 GND.n240 99.2212
R2789 GND.n1386 GND.n1385 98.1667
R2790 GND GND.n575 96.6896
R2791 GND GND.n571 96.6896
R2792 GND GND.n567 96.6896
R2793 GND GND.n563 96.6896
R2794 GND GND.n559 96.6896
R2795 GND GND.n555 96.6896
R2796 GND GND.n551 96.6896
R2797 GND GND.n547 96.6896
R2798 GND GND.n543 96.6896
R2799 GND.n1530 GND.n1529 96.4436
R2800 GND.n1317 GND.n1316 96.2411
R2801 GND.n1612 GND.t813 96.0899
R2802 GND.t417 GND.n1612 96.0899
R2803 GND.n1760 GND.t802 96.0899
R2804 GND.n1767 GND.t130 96.0899
R2805 GND.n1767 GND.t418 96.0899
R2806 GND.n336 GND.n320 96.0333
R2807 GND.n1448 GND.n288 95.2476
R2808 GND.t531 GND.t371 94.3121
R2809 GND.t743 GND.t557 94.3121
R2810 GND.t502 GND.t425 94.3121
R2811 GND.t71 GND.t128 91.6206
R2812 GND.t614 GND 89.9457
R2813 GND.n677 GND.n676 89.504
R2814 GND GND.t831 89.2144
R2815 GND.n1526 GND.n1525 88.9769
R2816 GND.n862 GND.n861 88.7516
R2817 GND.t91 GND.n1578 88.4193
R2818 GND.n1866 GND.t661 87.1513
R2819 GND.t509 GND 86.3761
R2820 GND.t848 GND 86.3761
R2821 GND.t894 GND 86.3761
R2822 GND.t483 GND 86.3761
R2823 GND.t689 GND 86.3761
R2824 GND.t856 GND 86.3761
R2825 GND.t380 GND 86.3761
R2826 GND.t674 GND 86.3761
R2827 GND.t852 GND 86.3761
R2828 GND.t941 GND 86.3761
R2829 GND.t882 GND 86.3761
R2830 GND.t890 GND 86.3761
R2831 GND.t817 GND 86.3761
R2832 GND.t77 GND 86.3761
R2833 GND.t25 GND 86.3761
R2834 GND.t717 GND 86.3761
R2835 GND.t170 GND 86.3761
R2836 GND.t537 GND 86.3761
R2837 GND.t865 GND 86.3761
R2838 GND.t511 GND 86.3761
R2839 GND.n844 GND 86.3761
R2840 GND.n1832 GND.n134 86.0925
R2841 GND.n1591 GND.n190 85.6616
R2842 GND.n1364 GND.t0 85.3595
R2843 GND.n362 GND.n361 84.94
R2844 GND.t418 GND.t182 84.1718
R2845 GND.n144 GND.t876 83.4151
R2846 GND.n142 GND.t878 83.4151
R2847 GND.n141 GND.t880 83.4151
R2848 GND.n1826 GND.t879 83.4151
R2849 GND.n1339 GND.n1338 82.8067
R2850 GND.n1341 GND.n1340 80.6733
R2851 GND.n1809 GND.t98 80.6633
R2852 GND.n1819 GND.t803 80.6633
R2853 GND.n1395 GND.n332 80.0005
R2854 GND.n1402 GND.n1400 80.0005
R2855 GND GND.t522 77.5142
R2856 GND.t28 GND.t801 75.2333
R2857 GND.n1710 GND.n1617 74.7248
R2858 GND.n1617 GND.n1616 74.7248
R2859 GND.n1616 GND.n14 74.7248
R2860 GND.n1862 GND.n14 74.7248
R2861 GND.n1750 GND.n16 74.7248
R2862 GND.n1769 GND.n1750 74.7248
R2863 GND.n1770 GND.n1769 74.7248
R2864 GND.n1366 GND.t18 74.416
R2865 GND.n1786 GND.n1778 74.3199
R2866 GND.n1786 GND.n148 74.3199
R2867 GND.n1403 GND.n1402 74.0272
R2868 GND.n1861 GND.n16 73.514
R2869 GND.n186 GND.n184 73.1255
R2870 GND.n192 GND.n184 73.1255
R2871 GND.n1589 GND.n191 73.1255
R2872 GND.t135 GND.t117 72.1616
R2873 GND.t136 GND.t166 72.1616
R2874 GND.t156 GND.t136 72.1616
R2875 GND.t164 GND.t156 72.1616
R2876 GND.t158 GND.t164 72.1616
R2877 GND.t116 GND.t158 72.1616
R2878 GND.t160 GND.t116 72.1616
R2879 GND.t160 GND.t118 72.1616
R2880 GND.t118 GND.t165 72.1616
R2881 GND.t165 GND.t159 72.1616
R2882 GND.t159 GND.t163 72.1616
R2883 GND.t161 GND.t119 72.1616
R2884 GND.t119 GND.t162 72.1616
R2885 GND.t162 GND.t157 72.1616
R2886 GND.t737 GND.t404 72.1616
R2887 GND.t404 GND.t114 72.1616
R2888 GND.t114 GND.t707 72.1616
R2889 GND.t403 GND.t702 72.1616
R2890 GND.t792 GND.t779 72.1616
R2891 GND.t779 GND.t783 72.1616
R2892 GND.t783 GND.t791 72.1616
R2893 GND.n1384 GND.n1383 72.14
R2894 GND.n1382 GND.n1381 72.14
R2895 GND.n341 GND.n340 72.14
R2896 GND.n247 GND.n245 70.4005
R2897 GND.n1496 GND.n247 70.4005
R2898 GND.n1489 GND.n249 70.4005
R2899 GND.n1495 GND.n249 70.4005
R2900 GND.n1136 GND.n1135 70.4005
R2901 GND.n1135 GND.n251 70.4005
R2902 GND.n1508 GND.n1507 70.4005
R2903 GND.n1508 GND.n218 70.4005
R2904 GND.n1536 GND.n217 70.4005
R2905 GND.n1542 GND.n217 70.4005
R2906 GND.n216 GND.n212 70.4005
R2907 GND.n1545 GND.n211 70.4005
R2908 GND.n1552 GND.n211 70.4005
R2909 GND.n1403 GND.n318 70.4005
R2910 GND.n326 GND.n325 70.4005
R2911 GND.n325 GND.n319 70.4005
R2912 GND.n1420 GND.n303 70.4005
R2913 GND.n1420 GND.n1419 70.4005
R2914 GND.n310 GND.n305 70.4005
R2915 GND.n1418 GND.n305 70.4005
R2916 GND.n1411 GND.n312 70.4005
R2917 GND.n312 GND.n306 70.4005
R2918 GND.n1410 GND.n1409 70.4005
R2919 GND.n1409 GND.n313 70.4005
R2920 GND.n431 GND.n261 70.4005
R2921 GND.n433 GND.n264 70.4005
R2922 GND.n1479 GND.n263 70.4005
R2923 GND.n1127 GND.n263 70.4005
R2924 GND.n1480 GND.n262 70.4005
R2925 GND.n262 GND.n257 70.4005
R2926 GND.n1487 GND.n256 70.4005
R2927 GND.n1129 GND.n265 70.4005
R2928 GND.n1137 GND.n1134 70.4005
R2929 GND.n1134 GND.n425 70.4005
R2930 GND.n1132 GND.n424 70.4005
R2931 GND.n1143 GND.n424 70.4005
R2932 GND.n1131 GND.n421 70.4005
R2933 GND.n1144 GND.n421 70.4005
R2934 GND.n1499 GND.n1498 70.4005
R2935 GND.t938 GND.t825 70.2016
R2936 GND.t466 GND.t614 70.2016
R2937 GND.n581 GND.n580 69.7769
R2938 GND.n388 GND.t541 69.7227
R2939 GND.n1217 GND 69.4703
R2940 GND.t166 GND.t167 69.0242
R2941 GND.n354 GND.n353 67.4467
R2942 GND.t27 GND.t764 67.4335
R2943 GND.t547 GND.t120 67.4335
R2944 GND.t172 GND.t829 67.4335
R2945 GND.n1319 GND.n367 67.2766
R2946 GND.n1760 GND.t73 67.0396
R2947 GND.n1328 GND.n363 66.9708
R2948 GND.n1516 GND.n231 65.8868
R2949 GND.n338 GND.n337 65.3297
R2950 GND.n1343 GND.n1342 65.3133
R2951 GND.n356 GND.n355 65.3133
R2952 GND.n1101 GND.n447 65.1299
R2953 GND.n387 GND 65.0093
R2954 GND.n1436 GND.n1435 65.0005
R2955 GND.n1435 GND.n1434 65.0005
R2956 GND.t571 GND.t115 64.841
R2957 GND.t708 GND.t53 64.841
R2958 GND.t50 GND.t401 64.841
R2959 GND.t887 GND.n1733 64.7271
R2960 GND.n1456 GND.n285 64.377
R2961 GND.n446 GND.n271 64.0005
R2962 GND.n442 GND.n437 64.0005
R2963 GND.n442 GND.n280 64.0005
R2964 GND.n1456 GND.n281 64.0005
R2965 GND.n1117 GND.n272 64.0005
R2966 GND.n446 GND.n437 63.624
R2967 GND.n1117 GND.n1116 63.624
R2968 GND.t813 GND.t260 63.3152
R2969 GND.n1346 GND.n1345 63.18
R2970 GND.n345 GND.n344 63.18
R2971 GND.t177 GND.t938 61.4265
R2972 GND.t561 GND.t466 61.4265
R2973 GND.t864 GND.t956 61.4265
R2974 GND.t831 GND.t549 61.4265
R2975 GND.n1378 GND.n1377 61.0467
R2976 GND.n1376 GND.n1375 61.0467
R2977 GND.n343 GND.n342 61.0467
R2978 GND.n1442 GND.n296 60.6123
R2979 GND.n1367 GND.t19 60.5543
R2980 GND.n1102 GND.n280 60.2358
R2981 GND.t51 GND.n235 60.1348
R2982 GND.n1742 GND.t927 59.6649
R2983 GND.n1739 GND.t507 59.6649
R2984 GND.n1803 GND.t249 59.4285
R2985 GND.n147 GND.t252 59.4285
R2986 GND.n1823 GND.t234 59.4285
R2987 GND.n1791 GND.t230 59.4285
R2988 GND.n1348 GND.n1347 58.9133
R2989 GND.n352 GND.n351 58.9133
R2990 GND.n350 GND.n349 58.9133
R2991 GND.t90 GND.t377 58.8459
R2992 GND.n1831 GND.n1830 58.5005
R2993 GND.n1832 GND.n1831 58.5005
R2994 GND.n1818 GND.n1817 58.5005
R2995 GND.n1819 GND.n1818 58.5005
R2996 GND.n1836 GND.n1835 58.5005
R2997 GND.n1835 GND.n1834 58.5005
R2998 GND.n1869 GND.n1868 58.5005
R2999 GND.n1868 GND.n1867 58.5005
R3000 GND.t706 GND.t630 57.5203
R3001 GND.t113 GND.t534 57.5203
R3002 GND.t402 GND.t683 57.5203
R3003 GND.t112 GND.t533 57.5203
R3004 GND.t622 GND.t915 56.9878
R3005 GND.n1350 GND.n1349 56.78
R3006 GND.t872 GND.n161 56.2845
R3007 GND.n1515 GND.t117 55.6901
R3008 GND.t157 GND.n1510 55.6901
R3009 GND.n501 GND 55.5764
R3010 GND.t15 GND.n666 55.0318
R3011 GND.n666 GND.t638 55.0318
R3012 GND.n853 GND.t896 55.0318
R3013 GND.n853 GND.t382 55.0318
R3014 GND.t568 GND.n852 55.0318
R3015 GND.n852 GND.t691 55.0318
R3016 GND.t1 GND.n851 55.0318
R3017 GND.n851 GND.t869 55.0318
R3018 GND.n475 GND.t773 55.0318
R3019 GND.n475 GND.t842 55.0318
R3020 GND.n845 GND.t543 55.0318
R3021 GND.n845 GND.t943 55.0318
R3022 GND.t785 GND.t900 54.9057
R3023 GND.t790 GND.t84 54.9057
R3024 GND.n389 GND 54.7689
R3025 GND.n1374 GND.n1373 54.6467
R3026 GND.n1372 GND.n1371 54.6467
R3027 GND.n347 GND.n346 54.6467
R3028 GND.t36 GND.t662 54.3767
R3029 GND GND.n367 54.1138
R3030 GND.n1736 GND.n1730 53.1823
R3031 GND.n1736 GND.n1735 53.1823
R3032 GND.n1744 GND.n1732 53.1823
R3033 GND.n1735 GND.n1732 53.1823
R3034 GND.n137 GND.n135 53.1823
R3035 GND.n1579 GND.n135 53.1823
R3036 GND.n1828 GND.n136 53.1823
R3037 GND.n1580 GND.n136 53.1823
R3038 GND.t101 GND.n1580 52.7416
R3039 GND.n1352 GND.n1351 52.0867
R3040 GND.t780 GND.t693 52.0297
R3041 GND.t956 GND 51.1888
R3042 GND.t549 GND 51.1888
R3043 GND.t703 GND.t618 50.1996
R3044 GND.t914 GND.t786 50.1996
R3045 GND.t663 GND.t61 49.9074
R3046 GND.n1800 GND.n1793 49.3146
R3047 GND.n1798 GND.n1794 49.3146
R3048 GND.n1784 GND.n1781 49.3146
R3049 GND.n1788 GND.n1780 49.3146
R3050 GND.n1783 GND.n1782 49.1993
R3051 GND.n1801 GND.n1792 49.0972
R3052 GND.n1797 GND.n1795 49.0972
R3053 GND.n1789 GND.n1779 49.0972
R3054 GND.t875 GND.t101 47.3123
R3055 GND GND.t177 46.8012
R3056 GND GND.t561 46.8012
R3057 GND.n1452 GND.n288 46.3064
R3058 GND.t61 GND.n9 46.183
R3059 GND.t707 GND.t12 46.0163
R3060 GND.t660 GND.t95 45.7611
R3061 GND.t501 GND.t91 45.7611
R3062 GND.n675 GND.n672 45.7159
R3063 GND.n456 GND.n454 45.7159
R3064 GND.n855 GND.n854 45.7159
R3065 GND.n464 GND.n457 45.7159
R3066 GND.n850 GND.n849 45.7159
R3067 GND.n848 GND.n461 45.7159
R3068 GND.n847 GND.n846 45.7159
R3069 GND.n483 GND.n473 45.7159
R3070 GND.n841 GND.n840 45.7159
R3071 GND.n839 GND.n480 45.7159
R3072 GND.n1452 GND.n285 45.5534
R3073 GND.n666 GND.n456 45.0005
R3074 GND.n854 GND.n853 45.0005
R3075 GND.n852 GND.n457 45.0005
R3076 GND.n851 GND.n850 45.0005
R3077 GND.n475 GND.n461 45.0005
R3078 GND.n846 GND.n845 45.0005
R3079 GND.n857 GND.n451 45.0005
R3080 GND.n666 GND.n451 45.0005
R3081 GND.n458 GND.n452 45.0005
R3082 GND.n853 GND.n458 45.0005
R3083 GND.n466 GND.n459 45.0005
R3084 GND.n852 GND.n459 45.0005
R3085 GND.n468 GND.n460 45.0005
R3086 GND.n851 GND.n460 45.0005
R3087 GND.n476 GND.n474 45.0005
R3088 GND.n476 GND.n475 45.0005
R3089 GND.n486 GND.n477 45.0005
R3090 GND.n845 GND.n477 45.0005
R3091 GND.n860 GND.n859 45.0005
R3092 GND.n1467 GND.n1466 45.0005
R3093 GND.n1466 GND.n1465 45.0005
R3094 GND.n843 GND.n473 45.0005
R3095 GND.n842 GND.n841 45.0005
R3096 GND.n484 GND.n480 45.0005
R3097 GND.n488 GND.n478 45.0005
R3098 GND.n843 GND.n478 45.0005
R3099 GND.n490 GND.n479 45.0005
R3100 GND.n842 GND.n479 45.0005
R3101 GND.n485 GND.n484 45.0005
R3102 GND.n1336 GND.t924 44.7381
R3103 GND.n1334 GND.t923 44.7381
R3104 GND.n1556 GND.t780 44.709
R3105 GND.t955 GND.t794 44.6706
R3106 GND.t142 GND.t554 44.6706
R3107 GND.n1422 GND.t861 44.5993
R3108 GND.t22 GND.t789 44.1861
R3109 GND.n538 GND.n537 43.9358
R3110 GND.t781 GND.t931 43.9247
R3111 GND.t782 GND.t917 43.9247
R3112 GND.n677 GND.n672 43.7886
R3113 GND.n861 GND.n860 43.7516
R3114 GND.t624 GND.n1088 42.9475
R3115 GND.t529 GND.t591 42.8789
R3116 GND.n158 GND.n139 41.7887
R3117 GND.n1701 GND.n29 41.7862
R3118 GND.n1854 GND.n1853 41.7862
R3119 GND.n1853 GND.n1852 41.7862
R3120 GND.n1703 GND.n1602 41.7862
R3121 GND.n1713 GND.n1602 41.7862
R3122 GND.n1857 GND.n1856 41.7862
R3123 GND.n1858 GND.n1857 41.7862
R3124 GND.n1109 GND.n1108 41.7862
R3125 GND.n1110 GND.n1109 41.7862
R3126 GND.n694 GND.n612 41.7076
R3127 GND.n710 GND.n604 39.8486
R3128 GND.n691 GND.n616 39.8486
R3129 GND.n640 GND.n625 39.8486
R3130 GND.n1506 GND.t737 39.7414
R3131 GND.n1549 GND.t52 39.7414
R3132 GND.t613 GND.n221 39.7414
R3133 GND.n1352 GND.t169 39.3159
R3134 GND.n1351 GND.t168 39.3159
R3135 GND.n1350 GND.t899 39.3159
R3136 GND.n1349 GND.t898 39.3159
R3137 GND.n1348 GND.t732 39.3159
R3138 GND.n1347 GND.t731 39.3159
R3139 GND.n1346 GND.t575 39.3159
R3140 GND.n1345 GND.t574 39.3159
R3141 GND.n1343 GND.t480 39.3159
R3142 GND.n1342 GND.t479 39.3159
R3143 GND.n1341 GND.t808 39.3159
R3144 GND.n1340 GND.t807 39.3159
R3145 GND.n1339 GND.t975 39.3159
R3146 GND.n1338 GND.t974 39.3159
R3147 GND.n1388 GND.t970 39.3159
R3148 GND.n1387 GND.t971 39.3159
R3149 GND.n1386 GND.t632 39.3159
R3150 GND.n1385 GND.t633 39.3159
R3151 GND.n1384 GND.t369 39.3159
R3152 GND.n1383 GND.t370 39.3159
R3153 GND.n1382 GND.t411 39.3159
R3154 GND.n1381 GND.t412 39.3159
R3155 GND.n1378 GND.t972 39.3159
R3156 GND.n1377 GND.t973 39.3159
R3157 GND.n1376 GND.t388 39.3159
R3158 GND.n1375 GND.t389 39.3159
R3159 GND.n1374 GND.t709 39.3159
R3160 GND.n1373 GND.t710 39.3159
R3161 GND.n1372 GND.t42 39.3159
R3162 GND.n1371 GND.t43 39.3159
R3163 GND.n197 GND.t776 39.3159
R3164 GND.n580 GND.t775 39.3159
R3165 GND.n579 GND.t659 39.3159
R3166 GND.n198 GND.t658 39.3159
R3167 GND.n1570 GND.t758 39.3159
R3168 GND.n1571 GND.t759 39.3159
R3169 GND.n1573 GND.t566 39.3159
R3170 GND.n1574 GND.t567 39.3159
R3171 GND.n1562 GND.t695 39.3159
R3172 GND.n201 GND.t8 39.3159
R3173 GND.n588 GND.t7 39.3159
R3174 GND.n589 GND.t647 39.3159
R3175 GND.n590 GND.t646 39.3159
R3176 GND.n591 GND.t573 39.3159
R3177 GND.n592 GND.t572 39.3159
R3178 GND.n593 GND.t83 39.3159
R3179 GND.n586 GND.t82 39.3159
R3180 GND.n585 GND.t546 39.3159
R3181 GND.n584 GND.t545 39.3159
R3182 GND.n583 GND.t965 39.3159
R3183 GND.n230 GND.t964 39.3159
R3184 GND.n1519 GND.t423 39.3159
R3185 GND.n1521 GND.t424 39.3159
R3186 GND.n1522 GND.t652 39.3159
R3187 GND.n1524 GND.t653 39.3159
R3188 GND.n1525 GND.t656 39.3159
R3189 GND.n1528 GND.t657 39.3159
R3190 GND.n1529 GND.t921 39.3159
R3191 GND.n1531 GND.t922 39.3159
R3192 GND.n1532 GND.t854 39.3159
R3193 GND.n1533 GND.t855 39.3159
R3194 GND.n202 GND.t694 39.3159
R3195 GND.n1398 GND.t665 39.3159
R3196 GND.n1397 GND.t741 39.3159
R3197 GND.n1396 GND.t742 39.3159
R3198 GND.n333 GND.t714 39.3159
R3199 GND.n358 GND.t713 39.3159
R3200 GND.n359 GND.t761 39.3159
R3201 GND.n360 GND.t760 39.3159
R3202 GND.n361 GND.t739 39.3159
R3203 GND.n362 GND.t738 39.3159
R3204 GND.n363 GND.t933 39.3159
R3205 GND.n357 GND.t932 39.3159
R3206 GND.n356 GND.t967 39.3159
R3207 GND.n355 GND.t966 39.3159
R3208 GND.n354 GND.t536 39.3159
R3209 GND.n353 GND.t535 39.3159
R3210 GND.n352 GND.t363 39.3159
R3211 GND.n351 GND.t362 39.3159
R3212 GND.n350 GND.t730 39.3159
R3213 GND.n349 GND.t729 39.3159
R3214 GND.n347 GND.t751 39.3159
R3215 GND.n346 GND.t752 39.3159
R3216 GND.n345 GND.t442 39.3159
R3217 GND.n344 GND.t443 39.3159
R3218 GND.n343 GND.t676 39.3159
R3219 GND.n342 GND.t677 39.3159
R3220 GND.n341 GND.t648 39.3159
R3221 GND.n340 GND.t649 39.3159
R3222 GND.n339 GND.t762 39.3159
R3223 GND.n337 GND.t763 39.3159
R3224 GND.n336 GND.t962 39.3159
R3225 GND.n320 GND.t963 39.3159
R3226 GND.n1399 GND.t664 39.3159
R3227 GND.n1745 GND.n1731 39.0005
R3228 GND.n1733 GND.n1731 39.0005
R3229 GND.n1738 GND.n1737 39.0005
R3230 GND.n1737 GND.n161 39.0005
R3231 GND.n1712 GND.n1711 39.0005
R3232 GND.n1713 GND.n1712 39.0005
R3233 GND.n1615 GND.n1614 39.0005
R3234 GND.n1614 GND.n1613 39.0005
R3235 GND.n1864 GND.n1863 39.0005
R3236 GND.n1865 GND.n1864 39.0005
R3237 GND.n1758 GND.n1756 39.0005
R3238 GND.n1759 GND.n1758 39.0005
R3239 GND.n1754 GND.n1749 39.0005
R3240 GND.n1754 GND.n20 39.0005
R3241 GND.n1595 GND.n1594 39.0005
R3242 GND.n1590 GND.n187 39.0005
R3243 GND.n1591 GND.n1590 39.0005
R3244 GND.n1774 GND.n1773 39.0005
R3245 GND.n1775 GND.n1774 39.0005
R3246 GND.n1426 GND.n1425 39.0005
R3247 GND.n1425 GND.n1424 39.0005
R3248 GND.n1586 GND.n188 38.777
R3249 GND.t455 GND.n183 38.7342
R3250 GND.t38 GND.t161 38.4342
R3251 GND.n224 GND.t619 38.4342
R3252 GND.t778 GND.n223 38.4342
R3253 GND.n1573 GND.n1572 38.2036
R3254 GND.t138 GND.t105 37.9893
R3255 GND.n1091 GND.t608 37.5791
R3256 GND.n1594 GND.n1593 37.3282
R3257 GND.n1613 GND.t475 37.2444
R3258 GND.t777 GND.t768 36.604
R3259 GND.t784 GND.t681 36.604
R3260 GND.n1596 GND.n185 36.563
R3261 GND.n1807 GND.n1806 36.563
R3262 GND.n1808 GND.n1807 36.563
R3263 GND.n1821 GND.n1820 36.563
R3264 GND.n1433 GND.n1432 36.563
R3265 GND.n1434 GND.n1433 36.563
R3266 GND GND.t912 36.2742
R3267 GND.t913 GND 36.2742
R3268 GND.t394 GND 36.2742
R3269 GND.n1058 GND.n1056 36.1417
R3270 GND.n1059 GND.n1058 36.1417
R3271 GND.n1067 GND.n1065 36.1417
R3272 GND.n1068 GND.n1067 36.1417
R3273 GND.n1076 GND.n1074 36.1417
R3274 GND.n1077 GND.n1076 36.1417
R3275 GND.n1083 GND.n1043 36.1417
R3276 GND.n1093 GND.n1043 36.1417
R3277 GND.n1039 GND.n865 36.1417
R3278 GND.n1035 GND.n865 36.1417
R3279 GND.n1035 GND.n1034 36.1417
R3280 GND.n1034 GND.n1033 36.1417
R3281 GND.n1033 GND.n875 36.1417
R3282 GND.n1027 GND.n1026 36.1417
R3283 GND.n1026 GND.n1025 36.1417
R3284 GND.n1025 GND.n886 36.1417
R3285 GND.n1019 GND.n886 36.1417
R3286 GND.n1019 GND.n1018 36.1417
R3287 GND.n1013 GND.n897 36.1417
R3288 GND.n1007 GND.n897 36.1417
R3289 GND.n1007 GND.n1006 36.1417
R3290 GND.n1006 GND.n1005 36.1417
R3291 GND.n1005 GND.n907 36.1417
R3292 GND.n999 GND.n998 36.1417
R3293 GND.n998 GND.n997 36.1417
R3294 GND.n997 GND.n918 36.1417
R3295 GND.n991 GND.n918 36.1417
R3296 GND.n991 GND.n990 36.1417
R3297 GND.n985 GND.n929 36.1417
R3298 GND.n979 GND.n929 36.1417
R3299 GND.n979 GND.n978 36.1417
R3300 GND.n978 GND.n977 36.1417
R3301 GND.n977 GND.n939 36.1417
R3302 GND.n971 GND.n970 36.1417
R3303 GND.n970 GND.n969 36.1417
R3304 GND.n969 GND.n950 36.1417
R3305 GND.n963 GND.n950 36.1417
R3306 GND.n963 GND.n962 36.1417
R3307 GND.n1212 GND.n1211 36.1417
R3308 GND.n1211 GND.n1210 36.1417
R3309 GND.n1210 GND.n398 36.1417
R3310 GND.n1204 GND.n398 36.1417
R3311 GND.n1204 GND.n1203 36.1417
R3312 GND.n1198 GND.n409 36.1417
R3313 GND.n1192 GND.n409 36.1417
R3314 GND.n1187 GND.n414 36.1417
R3315 GND.n1150 GND.n414 36.1417
R3316 GND.n1179 GND.n1178 36.1417
R3317 GND.n1178 GND.n1177 36.1417
R3318 GND.n1172 GND.n1160 36.1417
R3319 GND.n1165 GND.n1160 36.1417
R3320 GND.t628 GND.n1090 36.1338
R3321 GND.t929 GND.t597 36.1338
R3322 GND.t704 GND.t60 35.8196
R3323 GND.t784 GND.t768 35.5582
R3324 GND.t681 GND.t781 35.5582
R3325 GND.n1336 GND.t409 35.1381
R3326 GND.n1334 GND.t408 35.1381
R3327 GND.n1593 GND.n185 34.9952
R3328 GND.n1223 GND.n385 34.6358
R3329 GND.n1227 GND.n1226 34.6358
R3330 GND.n1229 GND.n1227 34.6358
R3331 GND.n1263 GND.n1262 34.6358
R3332 GND.n1309 GND.n1306 34.6358
R3333 GND.n537 GND.n493 34.6358
R3334 GND.n533 GND.n493 34.6358
R3335 GND.n533 GND.n532 34.6358
R3336 GND.n532 GND.n531 34.6358
R3337 GND.n531 GND.n495 34.6358
R3338 GND.n526 GND.n496 34.6358
R3339 GND.n522 GND.n521 34.6358
R3340 GND.n521 GND.n498 34.6358
R3341 GND.n517 GND.n498 34.6358
R3342 GND.n514 GND.n502 34.6358
R3343 GND.n509 GND.n503 34.6358
R3344 GND.n627 GND.n608 34.6358
R3345 GND.n718 GND.n717 34.6358
R3346 GND.n708 GND.n606 34.6358
R3347 GND.n715 GND.n602 34.6358
R3348 GND.n642 GND.n622 34.6358
R3349 GND.n689 GND.n618 34.6358
R3350 GND.n654 GND.n653 34.6358
R3351 GND.n658 GND.n621 34.6358
R3352 GND.n636 GND.n634 34.6358
R3353 GND.t396 GND.t625 33.8625
R3354 GND.t163 GND.t38 33.728
R3355 GND.n224 GND.t901 33.728
R3356 GND.n223 GND.t788 33.728
R3357 GND.t410 GND.t795 33.717
R3358 GND.n687 GND.n619 33.5688
R3359 GND.n631 GND.n628 33.5688
R3360 GND.n706 GND.n607 33.5688
R3361 GND.n600 GND.n599 33.5688
R3362 GND.n651 GND.n650 33.5688
R3363 GND.n644 GND.n623 33.5688
R3364 GND.n1309 GND.n1308 32.7534
R3365 GND.n1445 GND.t515 32.6237
R3366 GND.n1427 GND.n300 32.5005
R3367 GND.n1126 GND.n300 32.5005
R3368 GND.n1598 GND.n1597 30.79
R3369 GND.n1599 GND.n1598 30.79
R3370 GND.n613 GND.n611 30.79
R3371 GND.n667 GND.n611 30.79
R3372 GND.n696 GND.n695 30.79
R3373 GND.n697 GND.n696 30.79
R3374 GND.n664 GND.n612 30.79
R3375 GND.n1447 GND.n1446 30.79
R3376 GND.n1446 GND.n1445 30.79
R3377 GND.n1829 GND.n139 30.1181
R3378 GND.n157 GND.n140 30.1181
R3379 GND.t928 GND.t458 29.9395
R3380 GND.n326 GND.n246 29.3652
R3381 GND.t786 GND.t529 29.2833
R3382 GND.t591 GND.t613 29.2833
R3383 GND.t73 GND.t89 29.0508
R3384 GND.t20 GND 29.0195
R3385 GND.t902 GND 29.0195
R3386 GND GND.t945 29.0195
R3387 GND.n1136 GND.n255 28.9887
R3388 GND.n1489 GND.n1488 28.9887
R3389 GND.n1089 GND.t624 28.4942
R3390 GND.n1140 GND.t771 28.4942
R3391 GND.t931 GND.t782 28.2375
R3392 GND.t917 GND.t787 28.2375
R3393 GND.n1618 GND.n17 27.8576
R3394 GND.n1713 GND.n17 27.8576
R3395 GND.n1859 GND.n19 27.8576
R3396 GND.n1859 GND.n1858 27.8576
R3397 GND.n159 GND.n158 27.8576
R3398 GND.n159 GND.n134 27.8576
R3399 GND.n1810 GND.n160 27.8576
R3400 GND.n1810 GND.n1809 27.8576
R3401 GND.n154 GND.n152 27.8576
R3402 GND.n1819 GND.n152 27.8576
R3403 GND.n1813 GND.n1812 27.8576
R3404 GND.n1812 GND.n134 27.8576
R3405 GND.n1777 GND.n156 27.8576
R3406 GND.n1809 GND.n156 27.8576
R3407 GND.n1816 GND.n1815 27.8576
R3408 GND.n1819 GND.n1816 27.8576
R3409 GND.t787 GND.n1556 27.4531
R3410 GND.t958 GND.n843 26.6966
R3411 GND.n843 GND.t520 26.6966
R3412 GND.t753 GND.n842 26.6966
R3413 GND.n842 GND.t809 26.6966
R3414 GND.n484 GND.t581 26.6966
R3415 GND.n484 GND.t725 26.6966
R3416 GND.n1714 GND.n182 26.5914
R3417 GND.n1714 GND.n1713 26.5914
R3418 GND.n179 GND.n21 26.5914
R3419 GND.n1858 GND.n21 26.5914
R3420 GND.n277 GND.n276 26.5914
R3421 GND.t45 GND.n277 26.5914
R3422 GND.t493 GND.t860 26.2229
R3423 GND.t12 GND.t403 26.1458
R3424 GND.n1262 GND.n1261 25.977
R3425 GND.n527 GND.n495 25.977
R3426 GND.n517 GND.n516 25.977
R3427 GND.n1473 GND.n1472 25.4353
R3428 GND.n1474 GND.n1473 25.4353
R3429 GND.t791 GND.n193 25.3615
R3430 GND.n727 GND.n577 25.224
R3431 GND.n731 GND.n577 25.224
R3432 GND.n733 GND.n732 25.224
R3433 GND.n733 GND.n574 25.224
R3434 GND.n738 GND.n573 25.224
R3435 GND.n742 GND.n573 25.224
R3436 GND.n744 GND.n743 25.224
R3437 GND.n744 GND.n570 25.224
R3438 GND.n749 GND.n569 25.224
R3439 GND.n753 GND.n569 25.224
R3440 GND.n755 GND.n754 25.224
R3441 GND.n755 GND.n566 25.224
R3442 GND.n760 GND.n565 25.224
R3443 GND.n764 GND.n565 25.224
R3444 GND.n766 GND.n765 25.224
R3445 GND.n766 GND.n562 25.224
R3446 GND.n771 GND.n561 25.224
R3447 GND.n775 GND.n561 25.224
R3448 GND.n777 GND.n776 25.224
R3449 GND.n777 GND.n558 25.224
R3450 GND.n782 GND.n557 25.224
R3451 GND.n786 GND.n557 25.224
R3452 GND.n788 GND.n787 25.224
R3453 GND.n788 GND.n554 25.224
R3454 GND.n793 GND.n553 25.224
R3455 GND.n797 GND.n553 25.224
R3456 GND.n799 GND.n798 25.224
R3457 GND.n799 GND.n550 25.224
R3458 GND.n804 GND.n549 25.224
R3459 GND.n808 GND.n549 25.224
R3460 GND.n810 GND.n809 25.224
R3461 GND.n810 GND.n546 25.224
R3462 GND.n815 GND.n545 25.224
R3463 GND.n819 GND.n545 25.224
R3464 GND.n821 GND.n820 25.224
R3465 GND.n821 GND.n542 25.224
R3466 GND.n827 GND.n826 25.224
R3467 GND.n827 GND.n540 25.224
R3468 GND.n832 GND.n831 25.224
R3469 GND.n833 GND.n832 25.224
R3470 GND.n839 GND.n492 25.1797
R3471 GND.n840 GND.n481 25.1797
R3472 GND.n483 GND.n482 25.1797
R3473 GND.n847 GND.n472 25.1797
R3474 GND.n848 GND.n470 25.1797
R3475 GND.n849 GND.n462 25.1797
R3476 GND.n464 GND.n463 25.1797
R3477 GND.n855 GND.n455 25.1797
R3478 GND.n454 GND.n453 25.1797
R3479 GND.n675 GND.n674 25.1797
R3480 GND.n676 GND.n673 25.1797
R3481 GND.n1549 GND.t111 25.1
R3482 GND.n610 GND.t407 25.0567
R3483 GND.t416 GND.t417 24.5815
R3484 GND.n1299 GND.n1298 24.4711
R3485 GND.n1298 GND.n1297 24.4711
R3486 GND.n1276 GND.n1275 24.4711
R3487 GND.n164 GND.n162 24.3755
R3488 GND.n1734 GND.n162 24.3755
R3489 GND.n1772 GND.n163 24.3755
R3490 GND.n1734 GND.n163 24.3755
R3491 GND.n1766 GND.n1765 24.3755
R3492 GND.n1767 GND.n1766 24.3755
R3493 GND.n1762 GND.n1761 24.3755
R3494 GND.n1761 GND.n1760 24.3755
R3495 GND.n1608 GND.n1607 24.3755
R3496 GND.n1608 GND.n9 24.3755
R3497 GND.n1605 GND.n1603 24.3755
R3498 GND.n1612 GND.n1603 24.3755
R3499 GND.n1769 GND.n1768 24.3755
R3500 GND.n1768 GND.n1767 24.3755
R3501 GND.n1757 GND.n16 24.3755
R3502 GND.n1760 GND.n1757 24.3755
R3503 GND.n1610 GND.n14 24.3755
R3504 GND.n1610 GND.n9 24.3755
R3505 GND.n1617 GND.n1604 24.3755
R3506 GND.n1612 GND.n1604 24.3755
R3507 GND.t627 GND.t968 24.3646
R3508 GND.n582 GND 24.3288
R3509 GND.n1263 GND.n1218 24.0946
R3510 GND.n527 GND.n526 24.0946
R3511 GND.n1248 GND.n1238 23.7181
R3512 GND.n1250 GND.n1235 23.7181
R3513 GND.n1270 GND.n385 23.7181
R3514 GND.n1267 GND.n1219 23.7181
R3515 GND.n1306 GND.n1305 23.7181
R3516 GND.n1314 GND.n370 23.7181
R3517 GND.n1304 GND.n373 23.7181
R3518 GND.n1294 GND.n1293 23.7181
R3519 GND.n1285 GND.n1284 23.7181
R3520 GND.n515 GND.n514 23.7181
R3521 GND.n510 GND.n509 23.7181
R3522 GND.n699 GND.n608 23.7181
R3523 GND.n718 GND.n597 23.7181
R3524 GND.n709 GND.n708 23.7181
R3525 GND.n716 GND.n715 23.7181
R3526 GND.n642 GND.n641 23.7181
R3527 GND.n690 GND.n689 23.7181
R3528 GND.n657 GND.n654 23.7181
R3529 GND.n662 GND.n621 23.7181
R3530 GND.n634 GND.n633 23.7181
R3531 GND.n1278 GND.n380 23.3417
R3532 GND.n1087 GND.t459 23.1258
R3533 GND.t916 GND.n416 22.7128
R3534 GND.n1464 GND.t685 22.5064
R3535 GND.n1244 GND.n1238 22.2123
R3536 GND.n1250 GND.n1249 22.2123
R3537 GND.n1305 GND.n1304 22.2123
R3538 GND.n1289 GND.n1288 22.2123
R3539 GND.n510 GND.n502 22.2123
R3540 GND.n505 GND.n503 22.2123
R3541 GND.n633 GND.n627 22.2123
R3542 GND.n717 GND.n716 22.2123
R3543 GND.n703 GND.n606 22.2123
R3544 GND.n710 GND.n709 22.2123
R3545 GND.n603 GND.n602 22.2123
R3546 GND.n647 GND.n622 22.2123
R3547 GND.n684 GND.n618 22.2123
R3548 GND.n691 GND.n690 22.2123
R3549 GND.n653 GND.n652 22.2123
R3550 GND.n658 GND.n657 22.2123
R3551 GND.n641 GND.n640 22.2123
R3552 GND.n636 GND.n635 22.2123
R3553 GND.t618 GND.t112 21.9626
R3554 GND.t901 GND.t703 21.9626
R3555 GND.t788 GND.t519 21.9626
R3556 GND.t789 GND.t914 21.9626
R3557 GND.t60 GND.t631 21.7011
R3558 GND.n613 GND 21.0039
R3559 GND.n1858 GND.n20 20.8571
R3560 GND.n1090 GND.t622 20.8546
R3561 GND.t459 GND.t930 20.8546
R3562 GND.t513 GND.t626 20.8546
R3563 GND.t597 GND.t145 20.8546
R3564 GND.t625 GND.t526 20.8546
R3565 GND.n699 GND 20.7453
R3566 GND GND.n597 20.7453
R3567 GND.n702 GND 20.7453
R3568 GND.n648 GND 20.7453
R3569 GND GND.n662 20.7453
R3570 GND.n683 GND 20.7453
R3571 GND.n732 GND.n731 20.3299
R3572 GND.n743 GND.n742 20.3299
R3573 GND.n754 GND.n753 20.3299
R3574 GND.n765 GND.n764 20.3299
R3575 GND.n776 GND.n775 20.3299
R3576 GND.n787 GND.n786 20.3299
R3577 GND.n798 GND.n797 20.3299
R3578 GND.n809 GND.n808 20.3299
R3579 GND.n820 GND.n819 20.3299
R3580 GND.n831 GND.n540 20.3299
R3581 GND.n1300 GND.n1299 19.9534
R3582 GND.n1434 GND.n231 19.8222
R3583 GND.n1110 GND.t623 19.4092
R3584 GND.t596 GND.n435 19.2028
R3585 GND.n1277 GND.n1276 19.2005
R3586 GND.n1414 GND.n1413 18.2817
R3587 GND.n1415 GND.n1414 18.2817
R3588 GND.n1417 GND.n1416 18.2817
R3589 GND.n1416 GND.n1415 18.2817
R3590 GND.n315 GND.n314 18.2817
R3591 GND.n1406 GND.n315 18.2817
R3592 GND.n1401 GND.n316 18.2817
R3593 GND.n1406 GND.n316 18.2817
R3594 GND.n328 GND.n327 18.2817
R3595 GND.n329 GND.n328 18.2817
R3596 GND.n331 GND.n330 18.2817
R3597 GND.n330 GND.n329 18.2817
R3598 GND.n1483 GND.n1482 18.2817
R3599 GND.n1484 GND.n1483 18.2817
R3600 GND.n1486 GND.n1485 18.2817
R3601 GND.n1485 GND.n1484 18.2817
R3602 GND.n1491 GND.n1490 18.2817
R3603 GND.n1492 GND.n1491 18.2817
R3604 GND.n1501 GND.n1500 18.2817
R3605 GND.n1502 GND.n1501 18.2817
R3606 GND.n1494 GND.n1493 18.2817
R3607 GND.n1493 GND.n1492 18.2817
R3608 GND.n1497 GND.n242 18.2817
R3609 GND.n1502 GND.n242 18.2817
R3610 GND.n422 GND.n301 18.2817
R3611 GND.n1113 GND.n301 18.2817
R3612 GND.n304 GND.n302 18.2817
R3613 GND.n1113 GND.n302 18.2817
R3614 GND.n419 GND.n417 18.2817
R3615 GND.n1089 GND.n417 18.2817
R3616 GND.n1145 GND.n418 18.2817
R3617 GND.n1089 GND.n418 18.2817
R3618 GND.n1139 GND.n1138 18.2817
R3619 GND.n1140 GND.n1139 18.2817
R3620 GND.n1142 GND.n1141 18.2817
R3621 GND.n1141 GND.n1140 18.2817
R3622 GND.n1477 GND.n1476 18.2817
R3623 GND.n1476 GND.n1475 18.2817
R3624 GND.n1128 GND.n268 18.2817
R3625 GND.n1475 GND.n268 18.2817
R3626 GND.t915 GND.t81 18.1704
R3627 GND.n727 GND.n726 17.3181
R3628 GND.n738 GND.n737 17.3181
R3629 GND.n749 GND.n748 17.3181
R3630 GND.n760 GND.n759 17.3181
R3631 GND.n771 GND.n770 17.3181
R3632 GND.n782 GND.n781 17.3181
R3633 GND.n793 GND.n792 17.3181
R3634 GND.n804 GND.n803 17.3181
R3635 GND.n815 GND.n814 17.3181
R3636 GND.n826 GND.n825 17.3181
R3637 GND.t619 GND.t785 17.2564
R3638 GND.t900 GND.t790 17.2564
R3639 GND.t84 GND.t778 17.2564
R3640 GND.t6 GND.t792 17.2564
R3641 GND.n1543 GND.n208 17.2064
R3642 GND.n221 GND.n208 17.2064
R3643 GND.n1553 GND.n209 17.2064
R3644 GND.n221 GND.n209 17.2064
R3645 GND.n1115 GND.n1114 17.2064
R3646 GND.n1114 GND.t396 17.2064
R3647 GND.t419 GND.n1759 16.3878
R3648 GND.n1510 GND.n1506 15.9492
R3649 GND.n737 GND.n574 15.8123
R3650 GND.n748 GND.n570 15.8123
R3651 GND.n759 GND.n566 15.8123
R3652 GND.n770 GND.n562 15.8123
R3653 GND.n781 GND.n558 15.8123
R3654 GND.n792 GND.n554 15.8123
R3655 GND.n803 GND.n550 15.8123
R3656 GND.n814 GND.n546 15.8123
R3657 GND.n825 GND.n542 15.8123
R3658 GND.n151 GND.n149 15.8113
R3659 GND.n151 GND.n134 15.8113
R3660 GND.n307 GND.t767 15.4862
R3661 GND.n1261 GND.n1233 15.4358
R3662 GND.n1279 GND.n1277 15.4358
R3663 GND.n1344 GND.n1343 15.0979
R3664 GND.n297 GND.n295 15.0005
R3665 GND.t968 GND.n295 15.0005
R3666 GND.t148 GND.n844 14.708
R3667 GND.t918 GND.t107 14.6603
R3668 GND.t630 GND.t111 14.6419
R3669 GND.t534 GND.t706 14.6419
R3670 GND.t631 GND.t113 14.6419
R3671 GND.t683 GND.t704 14.6419
R3672 GND.t533 GND.t402 14.6419
R3673 GND.t375 GND.t911 14.51
R3674 GND.t551 GND.t400 14.51
R3675 GND.t395 GND.t155 14.51
R3676 GND.t393 GND.t493 14.2473
R3677 GND.n1088 GND.t621 14.0409
R3678 GND.t458 GND.n1105 14.0409
R3679 GND.t859 GND.t391 14.0409
R3680 GND.t95 GND.n1832 13.9614
R3681 GND.n1434 GND.t391 13.8344
R3682 GND.n1381 GND.n1380 13.7851
R3683 GND.n1275 GND.n1274 13.5534
R3684 GND.n1564 GND.n1563 13.296
R3685 GND.n1565 GND.n1564 13.296
R3686 GND.n1576 GND.n1575 13.296
R3687 GND.n1577 GND.n1576 13.296
R3688 GND.n1569 GND.n1568 13.296
R3689 GND.n1568 GND.n1567 13.296
R3690 GND.n1394 GND.n1393 13.296
R3691 GND.n1393 GND.n1392 13.296
R3692 GND.n1370 GND.n1369 13.296
R3693 GND.n1369 GND.n1368 13.296
R3694 GND.n1390 GND.n1389 13.296
R3695 GND.n1391 GND.n1390 13.296
R3696 GND.n1518 GND.n1517 13.296
R3697 GND.n1517 GND.n1516 13.296
R3698 GND.n348 GND.n335 13.296
R3699 GND.n1045 GND.n335 13.296
R3700 GND.n1113 GND.t45 13.215
R3701 GND.n1257 GND.n1233 13.177
R3702 GND.n1300 GND.n373 13.177
R3703 GND.n516 GND.n515 13.177
R3704 GND.n681 GND.n596 13.0995
R3705 GND.n721 GND.n720 13.0995
R3706 GND.n1424 GND.t918 12.802
R3707 GND.n1243 GND.n1239 12.8005
R3708 GND.n1254 GND.n1234 12.8005
R3709 GND.n1289 GND.n377 12.8005
R3710 GND.n1283 GND.n380 12.8005
R3711 GND.n1320 GND.n366 12.8005
R3712 GND.n505 GND.n366 12.8005
R3713 GND.n703 GND.n702 12.8005
R3714 GND.n648 GND.n647 12.8005
R3715 GND.n684 GND.n683 12.8005
R3716 GND.n1463 GND.n1462 12.4473
R3717 GND.n1464 GND.n1463 12.4473
R3718 GND.n1120 GND.t627 12.389
R3719 GND.n1482 GND.n1481 12.0476
R3720 GND.n1325 GND.t772 11.8635
R3721 GND.n1833 GND.t660 11.6346
R3722 GND.n1578 GND.n134 11.6346
R3723 GND.n1045 GND.t916 11.3567
R3724 GND.n1244 GND.n1243 11.2946
R3725 GND.n1249 GND.n1248 11.2946
R3726 GND.n1254 GND.n1235 11.2946
R3727 GND.n1257 GND.n1234 11.2946
R3728 GND.n1293 GND.n377 11.2946
R3729 GND.n1284 GND.n1283 11.2946
R3730 GND.n1462 GND.n1461 11.2946
R3731 GND.n1472 GND.n1471 11.2946
R3732 GND.n1448 GND.n1447 11.2946
R3733 GND.n695 GND.n614 10.9181
R3734 GND.t686 GND.t110 10.7372
R3735 GND.n1223 GND.n1221 10.5417
R3736 GND.n1229 GND.n1228 10.5417
R3737 GND.n1294 GND.n376 10.5417
R3738 GND.n1285 GND.n378 10.5417
R3739 GND.n497 GND.n496 10.5417
R3740 GND.n1110 GND.t513 10.5308
R3741 GND.n1454 GND.t861 10.5308
R3742 GND.n1865 GND.n10 10.4288
R3743 GND.n1792 GND.t249 10.3318
R3744 GND.n1792 GND.t99 10.3318
R3745 GND.n1793 GND.t427 10.3318
R3746 GND.n1793 GND.t428 10.3318
R3747 GND.n1794 GND.t92 10.3318
R3748 GND.n1794 GND.t102 10.3318
R3749 GND.n1795 GND.t804 10.3318
R3750 GND.n1795 GND.t251 10.3318
R3751 GND.n1782 GND.t806 10.3318
R3752 GND.n1782 GND.t233 10.3318
R3753 GND.n1781 GND.t97 10.3318
R3754 GND.n1781 GND.t805 10.3318
R3755 GND.n1780 GND.t94 10.3318
R3756 GND.n1780 GND.t96 10.3318
R3757 GND.n1779 GND.t230 10.3318
R3758 GND.n1779 GND.t100 10.3318
R3759 GND.t81 GND.n1089 10.3243
R3760 GND.n1424 GND.n1423 10.3243
R3761 GND.n1329 GND.n357 10.1749
R3762 GND.n1785 GND.n134 10.0867
R3763 GND.n1786 GND.n1785 10.0867
R3764 GND GND.n614 10.0862
R3765 GND.n694 GND 10.0862
R3766 GND.n432 GND.n426 9.91575
R3767 GND.n428 GND.n426 9.91575
R3768 GND.n429 GND.n427 9.91575
R3769 GND.n429 GND.n428 9.91575
R3770 GND.n1056 GND.n1055 9.32838
R3771 GND.n720 GND.n597 9.3031
R3772 GND.n1096 GND.n447 9.3005
R3773 GND.n717 GND.n598 9.3005
R3774 GND.n719 GND.n718 9.3005
R3775 GND.n716 GND.n601 9.3005
R3776 GND.n713 GND.n602 9.3005
R3777 GND.n715 GND.n714 9.3005
R3778 GND.n700 GND.n699 9.3005
R3779 GND.n630 GND.n627 9.3005
R3780 GND.n629 GND.n608 9.3005
R3781 GND.n709 GND.n605 9.3005
R3782 GND.n704 GND.n703 9.3005
R3783 GND.n702 GND.n701 9.3005
R3784 GND.n705 GND.n606 9.3005
R3785 GND.n708 GND.n707 9.3005
R3786 GND.n711 GND.n710 9.3005
R3787 GND.n633 GND.n632 9.3005
R3788 GND.n662 GND.n661 9.3005
R3789 GND.n657 GND.n656 9.3005
R3790 GND.n653 GND.n615 9.3005
R3791 GND.n655 GND.n654 9.3005
R3792 GND.n659 GND.n658 9.3005
R3793 GND.n660 GND.n621 9.3005
R3794 GND.n647 GND.n646 9.3005
R3795 GND.n649 GND.n648 9.3005
R3796 GND.n645 GND.n622 9.3005
R3797 GND.n643 GND.n642 9.3005
R3798 GND.n641 GND.n624 9.3005
R3799 GND.n640 GND.n639 9.3005
R3800 GND.n637 GND.n636 9.3005
R3801 GND.n634 GND.n626 9.3005
R3802 GND.n690 GND.n617 9.3005
R3803 GND.n685 GND.n684 9.3005
R3804 GND.n686 GND.n618 9.3005
R3805 GND.n689 GND.n688 9.3005
R3806 GND.n692 GND.n691 9.3005
R3807 GND.n683 GND.n682 9.3005
R3808 GND.n1080 GND.n1079 9.3005
R3809 GND.n1081 GND.n1080 9.3005
R3810 GND.n1071 GND.n1070 9.3005
R3811 GND.n1072 GND.n1071 9.3005
R3812 GND.n1062 GND.n1061 9.3005
R3813 GND.n1063 GND.n1062 9.3005
R3814 GND.n1094 GND.n1093 9.3005
R3815 GND.n1043 GND.n1042 9.3005
R3816 GND.n1083 GND.n1082 9.3005
R3817 GND.n1078 GND.n1077 9.3005
R3818 GND.n1076 GND.n1052 9.3005
R3819 GND.n1074 GND.n1073 9.3005
R3820 GND.n1069 GND.n1068 9.3005
R3821 GND.n1067 GND.n1053 9.3005
R3822 GND.n1065 GND.n1064 9.3005
R3823 GND.n1060 GND.n1059 9.3005
R3824 GND.n1058 GND.n1054 9.3005
R3825 GND.n1162 GND.n1161 9.3005
R3826 GND.n1163 GND.n1162 9.3005
R3827 GND.n1174 GND.n1158 9.3005
R3828 GND.n1175 GND.n1174 9.3005
R3829 GND.n1153 GND.n1152 9.3005
R3830 GND.n1154 GND.n1153 9.3005
R3831 GND.n1189 GND.n412 9.3005
R3832 GND.n1190 GND.n1189 9.3005
R3833 GND.n1200 GND.n407 9.3005
R3834 GND.n1201 GND.n1200 9.3005
R3835 GND.n403 GND.n402 9.3005
R3836 GND.n404 GND.n403 9.3005
R3837 GND.n959 GND.n958 9.3005
R3838 GND.n960 GND.n959 9.3005
R3839 GND.n954 GND.n953 9.3005
R3840 GND.n955 GND.n954 9.3005
R3841 GND.n945 GND.n944 9.3005
R3842 GND.n946 GND.n945 9.3005
R3843 GND.n935 GND.n934 9.3005
R3844 GND.n936 GND.n935 9.3005
R3845 GND.n987 GND.n927 9.3005
R3846 GND.n988 GND.n987 9.3005
R3847 GND.n923 GND.n922 9.3005
R3848 GND.n924 GND.n923 9.3005
R3849 GND.n913 GND.n912 9.3005
R3850 GND.n914 GND.n913 9.3005
R3851 GND.n903 GND.n902 9.3005
R3852 GND.n904 GND.n903 9.3005
R3853 GND.n1015 GND.n895 9.3005
R3854 GND.n1016 GND.n1015 9.3005
R3855 GND.n891 GND.n890 9.3005
R3856 GND.n892 GND.n891 9.3005
R3857 GND.n881 GND.n880 9.3005
R3858 GND.n882 GND.n881 9.3005
R3859 GND.n871 GND.n870 9.3005
R3860 GND.n872 GND.n871 9.3005
R3861 GND.n1165 GND.n1164 9.3005
R3862 GND.n1160 GND.n1159 9.3005
R3863 GND.n1173 GND.n1172 9.3005
R3864 GND.n1177 GND.n1176 9.3005
R3865 GND.n1178 GND.n1156 9.3005
R3866 GND.n1179 GND.n1155 9.3005
R3867 GND.n1151 GND.n1150 9.3005
R3868 GND.n414 GND.n413 9.3005
R3869 GND.n1188 GND.n1187 9.3005
R3870 GND.n1192 GND.n1191 9.3005
R3871 GND.n409 GND.n408 9.3005
R3872 GND.n1199 GND.n1198 9.3005
R3873 GND.n1203 GND.n1202 9.3005
R3874 GND.n1204 GND.n406 9.3005
R3875 GND.n405 GND.n398 9.3005
R3876 GND.n1210 GND.n397 9.3005
R3877 GND.n1211 GND.n396 9.3005
R3878 GND.n1212 GND.n395 9.3005
R3879 GND.n962 GND.n961 9.3005
R3880 GND.n963 GND.n957 9.3005
R3881 GND.n956 GND.n950 9.3005
R3882 GND.n969 GND.n949 9.3005
R3883 GND.n970 GND.n948 9.3005
R3884 GND.n971 GND.n947 9.3005
R3885 GND.n943 GND.n939 9.3005
R3886 GND.n977 GND.n938 9.3005
R3887 GND.n978 GND.n937 9.3005
R3888 GND.n979 GND.n933 9.3005
R3889 GND.n929 GND.n928 9.3005
R3890 GND.n986 GND.n985 9.3005
R3891 GND.n990 GND.n989 9.3005
R3892 GND.n991 GND.n926 9.3005
R3893 GND.n925 GND.n918 9.3005
R3894 GND.n997 GND.n917 9.3005
R3895 GND.n998 GND.n916 9.3005
R3896 GND.n999 GND.n915 9.3005
R3897 GND.n911 GND.n907 9.3005
R3898 GND.n1005 GND.n906 9.3005
R3899 GND.n1006 GND.n905 9.3005
R3900 GND.n1007 GND.n901 9.3005
R3901 GND.n897 GND.n896 9.3005
R3902 GND.n1014 GND.n1013 9.3005
R3903 GND.n1018 GND.n1017 9.3005
R3904 GND.n1019 GND.n894 9.3005
R3905 GND.n893 GND.n886 9.3005
R3906 GND.n1025 GND.n885 9.3005
R3907 GND.n1026 GND.n884 9.3005
R3908 GND.n1027 GND.n883 9.3005
R3909 GND.n879 GND.n875 9.3005
R3910 GND.n1033 GND.n874 9.3005
R3911 GND.n1034 GND.n873 9.3005
R3912 GND.n1035 GND.n869 9.3005
R3913 GND.n865 GND.n864 9.3005
R3914 GND.n1040 GND.n1039 9.3005
R3915 GND.n504 GND.n366 9.3005
R3916 GND.n506 GND.n505 9.3005
R3917 GND.n507 GND.n503 9.3005
R3918 GND.n509 GND.n508 9.3005
R3919 GND.n511 GND.n510 9.3005
R3920 GND.n512 GND.n502 9.3005
R3921 GND.n514 GND.n513 9.3005
R3922 GND.n515 GND.n500 9.3005
R3923 GND.n516 GND.n499 9.3005
R3924 GND.n518 GND.n517 9.3005
R3925 GND.n519 GND.n498 9.3005
R3926 GND.n521 GND.n520 9.3005
R3927 GND.n523 GND.n522 9.3005
R3928 GND.n524 GND.n496 9.3005
R3929 GND.n526 GND.n525 9.3005
R3930 GND.n528 GND.n527 9.3005
R3931 GND.n529 GND.n495 9.3005
R3932 GND.n531 GND.n530 9.3005
R3933 GND.n532 GND.n494 9.3005
R3934 GND.n534 GND.n533 9.3005
R3935 GND.n535 GND.n493 9.3005
R3936 GND.n537 GND.n536 9.3005
R3937 GND.n1321 GND.n1320 9.3005
R3938 GND.n1274 GND.n1273 9.3005
R3939 GND.n1281 GND.n380 9.3005
R3940 GND.n1283 GND.n1282 9.3005
R3941 GND.n1293 GND.n1292 9.3005
R3942 GND.n1301 GND.n1300 9.3005
R3943 GND.n1302 GND.n373 9.3005
R3944 GND.n1311 GND.n370 9.3005
R3945 GND.n1314 GND.n1313 9.3005
R3946 GND.n1310 GND.n1309 9.3005
R3947 GND.n1306 GND.n371 9.3005
R3948 GND.n1305 GND.n372 9.3005
R3949 GND.n1304 GND.n1303 9.3005
R3950 GND.n1299 GND.n374 9.3005
R3951 GND.n1298 GND.n375 9.3005
R3952 GND.n1297 GND.n1296 9.3005
R3953 GND.n1295 GND.n1294 9.3005
R3954 GND.n1291 GND.n377 9.3005
R3955 GND.n1290 GND.n1289 9.3005
R3956 GND.n1288 GND.n1287 9.3005
R3957 GND.n1286 GND.n1285 9.3005
R3958 GND.n1284 GND.n379 9.3005
R3959 GND.n1280 GND.n1279 9.3005
R3960 GND.n1276 GND.n382 9.3005
R3961 GND.n1275 GND.n383 9.3005
R3962 GND.n1267 GND.n1266 9.3005
R3963 GND.n1261 GND.n1260 9.3005
R3964 GND.n1236 GND.n1234 9.3005
R3965 GND.n1254 GND.n1253 9.3005
R3966 GND.n1249 GND.n1237 9.3005
R3967 GND.n1245 GND.n1244 9.3005
R3968 GND.n1243 GND.n1242 9.3005
R3969 GND.n1241 GND.n1239 9.3005
R3970 GND.n1246 GND.n1238 9.3005
R3971 GND.n1248 GND.n1247 9.3005
R3972 GND.n1251 GND.n1250 9.3005
R3973 GND.n1252 GND.n1235 9.3005
R3974 GND.n1258 GND.n1257 9.3005
R3975 GND.n1259 GND.n1233 9.3005
R3976 GND.n1262 GND.n1232 9.3005
R3977 GND.n1264 GND.n1263 9.3005
R3978 GND.n1265 GND.n1218 9.3005
R3979 GND.n1231 GND.n1219 9.3005
R3980 GND.n1230 GND.n1229 9.3005
R3981 GND.n1227 GND.n1220 9.3005
R3982 GND.n1226 GND.n1225 9.3005
R3983 GND.n1224 GND.n1223 9.3005
R3984 GND.n1222 GND.n385 9.3005
R3985 GND.n1271 GND.n1270 9.3005
R3986 GND.n834 GND.n833 9.3005
R3987 GND.n832 GND.n539 9.3005
R3988 GND.n831 GND.n830 9.3005
R3989 GND.n829 GND.n540 9.3005
R3990 GND.n828 GND.n827 9.3005
R3991 GND.n826 GND.n541 9.3005
R3992 GND.n825 GND.n824 9.3005
R3993 GND.n823 GND.n542 9.3005
R3994 GND.n822 GND.n821 9.3005
R3995 GND.n820 GND.n544 9.3005
R3996 GND.n819 GND.n818 9.3005
R3997 GND.n817 GND.n545 9.3005
R3998 GND.n816 GND.n815 9.3005
R3999 GND.n814 GND.n813 9.3005
R4000 GND.n812 GND.n546 9.3005
R4001 GND.n811 GND.n810 9.3005
R4002 GND.n809 GND.n548 9.3005
R4003 GND.n808 GND.n807 9.3005
R4004 GND.n806 GND.n549 9.3005
R4005 GND.n805 GND.n804 9.3005
R4006 GND.n803 GND.n802 9.3005
R4007 GND.n801 GND.n550 9.3005
R4008 GND.n800 GND.n799 9.3005
R4009 GND.n798 GND.n552 9.3005
R4010 GND.n797 GND.n796 9.3005
R4011 GND.n795 GND.n553 9.3005
R4012 GND.n794 GND.n793 9.3005
R4013 GND.n792 GND.n791 9.3005
R4014 GND.n790 GND.n554 9.3005
R4015 GND.n789 GND.n788 9.3005
R4016 GND.n787 GND.n556 9.3005
R4017 GND.n786 GND.n785 9.3005
R4018 GND.n784 GND.n557 9.3005
R4019 GND.n783 GND.n782 9.3005
R4020 GND.n781 GND.n780 9.3005
R4021 GND.n779 GND.n558 9.3005
R4022 GND.n778 GND.n777 9.3005
R4023 GND.n776 GND.n560 9.3005
R4024 GND.n775 GND.n774 9.3005
R4025 GND.n773 GND.n561 9.3005
R4026 GND.n772 GND.n771 9.3005
R4027 GND.n770 GND.n769 9.3005
R4028 GND.n768 GND.n562 9.3005
R4029 GND.n767 GND.n766 9.3005
R4030 GND.n765 GND.n564 9.3005
R4031 GND.n764 GND.n763 9.3005
R4032 GND.n762 GND.n565 9.3005
R4033 GND.n761 GND.n760 9.3005
R4034 GND.n759 GND.n758 9.3005
R4035 GND.n757 GND.n566 9.3005
R4036 GND.n756 GND.n755 9.3005
R4037 GND.n754 GND.n568 9.3005
R4038 GND.n753 GND.n752 9.3005
R4039 GND.n751 GND.n569 9.3005
R4040 GND.n750 GND.n749 9.3005
R4041 GND.n748 GND.n747 9.3005
R4042 GND.n746 GND.n570 9.3005
R4043 GND.n745 GND.n744 9.3005
R4044 GND.n743 GND.n572 9.3005
R4045 GND.n742 GND.n741 9.3005
R4046 GND.n740 GND.n573 9.3005
R4047 GND.n739 GND.n738 9.3005
R4048 GND.n737 GND.n736 9.3005
R4049 GND.n735 GND.n574 9.3005
R4050 GND.n734 GND.n733 9.3005
R4051 GND.n732 GND.n576 9.3005
R4052 GND.n731 GND.n730 9.3005
R4053 GND.n729 GND.n577 9.3005
R4054 GND.n728 GND.n727 9.3005
R4055 GND.n726 GND.n725 9.3005
R4056 GND.n1572 GND.n196 9.14112
R4057 GND.n1566 GND.n196 9.14112
R4058 GND.n581 GND.n195 9.14112
R4059 GND.n1566 GND.n195 9.14112
R4060 GND.n1267 GND.n1218 9.03579
R4061 GND.n339 GND.n338 8.94409
R4062 GND.n1866 GND.n9 8.93905
R4063 GND.t516 GND.t13 8.87896
R4064 GND.n54 GND.n53 8.85258
R4065 GND.n55 GND.n54 8.84842
R4066 GND.n619 GND.t86 8.7005
R4067 GND.n619 GND.t40 8.7005
R4068 GND.n628 GND.t744 8.7005
R4069 GND.n628 GND.t903 8.7005
R4070 GND.n607 GND.t834 8.7005
R4071 GND.n607 GND.t104 8.7005
R4072 GND.n599 GND.t532 8.7005
R4073 GND.n599 GND.t21 8.7005
R4074 GND.n650 GND.t426 8.7005
R4075 GND.n650 GND.t946 8.7005
R4076 GND.n623 GND.t926 8.7005
R4077 GND.n623 GND.t500 8.7005
R4078 GND.n205 GND.n203 8.47876
R4079 GND.t784 GND.n205 8.47876
R4080 GND.n1539 GND.n1538 8.47876
R4081 GND.t708 GND.n1539 8.47876
R4082 GND.n233 GND.n232 8.47876
R4083 GND.t160 GND.n233 8.47876
R4084 GND.n1557 GND.n207 8.47876
R4085 GND.n1557 GND.t784 8.47876
R4086 GND.n1541 GND.n1540 8.47876
R4087 GND.n1540 GND.t708 8.47876
R4088 GND.n1512 GND.n1511 8.47876
R4089 GND.n1511 GND.t160 8.47876
R4090 GND.n1120 GND.t514 8.46601
R4091 GND.n1423 GND.t686 8.46601
R4092 GND.n1444 GND.t767 8.46601
R4093 GND.n1475 GND.t145 7.64011
R4094 GND.t526 GND.n1113 7.64011
R4095 GND.t702 GND.t51 7.3212
R4096 GND.t705 GND.t571 7.3212
R4097 GND.t115 GND.t53 7.3212
R4098 GND.t708 GND.t50 7.3212
R4099 GND.t401 GND.t52 7.3212
R4100 GND.n1548 GND.n1547 7.13465
R4101 GND.n1549 GND.n1548 7.13465
R4102 GND.n1551 GND.n1550 7.13465
R4103 GND.n1550 GND.n1549 7.13465
R4104 GND.t968 GND.n1119 7.02068
R4105 GND.t621 GND.n1087 6.8142
R4106 GND.n1226 GND.n1221 6.77697
R4107 GND.n1228 GND.n1219 6.77697
R4108 GND.n1297 GND.n376 6.77697
R4109 GND.n1288 GND.n378 6.77697
R4110 GND.n522 GND.n497 6.77697
R4111 GND.n1122 GND.n231 6.44556
R4112 GND.n133 GND 6.4005
R4113 GND.n1528 GND.n1527 6.31845
R4114 GND.t608 GND.n1045 6.19477
R4115 GND.t930 GND.t623 6.19477
R4116 GND.t626 GND.t928 6.19477
R4117 GND.t107 GND.t525 6.19477
R4118 GND.t519 GND.t22 6.01393
R4119 GND.n1474 GND.t361 5.9883
R4120 GND.n492 GND.t582 5.8005
R4121 GND.n492 GND.t726 5.8005
R4122 GND.n481 GND.t754 5.8005
R4123 GND.n481 GND.t810 5.8005
R4124 GND.n482 GND.t959 5.8005
R4125 GND.n482 GND.t521 5.8005
R4126 GND.n472 GND.t544 5.8005
R4127 GND.n472 GND.t944 5.8005
R4128 GND.n470 GND.t774 5.8005
R4129 GND.n470 GND.t843 5.8005
R4130 GND.n462 GND.t2 5.8005
R4131 GND.n462 GND.t870 5.8005
R4132 GND.n463 GND.t569 5.8005
R4133 GND.n463 GND.t692 5.8005
R4134 GND.n455 GND.t897 5.8005
R4135 GND.n455 GND.t383 5.8005
R4136 GND.n453 GND.t16 5.8005
R4137 GND.n453 GND.t639 5.8005
R4138 GND.n674 GND.t505 5.8005
R4139 GND.n674 GND.t881 5.8005
R4140 GND.n673 GND.t740 5.8005
R4141 GND.n673 GND.t793 5.8005
R4142 GND.n1861 GND.n1860 5.79258
R4143 GND.n1860 GND.n10 5.79258
R4144 GND.n1851 GND.n1847 5.79258
R4145 GND.n1851 GND.n1850 5.79258
R4146 GND.t771 GND.n1126 5.78182
R4147 GND.n132 GND.t271 5.6932
R4148 GND.n1600 GND.n27 5.68011
R4149 GND.n1600 GND.n10 5.68011
R4150 GND.n1699 GND.n1673 5.68011
R4151 GND.n1673 GND.n10 5.68011
R4152 GND.n1717 GND.n1716 5.68011
R4153 GND.n1716 GND.n10 5.68011
R4154 GND.t367 GND.t929 5.36887
R4155 GND.n604 GND.n603 5.21334
R4156 GND.n652 GND.n616 5.21334
R4157 GND.n635 GND.n625 5.21334
R4158 GND.n1465 GND.t629 4.95592
R4159 GND.n1432 GND.n1431 4.89462
R4160 GND.n1437 GND.n1436 4.89462
R4161 GND.n1442 GND.n1441 4.89462
R4162 GND.n1102 GND.n1101 4.89462
R4163 GND.n1108 GND.n1107 4.89462
R4164 GND.n1748 GND.n19 4.89462
R4165 GND.n1709 GND.n1618 4.89462
R4166 GND.n1854 GND.n28 4.89462
R4167 GND.n1701 GND.n30 4.89462
R4168 GND.n1620 GND.n15 4.86612
R4169 GND.n166 GND.n15 4.86612
R4170 GND.n1718 GND.n177 4.57238
R4171 GND.n1727 GND.n1718 4.57238
R4172 GND.t684 GND.t596 4.54297
R4173 GND.t525 GND.t685 4.54297
R4174 GND.n1140 GND.t516 4.54297
R4175 GND.n234 GND.t705 4.44521
R4176 GND.n6 GND.n4 4.36617
R4177 GND.n1848 GND.n6 4.36617
R4178 GND.n5 GND.n3 4.36617
R4179 GND.n1849 GND.n5 4.36617
R4180 GND.n1323 GND.n1322 4.33704
R4181 GND.n837 GND.n836 4.33704
R4182 GND.t13 GND.t108 4.33649
R4183 GND.n1126 GND.t698 4.33649
R4184 GND.t919 GND.t506 4.2218
R4185 GND.n1735 GND.n1734 4.2218
R4186 GND.t462 GND.t920 4.2218
R4187 GND.n1337 GND.n1336 4.17828
R4188 GND.n1335 GND.n1334 4.17828
R4189 GND.n722 GND.n595 4.14696
R4190 GND.n1465 GND.n1464 4.13002
R4191 GND.n1273 GND.n1272 4.00641
R4192 GND.t515 GND.n1444 3.92354
R4193 GND.n1840 GND.n1839 3.91726
R4194 GND.t139 GND.t130 3.72489
R4195 GND.n863 GND.n448 3.71362
R4196 GND.n1380 GND.n1379 3.52871
R4197 GND.n1329 GND.n1328 3.52871
R4198 GND.n1825 GND 3.2614
R4199 GND.t167 GND.t135 3.13794
R4200 GND.n221 GND.t777 3.13794
R4201 GND.n1272 GND.n1271 3.13461
R4202 GND.n1452 GND.n1451 3.1005
R4203 GND.n1380 GND.n1333 3.09574
R4204 GND.n1365 GND.n1333 3.09574
R4205 GND.n1344 GND.n1332 3.09574
R4206 GND.n1365 GND.n1332 3.09574
R4207 GND.n1331 GND.n1329 2.9255
R4208 GND.n1331 GND.n1330 2.9255
R4209 GND.n338 GND.n334 2.9255
R4210 GND.n1330 GND.n334 2.9255
R4211 GND.n594 GND.n593 2.87229
R4212 GND.n1322 GND 2.85076
R4213 GND GND.n1312 2.85076
R4214 GND GND.n365 2.85076
R4215 GND.n1327 GND.n1324 2.82946
R4216 GND.t80 GND.t6 2.61503
R4217 GND.n721 GND.n596 2.5255
R4218 GND.n1527 GND.n200 2.51123
R4219 GND.n234 GND.n200 2.51123
R4220 GND.n587 GND.n199 2.51123
R4221 GND.n235 GND.n199 2.51123
R4222 GND.n1460 GND.n282 2.50988
R4223 GND.t860 GND.t859 2.47821
R4224 GND.n1771 GND.n1770 2.42212
R4225 GND.n1122 GND.t635 2.41134
R4226 GND.n582 GND.n581 2.33946
R4227 GND.n595 GND.n594 2.33946
R4228 GND.n1379 GND.n0 2.33915
R4229 GND.n1328 GND.n1327 2.33915
R4230 GND.n722 GND.n721 2.33654
R4231 GND GND.n1872 2.27362
R4232 GND.n595 GND.n582 2.25133
R4233 GND.n838 GND.n837 2.2505
R4234 GND.n1096 GND.n1095 2.23675
R4235 GND.n723 GND.n722 2.20779
R4236 GND.n1400 GND.n1399 2.13383
R4237 GND.t396 GND.t799 2.06526
R4238 GND.n712 GND.n604 2.04483
R4239 GND.n638 GND.n625 2.04483
R4240 GND.n693 GND.n616 2.04483
R4241 GND.n836 GND.n835 1.9555
R4242 GND.n1324 GND.n364 1.94363
R4243 GND.n1106 GND.n275 1.92706
R4244 GND.n1468 GND.n275 1.92706
R4245 GND.n1098 GND.n1097 1.92081
R4246 GND.n1099 GND.n1098 1.89738
R4247 GND GND.n186 1.89588
R4248 GND.n1428 GND.n289 1.87081
R4249 GND.n446 GND.n445 1.8605
R4250 GND.n443 GND.n442 1.8605
R4251 GND.n1101 GND.n1100 1.8605
R4252 GND.n1441 GND.n1440 1.8605
R4253 GND.n1457 GND.n1456 1.8605
R4254 GND.n1117 GND.n274 1.8605
R4255 GND.n1091 GND.t628 1.85878
R4256 GND GND.n491 1.85258
R4257 GND.n489 GND 1.85258
R4258 GND.n487 GND 1.85258
R4259 GND GND.n471 1.85258
R4260 GND GND.n469 1.85258
R4261 GND.n467 GND 1.85258
R4262 GND.n465 GND 1.85258
R4263 GND.n856 GND 1.85258
R4264 GND.n858 GND 1.85258
R4265 GND GND.n449 1.85258
R4266 GND.n1326 GND.n0 1.84196
R4267 GND.n444 GND.n440 1.788
R4268 GND.n1872 GND.n1871 1.7528
R4269 GND.n435 GND.t629 1.65231
R4270 GND.t110 GND.n1422 1.65231
R4271 GND.t877 GND.t501 1.55171
R4272 GND.n836 GND 1.52425
R4273 GND.n1872 GND.n0 1.51654
R4274 GND.n723 GND.n364 1.48404
R4275 GND.n1450 GND.n289 1.4755
R4276 GND.t548 GND.t387 1.45963
R4277 GND.n1741 GND.n1740 1.44894
R4278 GND.n1105 GND.t367 1.44583
R4279 GND.n1475 GND.n1474 1.44583
R4280 GND.n438 GND.n284 1.3755
R4281 GND.n1805 GND.n1791 1.27784
R4282 GND.n1445 GND.t106 1.23936
R4283 GND.n1470 GND.n273 1.21613
R4284 GND.n1862 GND.n1861 1.21131
R4285 GND.n1041 GND.n863 1.17175
R4286 GND.n1041 GND.n1040 1.15253
R4287 GND GND.n838 1.13527
R4288 GND.n1308 GND.n1307 1.12991
R4289 GND.n1728 GND.n168 1.12238
R4290 GND.n1692 GND.n168 1.12238
R4291 GND.n1324 GND.n1323 1.10279
R4292 GND.n117 GND.t312 1.082
R4293 GND.n1327 GND.n1326 1.0655
R4294 GND.n1429 GND.n1428 1.04894
R4295 GND.n1742 GND.n1741 1.04581
R4296 GND.n1438 GND.n1437 1.03383
R4297 GND.n307 GND.t393 1.03288
R4298 GND.n1470 GND.n1469 0.984875
R4299 GND.n1095 GND 0.977696
R4300 GND.n1469 GND.n1468 0.942687
R4301 GND.n1837 GND.n1836 0.9305
R4302 GND.n1870 GND.n1869 0.9305
R4303 GND.n1679 GND.n1677 0.91925
R4304 GND.n1681 GND.n1679 0.91925
R4305 GND.n1683 GND.n1681 0.91925
R4306 GND.n1698 GND.n1697 0.91925
R4307 GND.n1697 GND.n1696 0.91925
R4308 GND.n1696 GND.n1695 0.91925
R4309 GND.n1695 GND.n1694 0.91925
R4310 GND.n1653 GND.n1652 0.91925
R4311 GND.n1652 GND.n1651 0.91925
R4312 GND.n1651 GND.n1650 0.91925
R4313 GND.n1658 GND.n1657 0.91925
R4314 GND.n1657 GND.n1656 0.91925
R4315 GND.n1656 GND.n1655 0.91925
R4316 GND.n126 GND.t301 0.909177
R4317 GND.n1822 GND.n147 0.908052
R4318 GND.n1837 GND.n132 0.873417
R4319 GND.n1322 GND.n365 0.872295
R4320 GND.n724 GND.n448 0.857375
R4321 GND.n838 GND.n538 0.856945
R4322 GND.n1312 GND 0.846654
R4323 GND.n1830 GND.n138 0.845955
R4324 GND.n1817 GND.n145 0.845955
R4325 GND.n1460 GND.n1459 0.839563
R4326 GND.n1823 GND.n1822 0.833625
R4327 GND.n142 GND.n138 0.8255
R4328 GND.n145 GND.n144 0.8255
R4329 GND.n1430 GND.n1429 0.822375
R4330 GND.n1430 GND.n299 0.822375
R4331 GND.n1784 GND.n1783 0.821833
R4332 GND.n1593 GND.n1592 0.810441
R4333 GND.n1801 GND.n1800 0.788781
R4334 GND.n1798 GND.n1797 0.788781
R4335 GND.n1789 GND.n1788 0.788781
R4336 GND.n1698 GND 0.780188
R4337 GND.n1744 GND.n1743 0.7755
R4338 GND.n1740 GND.n1730 0.7755
R4339 GND.n1828 GND.n1827 0.7755
R4340 GND.n143 GND.n137 0.7755
R4341 GND.n1307 GND.n370 0.753441
R4342 GND.n1095 GND.n1041 0.744875
R4343 GND.n1838 GND.n1837 0.74425
R4344 GND.n71 GND.t186 0.7295
R4345 GND.n73 GND.t343 0.7295
R4346 GND.n75 GND.t180 0.7295
R4347 GND.n77 GND.t330 0.7295
R4348 GND.n79 GND.t314 0.7295
R4349 GND.n81 GND.t305 0.7295
R4350 GND.n83 GND.t227 0.7295
R4351 GND.n85 GND.t254 0.7295
R4352 GND.n87 GND.t345 0.7295
R4353 GND.n94 GND.t221 0.7295
R4354 GND.n64 GND.t188 0.7295
R4355 GND.n63 GND.t281 0.7295
R4356 GND.n62 GND.t256 0.7295
R4357 GND.n61 GND.t200 0.7295
R4358 GND.n96 GND.t310 0.7295
R4359 GND.n98 GND.t303 0.7295
R4360 GND.n100 GND.t349 0.7295
R4361 GND.n102 GND.t198 0.7295
R4362 GND.n104 GND.t211 0.7295
R4363 GND.n106 GND.t245 0.7295
R4364 GND.n70 GND.t209 0.7295
R4365 GND.n69 GND.t325 0.7295
R4366 GND.n68 GND.t277 0.7295
R4367 GND.n59 GND.t213 0.7295
R4368 GND.n108 GND.t215 0.7295
R4369 GND.n110 GND.t247 0.7295
R4370 GND.n112 GND.t287 0.7295
R4371 GND.n114 GND.t354 0.7295
R4372 GND.n116 GND.t202 0.7295
R4373 GND.n127 GND.t285 0.7295
R4374 GND.n129 GND.t279 0.7295
R4375 GND.n120 GND.t347 0.7295
R4376 GND.n117 GND.t258 0.7295
R4377 GND.n118 GND.t204 0.7295
R4378 GND.n119 GND.t283 0.7295
R4379 GND.t271 GND.n131 0.7295
R4380 GND.n1107 GND.n1106 0.715885
R4381 GND.n1468 GND.n1467 0.715885
R4382 GND.n1856 GND.n26 0.715885
R4383 GND.n1704 GND.n1703 0.715885
R4384 GND.n50 GND.n28 0.715885
R4385 GND.n1623 GND.n30 0.715885
R4386 GND.n1106 GND.n273 0.711438
R4387 GND.n1692 GND.n26 0.709875
R4388 GND.n1636 GND.n26 0.709875
R4389 GND.n1636 GND.n50 0.709875
R4390 GND.n1840 GND.n50 0.709875
R4391 GND.n1741 GND.n1738 0.664786
R4392 GND.n1746 GND.n1745 0.664786
R4393 GND.n1272 GND 0.661558
R4394 GND.n676 GND 0.645031
R4395 GND GND.n675 0.645031
R4396 GND.n675 GND 0.645031
R4397 GND.n454 GND 0.645031
R4398 GND GND.n454 0.645031
R4399 GND GND.n855 0.645031
R4400 GND.n855 GND 0.645031
R4401 GND.n464 GND 0.645031
R4402 GND GND.n464 0.645031
R4403 GND.n849 GND 0.645031
R4404 GND.n849 GND 0.645031
R4405 GND GND.n848 0.645031
R4406 GND.n848 GND 0.645031
R4407 GND GND.n847 0.645031
R4408 GND.n847 GND 0.645031
R4409 GND.n483 GND 0.645031
R4410 GND GND.n483 0.645031
R4411 GND.n840 GND 0.645031
R4412 GND.n840 GND 0.645031
R4413 GND GND.n839 0.645031
R4414 GND GND.n1188 0.633946
R4415 GND.n1155 GND 0.633946
R4416 GND GND.n1173 0.633946
R4417 GND.n861 GND.n450 0.625711
R4418 GND.n1431 GND.n1430 0.6205
R4419 GND.n1426 GND.n289 0.6205
R4420 GND.t698 GND.t106 0.619928
R4421 GND.n167 GND.n166 0.615539
R4422 GND.n1743 GND.n1729 0.609875
R4423 GND.n839 GND 0.608898
R4424 GND.n678 GND.n677 0.607197
R4425 GND GND.n138 0.603625
R4426 GND.n1458 GND.n283 0.59425
R4427 GND.n299 GND.n291 0.59425
R4428 GND.n1728 GND.n1727 0.59425
R4429 GND.n1637 GND.n1636 0.59425
R4430 GND.n1822 GND.n1821 0.58175
R4431 GND.n1806 GND.n1805 0.58175
R4432 GND.n1439 GND.n1438 0.568786
R4433 GND.n1326 GND.n1325 0.555206
R4434 GND.n835 GND.n364 0.552583
R4435 GND.n724 GND.n723 0.552583
R4436 GND.n1323 GND 0.5405
R4437 GND.n1707 GND.n177 0.53175
R4438 GND.n1672 GND.n1671 0.53175
R4439 GND GND.n1199 0.51148
R4440 GND.n41 GND.n40 0.51137
R4441 GND.n42 GND.n41 0.51137
R4442 GND.n43 GND.n42 0.51137
R4443 GND.n1846 GND.n43 0.51137
R4444 GND.n1846 GND.n1845 0.51137
R4445 GND.n1843 GND.n1842 0.51137
R4446 GND.n1842 GND.n1841 0.51137
R4447 GND.n1449 GND.n1448 0.489974
R4448 GND.n1428 GND.n1427 0.489974
R4449 GND.n298 GND.n283 0.48175
R4450 GND.n1312 GND 0.473256
R4451 GND.n1655 GND.n1654 0.459875
R4452 GND.n1654 GND.n1653 0.459875
R4453 GND.n1438 GND.n299 0.448938
R4454 GND.n1748 GND.n1747 0.443357
R4455 GND.n179 GND.n168 0.443357
R4456 GND.n1706 GND.n182 0.443357
R4457 GND.n1709 GND.n1708 0.443357
R4458 GND.n1708 GND.n1620 0.429028
R4459 GND.n1871 GND.n1 0.4255
R4460 GND.n276 GND.n275 0.423227
R4461 GND.n1471 GND.n1470 0.423227
R4462 GND.n1743 GND.n1742 0.403625
R4463 GND.n1740 GND.n1739 0.403625
R4464 GND.n1800 GND.n1799 0.403625
R4465 GND.n1799 GND.n1798 0.403625
R4466 GND.n1827 GND.n141 0.403625
R4467 GND.n1827 GND.n1826 0.403625
R4468 GND.n143 GND.n142 0.403625
R4469 GND.n144 GND.n143 0.403625
R4470 GND.n1788 GND.n1787 0.403625
R4471 GND.n1787 GND.n1784 0.403625
R4472 GND.n1450 GND.n1449 0.395812
R4473 GND.n1804 GND 0.392688
R4474 GND.n883 GND 0.390703
R4475 GND GND.n1014 0.390703
R4476 GND.n915 GND 0.390703
R4477 GND GND.n986 0.390703
R4478 GND.n947 GND 0.390703
R4479 GND GND.n395 0.390703
R4480 GND.n1279 GND.n1278 0.376971
R4481 GND.n1804 GND.n1803 0.368469
R4482 GND.n132 GND.n57 0.360917
R4483 GND.n1805 GND.n1804 0.359875
R4484 GND.n64 GND.n63 0.353
R4485 GND.n63 GND.n62 0.353
R4486 GND.n62 GND.n61 0.353
R4487 GND.n70 GND.n69 0.353
R4488 GND.n69 GND.n68 0.353
R4489 GND.n68 GND.n59 0.353
R4490 GND.n118 GND.n117 0.353
R4491 GND.n119 GND.n118 0.353
R4492 GND.n1622 GND.n1621 0.338152
R4493 GND.n1620 GND.n1619 0.338152
R4494 GND.n166 GND.n165 0.338152
R4495 GND.n177 GND.n172 0.338152
R4496 GND.n177 GND.n176 0.338152
R4497 GND.n1727 GND.n1722 0.338152
R4498 GND.n1727 GND.n1726 0.338152
R4499 GND.n1693 GND.n1691 0.338152
R4500 GND.n1825 GND.n145 0.332591
R4501 GND.n1650 GND.n1637 0.33175
R4502 GND.n1671 GND.n1658 0.33175
R4503 GND.n87 GND.n64 0.3295
R4504 GND.n94 GND.n61 0.3295
R4505 GND.n75 GND.n70 0.3295
R4506 GND.n106 GND.n59 0.3295
R4507 GND.n120 GND.n119 0.3295
R4508 GND.n1841 GND.n1840 0.314359
R4509 GND.n1693 GND.n1692 0.3005
R4510 GND.n1679 GND.n1678 0.291659
R4511 GND.n1681 GND.n1680 0.291659
R4512 GND.n1683 GND.n1682 0.291659
R4513 GND.n1698 GND.n1684 0.291659
R4514 GND.n1697 GND.n1685 0.291659
R4515 GND.n1696 GND.n1686 0.291659
R4516 GND.n1695 GND.n1687 0.291659
R4517 GND.n1653 GND.n1630 0.291659
R4518 GND.n1653 GND.n1631 0.291659
R4519 GND.n1652 GND.n1632 0.291659
R4520 GND.n1652 GND.n1633 0.291659
R4521 GND.n1651 GND.n1634 0.291659
R4522 GND.n1651 GND.n1635 0.291659
R4523 GND.n1657 GND.n1624 0.291659
R4524 GND.n1657 GND.n1625 0.291659
R4525 GND.n1656 GND.n1626 0.291659
R4526 GND.n1656 GND.n1627 0.291659
R4527 GND.n1655 GND.n1628 0.291659
R4528 GND.n1655 GND.n1629 0.291659
R4529 GND.n1115 GND.n440 0.291125
R4530 GND.n1670 GND.n1665 0.288543
R4531 GND.n37 GND.n35 0.288543
R4532 GND.n49 GND.n47 0.288543
R4533 GND.n1676 GND.n1674 0.288543
R4534 GND.n176 GND.n173 0.288543
R4535 GND.n176 GND.n174 0.288543
R4536 GND.n172 GND.n169 0.288543
R4537 GND.n172 GND.n170 0.288543
R4538 GND.n1726 GND.n1723 0.288543
R4539 GND.n1726 GND.n1724 0.288543
R4540 GND.n1722 GND.n1719 0.288543
R4541 GND.n1722 GND.n1720 0.288543
R4542 GND.n1690 GND.n1688 0.288543
R4543 GND.n1646 GND.n1644 0.288543
R4544 GND.n1649 GND.n1647 0.288543
R4545 GND.n1647 GND.n1646 0.288543
R4546 GND.n1641 GND.n1639 0.288543
R4547 GND.n1643 GND.n1642 0.288543
R4548 GND.n1642 GND.n1641 0.288543
R4549 GND.n1664 GND.n1661 0.288543
R4550 GND.n1661 GND.n1660 0.288543
R4551 GND.n1664 GND.n1662 0.288543
R4552 GND.n1670 GND.n1669 0.288543
R4553 GND.n1669 GND.n1668 0.288543
R4554 GND.n67 GND.t208 0.28175
R4555 GND.n66 GND.t324 0.28175
R4556 GND.n65 GND.t276 0.28175
R4557 GND.n60 GND.t212 0.28175
R4558 GND.n130 GND.t278 0.28175
R4559 GND.n128 GND.t284 0.28175
R4560 GND.n126 GND.t300 0.28175
R4561 GND.n125 GND.t311 0.28175
R4562 GND.n124 GND.t257 0.28175
R4563 GND.n123 GND.t203 0.28175
R4564 GND.n122 GND.t282 0.28175
R4565 GND.n121 GND.t346 0.28175
R4566 GND.n115 GND.t201 0.28175
R4567 GND.n113 GND.t353 0.28175
R4568 GND.n111 GND.t286 0.28175
R4569 GND.n109 GND.t246 0.28175
R4570 GND.n107 GND.t214 0.28175
R4571 GND.n105 GND.t244 0.28175
R4572 GND.n103 GND.t210 0.28175
R4573 GND.n101 GND.t197 0.28175
R4574 GND.n99 GND.t348 0.28175
R4575 GND.n97 GND.t302 0.28175
R4576 GND.n95 GND.t309 0.28175
R4577 GND.n93 GND.t220 0.28175
R4578 GND.n92 GND.t199 0.28175
R4579 GND.n91 GND.t255 0.28175
R4580 GND.n90 GND.t280 0.28175
R4581 GND.n89 GND.t187 0.28175
R4582 GND.n88 GND.t344 0.28175
R4583 GND.n86 GND.t253 0.28175
R4584 GND.n84 GND.t226 0.28175
R4585 GND.n82 GND.t304 0.28175
R4586 GND.n80 GND.t313 0.28175
R4587 GND.n78 GND.t329 0.28175
R4588 GND.n76 GND.t179 0.28175
R4589 GND.n74 GND.t342 0.28175
R4590 GND.n72 GND.t185 0.28175
R4591 GND.n58 GND.t270 0.28175
R4592 GND.n1839 GND 0.271125
R4593 GND.n1845 GND.n1844 0.263408
R4594 GND.n235 GND.n234 0.261953
R4595 GND.t693 GND.t80 0.261953
R4596 GND.n1846 GND.n31 0.261171
R4597 GND.n41 GND.n34 0.261171
R4598 GND.n42 GND.n33 0.261171
R4599 GND.n43 GND.n32 0.261171
R4600 GND.n1845 GND.n44 0.261171
R4601 GND.n1843 GND.n45 0.261171
R4602 GND.n1842 GND.n46 0.261171
R4603 GND.n1100 GND.n1099 0.259875
R4604 GND.n1799 GND.n149 0.251851
R4605 GND.n1787 GND.n1786 0.251851
R4606 GND.n1844 GND.n1843 0.248462
R4607 GND.n67 GND.n66 0.242354
R4608 GND.n66 GND.n65 0.242354
R4609 GND.n65 GND.n60 0.242354
R4610 GND.n125 GND.n124 0.242354
R4611 GND.n124 GND.n123 0.242354
R4612 GND.n123 GND.n122 0.242354
R4613 GND.n92 GND.n91 0.242354
R4614 GND.n91 GND.n90 0.242354
R4615 GND.n90 GND.n89 0.242354
R4616 GND.n1098 GND.n297 0.238962
R4617 GND.n1705 GND.n1622 0.238
R4618 GND.n1100 GND.n282 0.236438
R4619 GND.n444 GND.n443 0.23175
R4620 GND.n1457 GND.n284 0.23175
R4621 GND.n443 GND.n282 0.230187
R4622 GND.n445 GND.n273 0.230187
R4623 GND.n1458 GND.n1457 0.230187
R4624 GND.n1469 GND.n274 0.230187
R4625 GND.n445 GND.n444 0.228625
R4626 GND.n438 GND.n274 0.228625
R4627 GND.n1459 GND.n1458 0.227062
R4628 GND.n439 GND.n438 0.227062
R4629 GND.n141 GND 0.222375
R4630 GND.n76 GND.n67 0.218854
R4631 GND.n105 GND.n60 0.218854
R4632 GND.n126 GND.n125 0.218854
R4633 GND.n122 GND.n121 0.218854
R4634 GND.n93 GND.n92 0.218854
R4635 GND.n89 GND.n88 0.218854
R4636 GND.n837 GND 0.211237
R4637 GND.n1461 GND.n1460 0.207167
R4638 GND.t45 GND.t361 0.206976
R4639 GND.t799 GND.t514 0.206976
R4640 GND.n1119 GND.t684 0.206976
R4641 GND.n1454 GND.t108 0.206976
R4642 GND.n1739 GND.n167 0.20675
R4643 GND.n1826 GND.n1825 0.20675
R4644 GND.n131 GND.n130 0.205635
R4645 GND.n129 GND.n128 0.205635
R4646 GND.n127 GND.n126 0.205635
R4647 GND.n121 GND.n116 0.205635
R4648 GND.n115 GND.n114 0.205635
R4649 GND.n113 GND.n112 0.205635
R4650 GND.n111 GND.n110 0.205635
R4651 GND.n109 GND.n108 0.205635
R4652 GND.n107 GND.n106 0.205635
R4653 GND.n105 GND.n104 0.205635
R4654 GND.n103 GND.n102 0.205635
R4655 GND.n101 GND.n100 0.205635
R4656 GND.n99 GND.n98 0.205635
R4657 GND.n97 GND.n96 0.205635
R4658 GND.n95 GND.n94 0.205635
R4659 GND.n87 GND.n86 0.205635
R4660 GND.n85 GND.n84 0.205635
R4661 GND.n83 GND.n82 0.205635
R4662 GND.n81 GND.n80 0.205635
R4663 GND.n79 GND.n78 0.205635
R4664 GND.n77 GND.n76 0.205635
R4665 GND.n75 GND.n74 0.205635
R4666 GND.n73 GND.n72 0.205635
R4667 GND.n71 GND.n58 0.205635
R4668 GND.n1677 GND.n1676 0.204006
R4669 GND.n1694 GND.n1690 0.204006
R4670 GND.n1650 GND.n1643 0.204006
R4671 GND.n1650 GND.n1649 0.204006
R4672 GND.n1641 GND.n1637 0.204006
R4673 GND.n1646 GND.n1637 0.204006
R4674 GND.n1671 GND.n1664 0.204006
R4675 GND.n1671 GND.n1670 0.204006
R4676 GND.n1660 GND.n1658 0.204006
R4677 GND.n1668 GND.n1658 0.204006
R4678 GND.n1449 GND.n291 0.198937
R4679 GND.n596 GND.n448 0.196125
R4680 GND.n1708 GND.n1707 0.191528
R4681 GND.n1707 GND.n1706 0.191528
R4682 GND.n1706 GND.n1705 0.191528
R4683 GND.n440 GND.n439 0.186437
R4684 GND.n130 GND.n129 0.180177
R4685 GND.n128 GND.n127 0.180177
R4686 GND.n121 GND.n120 0.180177
R4687 GND.n116 GND.n115 0.180177
R4688 GND.n114 GND.n113 0.180177
R4689 GND.n112 GND.n111 0.180177
R4690 GND.n110 GND.n109 0.180177
R4691 GND.n108 GND.n107 0.180177
R4692 GND.n106 GND.n105 0.180177
R4693 GND.n104 GND.n103 0.180177
R4694 GND.n102 GND.n101 0.180177
R4695 GND.n100 GND.n99 0.180177
R4696 GND.n98 GND.n97 0.180177
R4697 GND.n96 GND.n95 0.180177
R4698 GND.n94 GND.n93 0.180177
R4699 GND.n88 GND.n87 0.180177
R4700 GND.n86 GND.n85 0.180177
R4701 GND.n84 GND.n83 0.180177
R4702 GND.n82 GND.n81 0.180177
R4703 GND.n80 GND.n79 0.180177
R4704 GND.n78 GND.n77 0.180177
R4705 GND.n76 GND.n75 0.180177
R4706 GND.n74 GND.n73 0.180177
R4707 GND.n72 GND.n71 0.180177
R4708 GND.n131 GND.n58 0.180177
R4709 GND.n39 GND.n2 0.175092
R4710 GND.n40 GND.n37 0.173518
R4711 GND.n1841 GND.n49 0.173518
R4712 GND.n594 GND.n587 0.164603
R4713 GND.n1097 GND.n283 0.164562
R4714 GND.n291 GND.n290 0.159799
R4715 GND.n1451 GND.n1450 0.15675
R4716 GND.n1451 GND.n284 0.155187
R4717 GND.n1729 GND.n1728 0.146789
R4718 GND GND.n1683 0.139562
R4719 GND.n1746 GND.n1729 0.139475
R4720 GND.n1623 GND.n2 0.138101
R4721 GND.n1747 GND.n167 0.1255
R4722 GND.n1705 GND.n1704 0.124996
R4723 GND.n1704 GND.n1672 0.124996
R4724 GND.n1672 GND.n1623 0.124996
R4725 GND.n719 GND.n598 0.120292
R4726 GND.n714 GND.n713 0.120292
R4727 GND.n711 GND.n605 0.120292
R4728 GND.n705 GND.n704 0.120292
R4729 GND.n630 GND.n629 0.120292
R4730 GND.n637 GND.n626 0.120292
R4731 GND.n639 GND.n624 0.120292
R4732 GND.n646 GND.n645 0.120292
R4733 GND.n660 GND.n659 0.120292
R4734 GND.n655 GND.n615 0.120292
R4735 GND.n692 GND.n617 0.120292
R4736 GND.n686 GND.n685 0.120292
R4737 GND.n536 GND.n535 0.120292
R4738 GND.n535 GND.n534 0.120292
R4739 GND.n534 GND.n494 0.120292
R4740 GND.n530 GND.n494 0.120292
R4741 GND.n530 GND.n529 0.120292
R4742 GND.n529 GND.n528 0.120292
R4743 GND.n525 GND.n524 0.120292
R4744 GND.n524 GND.n523 0.120292
R4745 GND.n520 GND.n519 0.120292
R4746 GND.n519 GND.n518 0.120292
R4747 GND.n518 GND.n499 0.120292
R4748 GND.n513 GND.n512 0.120292
R4749 GND.n512 GND.n511 0.120292
R4750 GND.n508 GND.n507 0.120292
R4751 GND.n507 GND.n506 0.120292
R4752 GND.n383 GND.n382 0.120292
R4753 GND.n1280 GND.n382 0.120292
R4754 GND.n1287 GND.n1286 0.120292
R4755 GND.n1296 GND.n1295 0.120292
R4756 GND.n375 GND.n374 0.120292
R4757 GND.n1301 GND.n374 0.120292
R4758 GND.n1303 GND.n372 0.120292
R4759 GND.n1310 GND.n371 0.120292
R4760 GND.n1311 GND.n1310 0.120292
R4761 GND.n1224 GND.n1222 0.120292
R4762 GND.n1225 GND.n1224 0.120292
R4763 GND.n1230 GND.n1220 0.120292
R4764 GND.n1231 GND.n1230 0.120292
R4765 GND.n1264 GND.n1232 0.120292
R4766 GND.n1260 GND.n1232 0.120292
R4767 GND.n1251 GND.n1237 0.120292
R4768 GND.n1246 GND.n1245 0.120292
R4769 GND.n1870 GND.n2 0.115506
R4770 GND.n1439 GND.n298 0.115419
R4771 GND.n40 GND.n39 0.112592
R4772 GND GND.n700 0.112479
R4773 GND.n661 GND 0.112479
R4774 GND.n713 GND.n712 0.109875
R4775 GND.n638 GND.n637 0.109875
R4776 GND.n693 GND.n615 0.109875
R4777 GND.n536 GND 0.105969
R4778 GND.n712 GND.n711 0.104667
R4779 GND.n639 GND.n638 0.104667
R4780 GND.n693 GND.n692 0.104667
R4781 GND.n835 GND 0.10425
R4782 GND.n1803 GND.n1802 0.101281
R4783 GND.n1802 GND.n1801 0.101281
R4784 GND.n1797 GND.n1796 0.101281
R4785 GND.n1796 GND.n147 0.101281
R4786 GND.n1791 GND.n1790 0.101281
R4787 GND.n1790 GND.n1789 0.101281
R4788 GND.n725 GND.n724 0.101125
R4789 GND.n1871 GND.n1870 0.100037
R4790 GND.n1861 GND.n15 0.0963763
R4791 GND.n1718 GND.n1717 0.0963763
R4792 GND.n1699 GND.n1698 0.0963763
R4793 GND.n1654 GND.n27 0.0963763
R4794 GND.n1847 GND.n1846 0.0963763
R4795 GND.n37 GND.n36 0.0881524
R4796 GND.n49 GND.n48 0.0881524
R4797 GND.n1676 GND.n1675 0.0881524
R4798 GND.n172 GND.n171 0.0881524
R4799 GND.n176 GND.n175 0.0881524
R4800 GND.n1722 GND.n1721 0.0881524
R4801 GND.n1726 GND.n1725 0.0881524
R4802 GND.n1690 GND.n1689 0.0881524
R4803 GND.n1643 GND.n1638 0.0881524
R4804 GND.n1649 GND.n1648 0.0881524
R4805 GND.n1641 GND.n1640 0.0881524
R4806 GND.n1646 GND.n1645 0.0881524
R4807 GND.n1664 GND.n1663 0.0881524
R4808 GND.n1670 GND.n1666 0.0881524
R4809 GND.n1660 GND.n1659 0.0881524
R4810 GND.n1668 GND.n1667 0.0881524
R4811 GND.n1061 GND 0.0866486
R4812 GND.n1060 GND.n1054 0.0815811
R4813 GND.n1069 GND.n1053 0.0815811
R4814 GND.n1078 GND.n1052 0.0815811
R4815 GND.n1094 GND.n1042 0.0815811
R4816 GND.n1040 GND.n864 0.0815811
R4817 GND.n874 GND.n873 0.0815811
R4818 GND.n884 GND.n883 0.0815811
R4819 GND.n894 GND.n893 0.0815811
R4820 GND.n1014 GND.n896 0.0815811
R4821 GND.n906 GND.n905 0.0815811
R4822 GND.n916 GND.n915 0.0815811
R4823 GND.n926 GND.n925 0.0815811
R4824 GND.n986 GND.n928 0.0815811
R4825 GND.n938 GND.n937 0.0815811
R4826 GND.n948 GND.n947 0.0815811
R4827 GND.n957 GND.n956 0.0815811
R4828 GND.n396 GND.n395 0.0815811
R4829 GND.n406 GND.n405 0.0815811
R4830 GND.n1199 GND.n408 0.0815811
R4831 GND.n1188 GND.n413 0.0815811
R4832 GND.n1156 GND.n1155 0.0815811
R4833 GND.n1173 GND.n1159 0.0815811
R4834 GND.n1070 GND 0.0807365
R4835 GND.n1079 GND 0.0807365
R4836 GND.n1824 GND.n1823 0.077375
R4837 GND.n600 GND.n598 0.0760208
R4838 GND.n706 GND.n705 0.0760208
R4839 GND.n631 GND.n630 0.0760208
R4840 GND.n645 GND.n644 0.0760208
R4841 GND.n659 GND.n651 0.0760208
R4842 GND.n687 GND.n686 0.0760208
R4843 GND.n1844 GND.n3 0.072593
R4844 GND.n54 GND.n4 0.072593
R4845 GND GND.n719 0.0603958
R4846 GND.n714 GND 0.0603958
R4847 GND.n707 GND 0.0603958
R4848 GND.n701 GND 0.0603958
R4849 GND.n629 GND 0.0603958
R4850 GND GND.n626 0.0603958
R4851 GND.n643 GND 0.0603958
R4852 GND.n649 GND 0.0603958
R4853 GND GND.n660 0.0603958
R4854 GND GND.n655 0.0603958
R4855 GND.n688 GND 0.0603958
R4856 GND.n525 GND 0.0603958
R4857 GND.n520 GND 0.0603958
R4858 GND.n500 GND 0.0603958
R4859 GND.n513 GND 0.0603958
R4860 GND.n508 GND 0.0603958
R4861 GND GND.n504 0.0603958
R4862 GND.n1321 GND 0.0603958
R4863 GND GND.n383 0.0603958
R4864 GND.n1281 GND 0.0603958
R4865 GND.n1282 GND 0.0603958
R4866 GND GND.n379 0.0603958
R4867 GND.n1286 GND 0.0603958
R4868 GND.n1290 GND 0.0603958
R4869 GND.n1291 GND 0.0603958
R4870 GND.n1292 GND 0.0603958
R4871 GND.n1295 GND 0.0603958
R4872 GND GND.n375 0.0603958
R4873 GND.n1302 GND 0.0603958
R4874 GND.n1303 GND 0.0603958
R4875 GND GND.n371 0.0603958
R4876 GND.n1313 GND 0.0603958
R4877 GND.n1222 GND 0.0603958
R4878 GND GND.n1220 0.0603958
R4879 GND.n1266 GND 0.0603958
R4880 GND GND.n1265 0.0603958
R4881 GND GND.n1264 0.0603958
R4882 GND GND.n1259 0.0603958
R4883 GND GND.n1258 0.0603958
R4884 GND.n1236 GND 0.0603958
R4885 GND.n1253 GND 0.0603958
R4886 GND GND.n1252 0.0603958
R4887 GND GND.n1251 0.0603958
R4888 GND.n1247 GND 0.0603958
R4889 GND GND.n1246 0.0603958
R4890 GND.n1242 GND 0.0603958
R4891 GND GND.n1241 0.0603958
R4892 GND.n57 GND.n56 0.0591735
R4893 GND.n52 GND.n1 0.0591735
R4894 GND.n729 GND.n728 0.058
R4895 GND.n730 GND.n729 0.058
R4896 GND.n734 GND.n576 0.058
R4897 GND.n735 GND.n734 0.058
R4898 GND.n740 GND.n739 0.058
R4899 GND.n741 GND.n740 0.058
R4900 GND.n745 GND.n572 0.058
R4901 GND.n746 GND.n745 0.058
R4902 GND.n751 GND.n750 0.058
R4903 GND.n752 GND.n751 0.058
R4904 GND.n756 GND.n568 0.058
R4905 GND.n757 GND.n756 0.058
R4906 GND.n762 GND.n761 0.058
R4907 GND.n763 GND.n762 0.058
R4908 GND.n767 GND.n564 0.058
R4909 GND.n768 GND.n767 0.058
R4910 GND.n773 GND.n772 0.058
R4911 GND.n774 GND.n773 0.058
R4912 GND.n778 GND.n560 0.058
R4913 GND.n779 GND.n778 0.058
R4914 GND.n784 GND.n783 0.058
R4915 GND.n785 GND.n784 0.058
R4916 GND.n789 GND.n556 0.058
R4917 GND.n790 GND.n789 0.058
R4918 GND.n795 GND.n794 0.058
R4919 GND.n796 GND.n795 0.058
R4920 GND.n800 GND.n552 0.058
R4921 GND.n801 GND.n800 0.058
R4922 GND.n806 GND.n805 0.058
R4923 GND.n807 GND.n806 0.058
R4924 GND.n811 GND.n548 0.058
R4925 GND.n812 GND.n811 0.058
R4926 GND.n817 GND.n816 0.058
R4927 GND.n818 GND.n817 0.058
R4928 GND.n822 GND.n544 0.058
R4929 GND.n823 GND.n822 0.058
R4930 GND.n828 GND.n541 0.058
R4931 GND.n829 GND.n828 0.058
R4932 GND.n830 GND.n539 0.058
R4933 GND.n834 GND.n539 0.058
R4934 GND.n681 GND 0.0577917
R4935 GND.n1064 GND.n1063 0.0553986
R4936 GND.n1073 GND.n1072 0.0553986
R4937 GND.n1082 GND.n1081 0.0553986
R4938 GND.n870 GND.n869 0.0553986
R4939 GND.n880 GND.n879 0.0553986
R4940 GND.n890 GND.n885 0.0553986
R4941 GND.n1017 GND.n895 0.0553986
R4942 GND.n902 GND.n901 0.0553986
R4943 GND.n912 GND.n911 0.0553986
R4944 GND.n922 GND.n917 0.0553986
R4945 GND.n989 GND.n927 0.0553986
R4946 GND.n934 GND.n933 0.0553986
R4947 GND.n944 GND.n943 0.0553986
R4948 GND.n953 GND.n949 0.0553986
R4949 GND.n961 GND.n958 0.0553986
R4950 GND.n402 GND.n397 0.0553986
R4951 GND.n1202 GND.n407 0.0553986
R4952 GND.n1191 GND.n412 0.0553986
R4953 GND.n1152 GND.n1151 0.0553986
R4954 GND.n1176 GND.n1158 0.0553986
R4955 GND.n1164 GND.n1161 0.0553986
R4956 GND.n1055 GND.n1054 0.0545423
R4957 GND.t636 GND.n1122 0.0500323
R4958 GND.n56 GND.n55 0.0489694
R4959 GND.n53 GND.n52 0.0489694
R4960 GND.n601 GND.n600 0.0447708
R4961 GND.n707 GND.n706 0.0447708
R4962 GND.n632 GND.n631 0.0447708
R4963 GND.n644 GND.n643 0.0447708
R4964 GND.n656 GND.n651 0.0447708
R4965 GND.n688 GND.n687 0.0447708
R4966 GND GND.n1060 0.0410405
R4967 GND GND.n1069 0.0410405
R4968 GND GND.n1078 0.0410405
R4969 GND GND.n1094 0.0410405
R4970 GND.n873 GND 0.0410405
R4971 GND.n893 GND 0.0410405
R4972 GND.n905 GND 0.0410405
R4973 GND.n925 GND 0.0410405
R4974 GND.n937 GND 0.0410405
R4975 GND.n956 GND 0.0410405
R4976 GND.n405 GND 0.0410405
R4977 GND GND.n1824 0.0390417
R4978 GND.n1677 GND.n1622 0.038
R4979 GND.n1694 GND.n1693 0.038
R4980 GND GND.n872 0.0351284
R4981 GND GND.n892 0.0351284
R4982 GND GND.n904 0.0351284
R4983 GND GND.n924 0.0351284
R4984 GND GND.n936 0.0351284
R4985 GND GND.n955 0.0351284
R4986 GND GND.n404 0.0351284
R4987 GND.n1190 GND 0.0351284
R4988 GND GND.n1154 0.0351284
R4989 GND.n1175 GND 0.0351284
R4990 GND.n1163 GND 0.0351284
R4991 GND.n712 GND 0.0343542
R4992 GND.n638 GND 0.0343542
R4993 GND.n693 GND 0.0343542
R4994 GND GND.n1291 0.0343542
R4995 GND.n1783 GND.n146 0.03425
R4996 GND GND.n500 0.0330521
R4997 GND.n504 GND 0.0330521
R4998 GND GND.n1321 0.0330521
R4999 GND.n1273 GND 0.0330521
R5000 GND GND.n1281 0.0330521
R5001 GND.n1282 GND 0.0330521
R5002 GND GND.n1302 0.0330521
R5003 GND.n1313 GND 0.0330521
R5004 GND.n1271 GND 0.0330521
R5005 GND.n1266 GND 0.0330521
R5006 GND.n1258 GND 0.0330521
R5007 GND.n1253 GND 0.0330521
R5008 GND.n1241 GND 0.0330521
R5009 GND.n728 GND 0.02925
R5010 GND GND.n576 0.02925
R5011 GND.n736 GND 0.02925
R5012 GND.n739 GND 0.02925
R5013 GND GND.n572 0.02925
R5014 GND.n747 GND 0.02925
R5015 GND.n750 GND 0.02925
R5016 GND GND.n568 0.02925
R5017 GND.n758 GND 0.02925
R5018 GND.n761 GND 0.02925
R5019 GND GND.n564 0.02925
R5020 GND.n769 GND 0.02925
R5021 GND.n772 GND 0.02925
R5022 GND GND.n560 0.02925
R5023 GND.n780 GND 0.02925
R5024 GND.n783 GND 0.02925
R5025 GND GND.n556 0.02925
R5026 GND.n791 GND 0.02925
R5027 GND.n794 GND 0.02925
R5028 GND GND.n552 0.02925
R5029 GND.n802 GND 0.02925
R5030 GND.n805 GND 0.02925
R5031 GND GND.n548 0.02925
R5032 GND.n813 GND 0.02925
R5033 GND.n816 GND 0.02925
R5034 GND GND.n544 0.02925
R5035 GND.n824 GND 0.02925
R5036 GND GND.n541 0.02925
R5037 GND.n830 GND 0.02925
R5038 GND.n1429 GND 0.0270625
R5039 GND.n1063 GND.n1053 0.0266824
R5040 GND.n1072 GND.n1052 0.0266824
R5041 GND.n1081 GND.n1042 0.0266824
R5042 GND.n870 GND.n864 0.0266824
R5043 GND.n880 GND.n874 0.0266824
R5044 GND.n890 GND.n884 0.0266824
R5045 GND.n895 GND.n894 0.0266824
R5046 GND.n902 GND.n896 0.0266824
R5047 GND.n912 GND.n906 0.0266824
R5048 GND.n922 GND.n916 0.0266824
R5049 GND.n927 GND.n926 0.0266824
R5050 GND.n934 GND.n928 0.0266824
R5051 GND.n944 GND.n938 0.0266824
R5052 GND.n953 GND.n948 0.0266824
R5053 GND.n958 GND.n957 0.0266824
R5054 GND.n402 GND.n396 0.0266824
R5055 GND.n407 GND.n406 0.0266824
R5056 GND.n412 GND.n408 0.0266824
R5057 GND.n1152 GND.n413 0.0266824
R5058 GND.n1158 GND.n1156 0.0266824
R5059 GND.n1161 GND.n1159 0.0266824
R5060 GND GND.n365 0.026141
R5061 GND GND.n882 0.0249932
R5062 GND.n1016 GND 0.0249932
R5063 GND GND.n914 0.0249932
R5064 GND.n988 GND 0.0249932
R5065 GND GND.n946 0.0249932
R5066 GND.n960 GND 0.0249932
R5067 GND.n1201 GND 0.0249932
R5068 GND GND.n601 0.0239375
R5069 GND GND.n605 0.0239375
R5070 GND.n704 GND 0.0239375
R5071 GND.n701 GND 0.0239375
R5072 GND.n700 GND 0.0239375
R5073 GND.n632 GND 0.0239375
R5074 GND.n624 GND 0.0239375
R5075 GND.n646 GND 0.0239375
R5076 GND GND.n649 0.0239375
R5077 GND.n661 GND 0.0239375
R5078 GND.n656 GND 0.0239375
R5079 GND GND.n617 0.0239375
R5080 GND.n685 GND 0.0239375
R5081 GND.n682 GND 0.0239375
R5082 GND.n511 GND 0.0239375
R5083 GND.n506 GND 0.0239375
R5084 GND.n379 GND 0.0239375
R5085 GND GND.n1290 0.0239375
R5086 GND.n1292 GND 0.0239375
R5087 GND.n372 GND 0.0239375
R5088 GND GND.n1236 0.0239375
R5089 GND.n1252 GND 0.0239375
R5090 GND GND.n1237 0.0239375
R5091 GND.n1247 GND 0.0239375
R5092 GND.n1245 GND 0.0239375
R5093 GND.n1242 GND 0.0239375
R5094 GND.n523 GND 0.0226354
R5095 GND.n1287 GND 0.0226354
R5096 GND.n1296 GND 0.0226354
R5097 GND GND.n1231 0.0226354
R5098 GND.n720 GND 0.0213333
R5099 GND.n528 GND 0.0213333
R5100 GND GND.n499 0.0213333
R5101 GND GND.n1280 0.0213333
R5102 GND GND.n1301 0.0213333
R5103 GND GND.n1311 0.0213333
R5104 GND.n1265 GND 0.0213333
R5105 GND.n1260 GND 0.0213333
R5106 GND.n1259 GND 0.0213333
R5107 GND.n712 GND 0.0194732
R5108 GND.n638 GND 0.0194732
R5109 GND GND.n693 0.0194732
R5110 GND.n1225 GND 0.016125
R5111 GND.n725 GND 0.016125
R5112 GND.n736 GND 0.016125
R5113 GND.n747 GND 0.016125
R5114 GND.n758 GND 0.016125
R5115 GND.n769 GND 0.016125
R5116 GND.n780 GND 0.016125
R5117 GND.n791 GND 0.016125
R5118 GND.n802 GND 0.016125
R5119 GND.n813 GND 0.016125
R5120 GND.n824 GND 0.016125
R5121 GND.n538 GND 0.0148229
R5122 GND.n1747 GND.n1746 0.0144752
R5123 GND.n1099 GND.n1096 0.01175
R5124 GND.n1440 GND.n283 0.011346
R5125 GND.n730 GND 0.011125
R5126 GND GND.n735 0.011125
R5127 GND.n741 GND 0.011125
R5128 GND GND.n746 0.011125
R5129 GND.n752 GND 0.011125
R5130 GND GND.n757 0.011125
R5131 GND.n763 GND 0.011125
R5132 GND GND.n768 0.011125
R5133 GND.n774 GND 0.011125
R5134 GND GND.n779 0.011125
R5135 GND.n785 GND 0.011125
R5136 GND GND.n790 0.011125
R5137 GND.n796 GND 0.011125
R5138 GND GND.n801 0.011125
R5139 GND.n807 GND 0.011125
R5140 GND GND.n812 0.011125
R5141 GND.n818 GND 0.011125
R5142 GND GND.n823 0.011125
R5143 GND GND.n829 0.011125
R5144 GND GND.n834 0.011125
R5145 GND.n1839 GND.n1838 0.009875
R5146 GND.n1838 GND.n51 0.00912069
R5147 GND.n39 GND.n38 0.00912069
R5148 GND.n1440 GND.n1439 0.00646529
R5149 GND.n1064 GND.n1061 0.00641216
R5150 GND.n1073 GND.n1070 0.00641216
R5151 GND.n1082 GND.n1079 0.00641216
R5152 GND.n872 GND.n869 0.00641216
R5153 GND.n882 GND.n879 0.00641216
R5154 GND.n892 GND.n885 0.00641216
R5155 GND.n1017 GND.n1016 0.00641216
R5156 GND.n904 GND.n901 0.00641216
R5157 GND.n914 GND.n911 0.00641216
R5158 GND.n924 GND.n917 0.00641216
R5159 GND.n989 GND.n988 0.00641216
R5160 GND.n936 GND.n933 0.00641216
R5161 GND.n946 GND.n943 0.00641216
R5162 GND.n955 GND.n949 0.00641216
R5163 GND.n961 GND.n960 0.00641216
R5164 GND.n404 GND.n397 0.00641216
R5165 GND.n1202 GND.n1201 0.00641216
R5166 GND.n1191 GND.n1190 0.00641216
R5167 GND.n1154 GND.n1151 0.00641216
R5168 GND.n1176 GND.n1175 0.00641216
R5169 GND.n1164 GND.n1163 0.00641216
R5170 GND.n1824 GND.n146 0.00425
R5171 GND.n682 GND.n681 0.00310417
R5172 a_45343_4538.t0 a_45343_4538.t1 49.8467
R5173 top_DAC_0/top_final_switch_0.VOUT[1].n2 top_DAC_0/top_final_switch_0.VOUT[1].n0 603.66
R5174 top_DAC_0/top_final_switch_0.VOUT[1].n2 top_DAC_0/top_final_switch_0.VOUT[1].n1 202.21
R5175 top_DAC_0/top_final_switch_0.VOUT[1].n3 top_DAC_0/top_final_switch_0.VOUT[1].t9 172.237
R5176 top_DAC_0/top_final_switch_0.VOUT[1].n4 top_DAC_0/top_final_switch_0.VOUT[1].t5 171.161
R5177 top_DAC_0/top_final_switch_0.VOUT[1].n3 top_DAC_0/top_final_switch_0.VOUT[1].t7 170.625
R5178 top_DAC_0/top_final_switch_0.VOUT[1].n4 top_DAC_0/top_final_switch_0.VOUT[1].t11 170.625
R5179 top_DAC_0/top_final_switch_0.VOUT[1].n7 top_DAC_0/top_final_switch_0.VOUT[1].t8 121.868
R5180 top_DAC_0/top_final_switch_0.VOUT[1].n6 top_DAC_0/top_final_switch_0.VOUT[1].t4 120.793
R5181 top_DAC_0/top_final_switch_0.VOUT[1].n7 top_DAC_0/top_final_switch_0.VOUT[1].t6 120.255
R5182 top_DAC_0/top_final_switch_0.VOUT[1].n6 top_DAC_0/top_final_switch_0.VOUT[1].t10 120.255
R5183 top_DAC_0/top_final_switch_0.VOUT[1].n0 top_DAC_0/top_final_switch_0.VOUT[1].t2 65.941
R5184 top_DAC_0/top_final_switch_0.VOUT[1].n0 top_DAC_0/top_final_switch_0.VOUT[1].t3 65.941
R5185 top_DAC_0/top_final_switch_0.VOUT[1].n1 top_DAC_0/top_final_switch_0.VOUT[1].t0 39.3576
R5186 top_DAC_0/top_final_switch_0.VOUT[1].n1 top_DAC_0/top_final_switch_0.VOUT[1].t1 39.3576
R5187 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_final_switch_0.VOUT[1].n9 15.238
R5188 top_DAC_0/top_final_switch_0.VOUT[1].n5 top_DAC_0/top_final_switch_0.VOUT[1].n3 8.69842
R5189 top_DAC_0/top_final_switch_0.VOUT[1].n8 top_DAC_0/top_final_switch_0.VOUT[1].n6 7.53592
R5190 top_DAC_0/top_final_switch_0.VOUT[1].n10 top_DAC_0/top_final_switch_0.VOUT[1] 5.89065
R5191 top_DAC_0/top_final_switch_0.VOUT[1].n5 top_DAC_0/top_final_switch_0.VOUT[1].n4 5.82758
R5192 top_DAC_0/top_final_switch_0.VOUT[1].n8 top_DAC_0/top_final_switch_0.VOUT[1].n7 5.29008
R5193 top_DAC_0/top_final_switch_0.VOUT[1].n9 top_DAC_0/top_final_switch_0.VOUT[1].n5 1.13383
R5194 top_DAC_0/top_final_switch_0.VOUT[1].n9 top_DAC_0/top_final_switch_0.VOUT[1].n8 0.583833
R5195 top_DAC_0/top_final_switch_0.VOUT[1].n10 top_DAC_0/top_final_switch_0.VOUT[1].n2 0.233364
R5196 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_final_switch_0.VOUT[1].n10 0.0275606
R5197 a_6778_12595.n3 a_6778_12595.t6 236.924
R5198 a_6778_12595.n3 a_6778_12595.t9 235.214
R5199 a_6778_12595.n6 a_6778_12595.n5 71.3963
R5200 a_6778_12595.n2 a_6778_12595.n1 71.3963
R5201 a_6778_12595.n2 a_6778_12595.n0 71.3963
R5202 a_6778_12595.n7 a_6778_12595.n6 71.3963
R5203 a_6778_12595.n5 a_6778_12595.t1 16.5305
R5204 a_6778_12595.n5 a_6778_12595.t5 16.5305
R5205 a_6778_12595.n1 a_6778_12595.t3 16.5305
R5206 a_6778_12595.n1 a_6778_12595.t8 16.5305
R5207 a_6778_12595.n0 a_6778_12595.t7 16.5305
R5208 a_6778_12595.n0 a_6778_12595.t4 16.5305
R5209 a_6778_12595.n7 a_6778_12595.t2 16.5305
R5210 a_6778_12595.t0 a_6778_12595.n7 16.5305
R5211 a_6778_12595.n4 a_6778_12595.n3 4.7735
R5212 a_6778_12595.n6 a_6778_12595.n4 0.3505
R5213 a_6778_12595.n4 a_6778_12595.n2 0.3505
R5214 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t17 84.1846
R5215 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t5 83.2221
R5216 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t20 83.2221
R5217 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t21 83.2221
R5218 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t4 83.2221
R5219 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t1 83.2221
R5220 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t18 83.2221
R5221 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t2 83.2221
R5222 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t10 83.2221
R5223 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t14 83.2221
R5224 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n1 66.665
R5225 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n0 66.665
R5226 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n39 66.665
R5227 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n38 66.665
R5228 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n35 66.665
R5229 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t13 60.0431
R5230 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t12 55.7878
R5231 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t7 55.5545
R5232 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t8 49.6518
R5233 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n4 18.1401
R5234 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n23 16.8247
R5235 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t22 16.5305
R5236 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t23 16.5305
R5237 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t3 16.5305
R5238 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t6 16.5305
R5239 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t16 16.5305
R5240 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t19 16.5305
R5241 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t11 16.5305
R5242 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t9 16.5305
R5243 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t15 16.5305
R5244 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t0 16.5305
R5245 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n26 10.2109
R5246 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n30 10.2109
R5247 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n34 10.2109
R5248 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n40 10.2089
R5249 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n44 10.2089
R5250 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n24 7.49008
R5251 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n3 7.44425
R5252 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n2 7.39008
R5253 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 7.00883
R5254 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n28 6.00467
R5255 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n32 6.00467
R5256 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n42 6.00467
R5257 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n37 6.00467
R5258 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n25 4.5005
R5259 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n29 4.5005
R5260 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n33 4.5005
R5261 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n41 4.5005
R5262 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n45 4.5005
R5263 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n7 3.90596
R5264 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n18 3.90547
R5265 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n21 3.4105
R5266 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n14 3.4105
R5267 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n10 3.4105
R5268 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n27 0.962993
R5269 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n31 0.962993
R5270 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n43 0.962974
R5271 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n36 0.962974
R5272 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t41 0.523604
R5273 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t38 0.523604
R5274 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t30 0.523604
R5275 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t27 0.523604
R5276 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t24 0.523604
R5277 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n11 0.495958
R5278 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t42 0.402677
R5279 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t39 0.402677
R5280 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t31 0.402677
R5281 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t28 0.402677
R5282 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t25 0.402677
R5283 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n15 0.319708
R5284 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t35 0.28175
R5285 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t29 0.28175
R5286 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t33 0.28175
R5287 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t26 0.28175
R5288 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t43 0.28175
R5289 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t36 0.28175
R5290 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t40 0.28175
R5291 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t34 0.28175
R5292 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t37 0.28175
R5293 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t32 0.28175
R5294 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n5 0.242354
R5295 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n8 0.242354
R5296 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n12 0.242354
R5297 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n19 0.242354
R5298 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n16 0.242354
R5299 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n22 0.17724
R5300 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n6 0.121427
R5301 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n9 0.121427
R5302 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n13 0.121427
R5303 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n20 0.121427
R5304 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n17 0.121427
R5305 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.04425
R5306 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.04425
R5307 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.04425
R5308 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.04425
R5309 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n46 0.04425
R5310 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t1 334.771
R5311 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t18 213.218
R5312 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t14 213.218
R5313 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t5 213.218
R5314 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t22 212.895
R5315 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t23 212.554
R5316 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t2 212.554
R5317 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t3 212.554
R5318 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t20 212.554
R5319 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t17 212.554
R5320 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t16 212.554
R5321 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t21 212.554
R5322 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t12 212.554
R5323 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t9 212.554
R5324 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t15 212.554
R5325 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t4 212.554
R5326 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t10 212.554
R5327 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t8 212.554
R5328 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t6 208.054
R5329 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n21 152
R5330 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t7 126.278
R5331 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t19 125.566
R5332 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t11 125.566
R5333 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t13 114.031
R5334 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t0 87.8568
R5335 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t24 81.5883
R5336 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n20 43.6567
R5337 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n4 20.963
R5338 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n19 19.2422
R5339 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 15.6308
R5340 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n22 11.4706
R5341 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 7.31717
R5342 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n11 7.0755
R5343 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n3 5.04008
R5344 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 4.82262
R5345 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n2 4.68383
R5346 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 4.48881
R5347 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n23 1.01508
R5348 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n0 0.876942
R5349 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.7755
R5350 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n1 0.713
R5351 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n12 0.663962
R5352 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n13 0.663962
R5353 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n14 0.663962
R5354 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n15 0.663962
R5355 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n16 0.663962
R5356 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n17 0.663962
R5357 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n9 0.663962
R5358 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n8 0.663962
R5359 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n5 0.663962
R5360 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n6 0.663962
R5361 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n10 0.312199
R5362 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n7 0.312199
R5363 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n18 0.254667
R5364 a_30056_7686.n0 a_30056_7686.t3 246.061
R5365 a_30056_7686.t0 a_30056_7686.n2 240.989
R5366 a_30056_7686.n2 a_30056_7686.t2 240.81
R5367 a_30056_7686.n0 a_30056_7686.t1 238.775
R5368 a_30056_7686.n1 a_30056_7686.t4 238.775
R5369 a_30056_7686.n1 a_30056_7686.n0 6.788
R5370 a_30056_7686.n2 a_30056_7686.n1 4.54842
R5371 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.t1 249.345
R5372 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.t0 10.5773
R5373 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.t2 10.5739
R5374 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.n0 4.18158
R5375 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t4 221.851
R5376 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t2 221.851
R5377 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t5 140.244
R5378 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t0 140.056
R5379 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t18 122.656
R5380 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t9 122.656
R5381 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t17 122.656
R5382 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t8 122.656
R5383 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t11 122.656
R5384 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t15 122.656
R5385 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t16 122.656
R5386 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t6 122.656
R5387 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t10 122.656
R5388 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t13 122.656
R5389 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t7 122.656
R5390 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t14 122.656
R5391 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t3 108.365
R5392 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t1 108.365
R5393 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n17 14.4346
R5394 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t12 13.3032
R5395 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n18 12.8291
R5396 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n2 11.1702
R5397 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n20 4.63108
R5398 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n0 3.9493
R5399 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n19 3.4105
R5400 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n21 2.67342
R5401 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n4 2.26409
R5402 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n1 2.25675
R5403 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n5 0.742167
R5404 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n6 0.742167
R5405 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n7 0.742167
R5406 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n15 0.742167
R5407 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n14 0.742167
R5408 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n13 0.742167
R5409 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n11 0.742167
R5410 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n10 0.742167
R5411 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n9 0.742167
R5412 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n16 0.652583
R5413 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n12 0.652583
R5414 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n1 0.546515
R5415 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n3 0.527402
R5416 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.504667
R5417 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.0900833
R5418 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.0900833
R5419 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.0650833
R5420 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n22 0.063
R5421 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.0498421
R5422 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n8 0.0255
R5423 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t1 334.771
R5424 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t9 213.218
R5425 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t6 213.218
R5426 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t3 212.554
R5427 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t2 212.554
R5428 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t4 208.054
R5429 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t5 126.278
R5430 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t7 125.566
R5431 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t8 125.566
R5432 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t0 87.8568
R5433 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n3 65.2609
R5434 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n7 5.04008
R5435 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n6 4.68383
R5436 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n2 4.5005
R5437 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n4 0.876942
R5438 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n5 0.713
R5439 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n1 0.663962
R5440 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n0 0.363481
R5441 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.300981
R5442 a_44062_19517.t0 a_44062_19517.t1 129.28
R5443 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n1 863.124
R5444 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n0 585
R5445 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t0 495.469
R5446 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t15 217.555
R5447 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t10 217.555
R5448 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t12 216.893
R5449 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t11 216.893
R5450 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t8 216.893
R5451 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t6 216.893
R5452 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t4 216.893
R5453 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t9 216.893
R5454 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t7 216.893
R5455 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t5 216.893
R5456 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t3 216.893
R5457 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t2 216.893
R5458 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t16 216.893
R5459 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t14 216.893
R5460 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t13 216.893
R5461 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t17 216.893
R5462 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t1 141.189
R5463 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t0 140.738
R5464 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n18 101.117
R5465 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n19 13.9797
R5466 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n10 12.8332
R5467 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 11.6369
R5468 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 10.1408
R5469 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n20 8.14595
R5470 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n3 7.94225
R5471 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 6.20656
R5472 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 6.14988
R5473 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 2.16154
R5474 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec2b[0] 0.7755
R5475 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n2 0.665435
R5476 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n8 0.663962
R5477 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n7 0.663962
R5478 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n4 0.663962
R5479 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n5 0.663962
R5480 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n17 0.663962
R5481 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n16 0.663962
R5482 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n15 0.663962
R5483 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n14 0.663962
R5484 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n13 0.663962
R5485 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n12 0.663962
R5486 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n11 0.663962
R5487 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n9 0.320692
R5488 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n6 0.320692
R5489 a_14331_6250.n2 a_14331_6250.t4 672.461
R5490 a_14331_6250.n0 a_14331_6250.t3 672.087
R5491 a_14331_6250.n1 a_14331_6250.t1 671.755
R5492 a_14331_6250.n0 a_14331_6250.t2 665.667
R5493 a_14331_6250.t0 a_14331_6250.n2 665.667
R5494 a_14331_6250.n2 a_14331_6250.n1 5.39008
R5495 a_14331_6250.n1 a_14331_6250.n0 1.17133
R5496 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t1 673.192
R5497 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t2 10.7568
R5498 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t0 10.6545
R5499 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.n0 0.67884
R5500 VDDH.n398 VDDH.n397 10828.8
R5501 VDDH.n399 VDDH.n398 10828.8
R5502 VDDH.n535 VDDH.n185 10344.7
R5503 VDDH.n254 VDDH.n185 10344.7
R5504 VDDH.n577 VDDH.n178 9916.1
R5505 VDDH.n196 VDDH.n180 9916.1
R5506 VDDH.n530 VDDH.n178 9914.2
R5507 VDDH.n446 VDDH.n196 9914.2
R5508 VDDH.n573 VDDH.n187 9786.51
R5509 VDDH.n573 VDDH.n188 9786.51
R5510 VDDH.n526 VDDH.n179 8757.1
R5511 VDDH.n526 VDDH.n447 8755.2
R5512 VDDH.n285 VDDH.n184 8715.3
R5513 VDDH.n228 VDDH.n184 8715.3
R5514 VDDH.n253 VDDH.n186 8715.3
R5515 VDDH.n532 VDDH.n186 8715.3
R5516 VDDH.n252 VDDH.n183 8715.3
R5517 VDDH.n444 VDDH.n183 8715.3
R5518 VDDH.n392 VDDH.n189 7193.6
R5519 VDDH.n393 VDDH.n392 7193.6
R5520 VDDH.n143 VDDH.n141 5941.3
R5521 VDDH.n143 VDDH.n94 5941.3
R5522 VDDH.n166 VDDH.n141 5939.4
R5523 VDDH.n111 VDDH.n109 5352.3
R5524 VDDH.n1050 VDDH.n1046 4436.17
R5525 VDDH.n1050 VDDH.n1047 4436.17
R5526 VDDH.n1052 VDDH.n1046 4436.17
R5527 VDDH.n1052 VDDH.n1047 4436.17
R5528 VDDH.n153 VDDH.n152 4157.2
R5529 VDDH.n490 VDDH.n464 4035.6
R5530 VDDH.n507 VDDH.n464 4035.6
R5531 VDDH.n510 VDDH.n457 3731.6
R5532 VDDH.n510 VDDH.n509 3731.6
R5533 VDDH.n163 VDDH.n122 3638.5
R5534 VDDH.n671 VDDH.n122 3638.5
R5535 VDDH.n283 VDDH.n255 3420
R5536 VDDH.n283 VDDH.n256 3420
R5537 VDDH.n441 VDDH.n229 3420
R5538 VDDH.n441 VDDH.n230 3420
R5539 VDDH.n643 VDDH.n618 3298.14
R5540 VDDH.n646 VDDH.n618 3296.17
R5541 VDDH.n416 VDDH.n413 2996.3
R5542 VDDH.n418 VDDH.n413 2996.3
R5543 VDDH.n418 VDDH.n415 2996.3
R5544 VDDH.n416 VDDH.n415 2996.3
R5545 VDDH.n646 VDDH.n619 2942.38
R5546 VDDH.n653 VDDH.n611 2942.38
R5547 VDDH.n655 VDDH.n606 2942.38
R5548 VDDH.n656 VDDH.n606 2942.38
R5549 VDDH.n652 VDDH.n611 2942.38
R5550 VDDH.n643 VDDH.n620 2940.41
R5551 VDDH.n152 VDDH.n151 2855.7
R5552 VDDH.n715 VDDH.n714 2705.6
R5553 VDDH.n674 VDDH.n120 2692.3
R5554 VDDH.n1134 VDDH.n995 2671.14
R5555 VDDH.n1136 VDDH.n995 2671.14
R5556 VDDH.n1136 VDDH.n1133 2671.14
R5557 VDDH.n1134 VDDH.n1133 2671.14
R5558 VDDH.n1058 VDDH.n1030 2671.14
R5559 VDDH.n1058 VDDH.n1031 2671.14
R5560 VDDH.n1060 VDDH.n1030 2671.14
R5561 VDDH.n1060 VDDH.n1031 2671.14
R5562 VDDH.n1039 VDDH.n1035 2671.14
R5563 VDDH.n1041 VDDH.n1035 2671.14
R5564 VDDH.n1041 VDDH.n1037 2671.14
R5565 VDDH.n1039 VDDH.n1037 2671.14
R5566 VDDH.n1125 VDDH.n1000 2671.14
R5567 VDDH.n1125 VDDH.n1001 2671.14
R5568 VDDH.n1127 VDDH.n1000 2671.14
R5569 VDDH.n1127 VDDH.n1001 2671.14
R5570 VDDH.n1118 VDDH.n1005 2671.14
R5571 VDDH.n1118 VDDH.n1006 2671.14
R5572 VDDH.n1116 VDDH.n1006 2671.14
R5573 VDDH.n1116 VDDH.n1005 2671.14
R5574 VDDH.n1071 VDDH.n1065 2671.14
R5575 VDDH.n1071 VDDH.n1067 2671.14
R5576 VDDH.n1069 VDDH.n1067 2671.14
R5577 VDDH.n1069 VDDH.n1065 2671.14
R5578 VDDH.n1078 VDDH.n1024 2671.14
R5579 VDDH.n1078 VDDH.n1025 2671.14
R5580 VDDH.n1080 VDDH.n1025 2671.14
R5581 VDDH.n1080 VDDH.n1024 2671.14
R5582 VDDH.n1111 VDDH.n1011 2671.14
R5583 VDDH.n1111 VDDH.n1012 2671.14
R5584 VDDH.n1109 VDDH.n1012 2671.14
R5585 VDDH.n1109 VDDH.n1011 2671.14
R5586 VDDH.n1100 VDDH.n1016 2671.14
R5587 VDDH.n1100 VDDH.n1017 2671.14
R5588 VDDH.n1102 VDDH.n1017 2671.14
R5589 VDDH.n1102 VDDH.n1016 2671.14
R5590 VDDH.n1091 VDDH.n1084 2671.14
R5591 VDDH.n1091 VDDH.n1085 2671.14
R5592 VDDH.n1089 VDDH.n1085 2671.14
R5593 VDDH.n1089 VDDH.n1084 2671.14
R5594 VDDH.n490 VDDH.n487 2612.5
R5595 VDDH.n468 VDDH.n463 2612.5
R5596 VDDH.n469 VDDH.n468 2612.5
R5597 VDDH.n507 VDDH.n469 2612.5
R5598 VDDH.n488 VDDH.n462 2612.5
R5599 VDDH.n488 VDDH.n487 2612.5
R5600 VDDH.n654 VDDH.n653 2588.59
R5601 VDDH.n655 VDDH.n654 2588.59
R5602 VDDH.n652 VDDH.n609 2588.59
R5603 VDDH.n656 VDDH.n609 2588.59
R5604 VDDH.n674 VDDH.n121 2513.7
R5605 VDDH.n592 VDDH.n591 2411.69
R5606 VDDH.n462 VDDH.n457 2308.5
R5607 VDDH.n509 VDDH.n463 2308.5
R5608 VDDH.n494 VDDH.n474 2283.8
R5609 VDDH.n495 VDDH.n474 2283.8
R5610 VDDH.n496 VDDH.n495 2283.8
R5611 VDDH.n496 VDDH.n494 2283.8
R5612 VDDH.n156 VDDH.n109 2129.9
R5613 VDDH.n159 VDDH.n156 2069.1
R5614 VDDH.n121 VDDH.n111 1983.6
R5615 VDDH.n579 VDDH.n176 1964.8
R5616 VDDH.n520 VDDH.n176 1964.42
R5617 VDDH.n569 VDDH.n568 1964.42
R5618 VDDH.n592 VDDH.n588 1934.07
R5619 VDDH.n572 VDDH.n190 1932.05
R5620 VDDH.n572 VDDH.n189 1931.86
R5621 VDDH.n762 VDDH.n744 1881
R5622 VDDH.n829 VDDH.n744 1881
R5623 VDDH.n829 VDDH.n41 1881
R5624 VDDH.n893 VDDH.n41 1881
R5625 VDDH.n894 VDDH.n893 1881
R5626 VDDH.n894 VDDH.n11 1881
R5627 VDDH.n973 VDDH.n11 1881
R5628 VDDH.n973 VDDH.n5 1881
R5629 VDDH.n977 VDDH.n5 1881
R5630 VDDH.n978 VDDH.n977 1881
R5631 VDDH.n634 VDDH.n628 1857.41
R5632 VDDH.n633 VDDH.n628 1857.41
R5633 VDDH.n591 VDDH.n584 1831.86
R5634 VDDH.n278 VDDH.n260 1778.4
R5635 VDDH.n278 VDDH.n261 1778.4
R5636 VDDH.n242 VDDH.n236 1778.4
R5637 VDDH.n242 VDDH.n234 1778.4
R5638 VDDH.n271 VDDH.n265 1778.4
R5639 VDDH.n271 VDDH.n269 1778.4
R5640 VDDH.n240 VDDH.n239 1778.4
R5641 VDDH.n239 VDDH.n235 1778.4
R5642 VDDH.n527 VDDH.n177 1735.15
R5643 VDDH.n528 VDDH.n527 1734.78
R5644 VDDH.n569 VDDH 1728.75
R5645 VDDH.n552 VDDH.n214 1726.87
R5646 VDDH.n538 VDDH.n537 1726.87
R5647 VDDH.n389 VDDH.n291 1726.87
R5648 VDDH.n248 VDDH.n214 1726.5
R5649 VDDH.n538 VDDH.n226 1726.49
R5650 VDDH.n391 VDDH.n389 1726.49
R5651 VDDH.n260 VDDH.n255 1641.6
R5652 VDDH.n275 VDDH.n260 1641.6
R5653 VDDH.n275 VDDH.n265 1641.6
R5654 VDDH.n265 VDDH.n264 1641.6
R5655 VDDH.n264 VDDH.n236 1641.6
R5656 VDDH.n434 VDDH.n236 1641.6
R5657 VDDH.n434 VDDH.n240 1641.6
R5658 VDDH.n240 VDDH.n229 1641.6
R5659 VDDH.n261 VDDH.n256 1641.6
R5660 VDDH.n263 VDDH.n261 1641.6
R5661 VDDH.n269 VDDH.n263 1641.6
R5662 VDDH.n269 VDDH.n268 1641.6
R5663 VDDH.n268 VDDH.n234 1641.6
R5664 VDDH.n436 VDDH.n234 1641.6
R5665 VDDH.n436 VDDH.n235 1641.6
R5666 VDDH.n235 VDDH.n230 1641.6
R5667 VDDH.n286 VDDH.n253 1629.41
R5668 VDDH.n533 VDDH.n532 1629.41
R5669 VDDH.n535 VDDH.n228 1578.31
R5670 VDDH.n286 VDDH.n285 1578.31
R5671 VDDH.n285 VDDH.n254 1578.31
R5672 VDDH.n533 VDDH.n228 1578.31
R5673 VDDH.n155 VDDH.n154 1506.3
R5674 VDDH.n638 VDDH.n619 1503.62
R5675 VDDH.n638 VDDH.n626 1503.62
R5676 VDDH.n634 VDDH.n626 1503.62
R5677 VDDH.n639 VDDH.n620 1503.62
R5678 VDDH.n639 VDDH.n623 1503.62
R5679 VDDH.n633 VDDH.n623 1503.62
R5680 VDDH.n487 VDDH.n465 1423.1
R5681 VDDH.n469 VDDH.n465 1423.1
R5682 VDDH.n512 VDDH.n462 1423.1
R5683 VDDH.n512 VDDH.n463 1423.1
R5684 VDDH.n596 VDDH.n588 1413.21
R5685 VDDH.n153 VDDH.n142 1407.9
R5686 VDDH.n696 VDDH.n93 1182.12
R5687 VDDH.n140 VDDH.n93 1182.12
R5688 VDDH.n167 VDDH.n140 1181.74
R5689 VDDH.n530 VDDH.n447 1109.6
R5690 VDDH.n577 VDDH.n179 1109.6
R5691 VDDH.n180 VDDH.n179 1109.6
R5692 VDDH.n447 VDDH.n446 1109.6
R5693 VDDH.n532 VDDH.n445 1071.21
R5694 VDDH.n288 VDDH.n253 1071.21
R5695 VDDH.n600 VDDH.n584 1027.97
R5696 VDDH.n445 VDDH.n444 1020.1
R5697 VDDH.n252 VDDH.n187 1020.1
R5698 VDDH.n288 VDDH.n252 1020.1
R5699 VDDH.n444 VDDH.n188 1020.1
R5700 VDDH.n163 VDDH.n120 986.101
R5701 VDDH.n671 VDDH.n121 986.101
R5702 VDDH.n1043 VDDH.n1032 883.577
R5703 VDDH.n1062 VDDH.n1028 883.577
R5704 VDDH.n1049 VDDH.n1033 854.212
R5705 VDDH.n1049 VDDH.n1048 854.212
R5706 VDDH.t141 VDDH.t457 824.275
R5707 VDDH.n695 VDDH.n694 823.718
R5708 VDDH.n1053 VDDH.n1045 781.929
R5709 VDDH.n1054 VDDH.n1053 781.929
R5710 VDDH.n589 VDDH.n586 772.448
R5711 VDDH.n443 VDDH.t82 759.42
R5712 VDDH.n492 VDDH.n491 756.33
R5713 VDDH.n466 VDDH.n456 744.283
R5714 VDDH.n515 VDDH.n456 744.283
R5715 VDDH.t382 VDDH.t425 740.356
R5716 VDDH.t456 VDDH.n181 734.784
R5717 VDDH.n687 VDDH.n686 725.46
R5718 VDDH.n669 VDDH.n668 720.942
R5719 VDDH.n668 VDDH.n123 720.942
R5720 VDDH.n154 VDDH.n153 720.101
R5721 VDDH.n282 VDDH.n281 682.542
R5722 VDDH.n440 VDDH.n439 682.542
R5723 VDDH.n992 VDDH.t64 667.769
R5724 VDDH.n642 VDDH.n616 636.236
R5725 VDDH.t83 VDDH.n575 630.073
R5726 VDDH.n414 VDDH.n412 598.588
R5727 VDDH.n423 VDDH.n412 598.588
R5728 VDDH.n422 VDDH.n414 598.588
R5729 VDDH.n423 VDDH.n422 598.588
R5730 VDDH.t515 VDDH.t497 583.548
R5731 VDDH.t506 VDDH.t331 583.548
R5732 VDDH.t514 VDDH.t334 583.548
R5733 VDDH.n659 VDDH.n605 568.095
R5734 VDDH.n695 VDDH.n95 564.33
R5735 VDDH.n647 VDDH.n617 563.577
R5736 VDDH.n642 VDDH.n641 563.201
R5737 VDDH.t521 VDDH.t575 552.236
R5738 VDDH.n712 VDDH.n90 536.095
R5739 VDDH.n716 VDDH.n90 536.095
R5740 VDDH.n675 VDDH.n119 533.46
R5741 VDDH.n506 VDDH.n505 528.759
R5742 VDDH.t503 VDDH.t459 523.162
R5743 VDDH.t351 VDDH.t373 523.162
R5744 VDDH.t561 VDDH.t38 523.162
R5745 VDDH.t451 VDDH.t339 523.162
R5746 VDDH.t374 VDDH.t537 523.162
R5747 VDDH.t244 VDDH.t81 523.162
R5748 VDDH.n596 VDDH.n586 522.828
R5749 VDDH.n514 VDDH.n458 522.542
R5750 VDDH.n486 VDDH.n458 522.542
R5751 VDDH.n506 VDDH.n471 522.542
R5752 VDDH.n491 VDDH.n486 522.542
R5753 VDDH.n470 VDDH.n461 522.542
R5754 VDDH.n471 VDDH.n470 522.542
R5755 VDDH.n1038 VDDH.n1034 516.141
R5756 VDDH.n1124 VDDH.n998 516.141
R5757 VDDH.n1077 VDDH.n1023 516.141
R5758 VDDH.n1081 VDDH.n1023 516.141
R5759 VDDH.n1088 VDDH.n1086 516.141
R5760 VDDH.n1138 VDDH.n994 516.141
R5761 VDDH.n1138 VDDH.n1137 516.141
R5762 VDDH.n156 VDDH.n98 513
R5763 VDDH.n154 VDDH.n98 511.101
R5764 VDDH.n231 VDDH.n227 507.824
R5765 VDDH.n8 VDDH.t504 499.882
R5766 VDDH.n9 VDDH.t516 499.882
R5767 VDDH.n10 VDDH.t573 499.882
R5768 VDDH.n980 VDDH.t332 499.882
R5769 VDDH.n614 VDDH.n613 495.812
R5770 VDDH.n613 VDDH.n605 495.812
R5771 VDDH.n651 VDDH.n650 495.812
R5772 VDDH.n651 VDDH.n608 495.812
R5773 VDDH.n657 VDDH.n608 495.812
R5774 VDDH.n658 VDDH.n657 495.812
R5775 VDDH VDDH.n614 490.166
R5776 VDDH.n155 VDDH.n151 489.267
R5777 VDDH.n676 VDDH.n110 486.776
R5778 VDDH.n159 VDDH.n155 486.401
R5779 VDDH.t250 VDDH.t308 475
R5780 VDDH.t249 VDDH.t458 475
R5781 VDDH.t522 VDDH.t350 475
R5782 VDDH.t330 VDDH.t312 475
R5783 VDDH.t312 VDDH.t530 475
R5784 VDDH.t379 VDDH.t240 475
R5785 VDDH.t405 VDDH.t375 475
R5786 VDDH.t396 VDDH.t408 475
R5787 VDDH.n593 VDDH.n583 466.447
R5788 VDDH.n466 VDDH.n461 462.307
R5789 VDDH.n515 VDDH.n514 462.307
R5790 VDDH.n503 VDDH.n475 457.413
R5791 VDDH.n497 VDDH.n475 457.413
R5792 VDDH.n600 VDDH.t563 455.01
R5793 VDDH.n1057 VDDH.n1032 443.86
R5794 VDDH.n1036 VDDH.n1026 443.86
R5795 VDDH.n1036 VDDH.n1028 443.86
R5796 VDDH.n1062 VDDH.n1061 443.86
R5797 VDDH.n1061 VDDH.n1003 443.86
R5798 VDDH.n1072 VDDH.n1064 443.86
R5799 VDDH.n1119 VDDH.n1004 443.86
R5800 VDDH.n1124 VDDH.n1123 443.86
R5801 VDDH.n1082 VDDH.n1081 443.86
R5802 VDDH.n1068 VDDH.n1021 443.86
R5803 VDDH.n1068 VDDH.n1018 443.86
R5804 VDDH.n1115 VDDH.n1008 443.86
R5805 VDDH.n1115 VDDH.n1114 443.86
R5806 VDDH.n1128 VDDH.n999 443.86
R5807 VDDH.n1129 VDDH.n1128 443.86
R5808 VDDH.n1088 VDDH.n1087 443.86
R5809 VDDH.n1103 VDDH.n1015 443.86
R5810 VDDH.n1104 VDDH.n1103 443.86
R5811 VDDH.n1108 VDDH.n1105 443.86
R5812 VDDH.n1108 VDDH.n1107 443.86
R5813 VDDH.n1137 VDDH.n996 443.86
R5814 VDDH.t476 VDDH.t483 431.25
R5815 VDDH.t480 VDDH.t476 431.25
R5816 VDDH.t479 VDDH.t480 431.25
R5817 VDDH.t477 VDDH.t491 431.25
R5818 VDDH.t491 VDDH.t490 431.25
R5819 VDDH.t490 VDDH.t478 431.25
R5820 VDDH.t307 VDDH.t311 431.25
R5821 VDDH.t378 VDDH.t307 431.25
R5822 VDDH.t308 VDDH.t378 431.25
R5823 VDDH.t248 VDDH.t250 431.25
R5824 VDDH.t247 VDDH.t248 431.25
R5825 VDDH.t458 VDDH.t522 431.25
R5826 VDDH.t350 VDDH.t330 431.25
R5827 VDDH.t377 VDDH.t342 431.25
R5828 VDDH.t344 VDDH.t377 431.25
R5829 VDDH.t343 VDDH.t344 431.25
R5830 VDDH.t415 VDDH.t416 431.25
R5831 VDDH.t416 VDDH.t376 431.25
R5832 VDDH.t376 VDDH.t414 431.25
R5833 VDDH.t450 VDDH.t243 431.25
R5834 VDDH.t448 VDDH.t450 431.25
R5835 VDDH.t242 VDDH.t448 431.25
R5836 VDDH.t260 VDDH.t259 431.25
R5837 VDDH.t241 VDDH.t260 431.25
R5838 VDDH.t258 VDDH.t241 431.25
R5839 VDDH.t486 VDDH.t488 431.25
R5840 VDDH.t484 VDDH.t486 431.25
R5841 VDDH.t489 VDDH.t484 431.25
R5842 VDDH.t487 VDDH.t485 431.25
R5843 VDDH.t485 VDDH.t482 431.25
R5844 VDDH.t482 VDDH.t481 431.25
R5845 VDDH.t322 VDDH.t531 431.25
R5846 VDDH.t424 VDDH.t322 431.25
R5847 VDDH.t534 VDDH.t424 431.25
R5848 VDDH.t324 VDDH.t446 431.25
R5849 VDDH.t446 VDDH.t321 431.25
R5850 VDDH.t321 VDDH.t323 431.25
R5851 VDDH.t340 VDDH.t37 431.25
R5852 VDDH.t519 VDDH.t340 431.25
R5853 VDDH.t36 VDDH.t519 431.25
R5854 VDDH.t41 VDDH.t356 431.25
R5855 VDDH.t356 VDDH.t520 431.25
R5856 VDDH.t520 VDDH.t40 431.25
R5857 VDDH.t460 VDDH.t63 431.25
R5858 VDDH.t461 VDDH.t460 431.25
R5859 VDDH.t60 VDDH.t461 431.25
R5860 VDDH.t465 VDDH.t579 431.25
R5861 VDDH.t579 VDDH.t59 431.25
R5862 VDDH.t59 VDDH.t61 431.25
R5863 VDDH.t421 VDDH.t532 431.25
R5864 VDDH.t422 VDDH.t421 431.25
R5865 VDDH.t423 VDDH.t422 431.25
R5866 VDDH.t420 VDDH.t445 431.25
R5867 VDDH.t445 VDDH.t447 431.25
R5868 VDDH.t447 VDDH.t533 431.25
R5869 VDDH.t35 VDDH.t341 431.25
R5870 VDDH.t39 VDDH.t35 431.25
R5871 VDDH.t255 VDDH.t39 431.25
R5872 VDDH.t518 VDDH.t253 431.25
R5873 VDDH.t253 VDDH.t254 431.25
R5874 VDDH.t254 VDDH.t357 431.25
R5875 VDDH.t65 VDDH.t464 431.25
R5876 VDDH.t62 VDDH.t65 431.25
R5877 VDDH.t463 VDDH.t62 431.25
R5878 VDDH.t577 VDDH.t578 431.25
R5879 VDDH.t578 VDDH.t462 431.25
R5880 VDDH.t462 VDDH.t576 431.25
R5881 VDDH.t240 VDDH.t449 431.25
R5882 VDDH.t375 VDDH.t379 431.25
R5883 VDDH.t408 VDDH.t409 431.25
R5884 VDDH.t284 VDDH.t396 431.25
R5885 VDDH.t395 VDDH.t284 431.25
R5886 VDDH.t443 VDDH.t440 431.25
R5887 VDDH.t441 VDDH.t443 431.25
R5888 VDDH.t441 VDDH.t444 431.25
R5889 VDDH.t442 VDDH.t444 431.25
R5890 VDDH.t525 VDDH.t494 431.25
R5891 VDDH.t495 VDDH.t525 431.25
R5892 VDDH.t495 VDDH.t493 431.25
R5893 VDDH.t493 VDDH.t496 431.25
R5894 VDDH.t501 VDDH.t73 431.25
R5895 VDDH.t74 VDDH.t501 431.25
R5896 VDDH.t70 VDDH.t74 431.25
R5897 VDDH.t500 VDDH.t70 431.25
R5898 VDDH.t500 VDDH.t72 431.25
R5899 VDDH.t72 VDDH.t498 431.25
R5900 VDDH.t498 VDDH.t499 431.25
R5901 VDDH.t499 VDDH.t71 431.25
R5902 VDDH.t398 VDDH.t77 431.25
R5903 VDDH.t77 VDDH.t400 431.25
R5904 VDDH.t400 VDDH.t78 431.25
R5905 VDDH.t75 VDDH.t78 431.25
R5906 VDDH.t75 VDDH.t399 431.25
R5907 VDDH.t399 VDDH.t76 431.25
R5908 VDDH.t76 VDDH.t397 431.25
R5909 VDDH.t397 VDDH.t289 431.25
R5910 VDDH.n648 VDDH.n647 428.048
R5911 VDDH.n687 VDDH.n99 422.024
R5912 VDDH.n157 VDDH.n99 409.976
R5913 VDDH.n1120 VDDH.n1119 406.589
R5914 VDDH.n685 VDDH.n110 397.93
R5915 VDDH.n600 VDDH.n586 395.07
R5916 VDDH.t483 VDDH.n1133 379.062
R5917 VDDH.t478 VDDH.n995 379.062
R5918 VDDH.t311 VDDH.n1046 379.062
R5919 VDDH.t530 VDDH.n1047 379.062
R5920 VDDH.t342 VDDH.n1030 379.062
R5921 VDDH.t414 VDDH.n1031 379.062
R5922 VDDH.t243 VDDH.n1039 379.062
R5923 VDDH.n1041 VDDH.t258 379.062
R5924 VDDH.t488 VDDH.n1000 379.062
R5925 VDDH.t481 VDDH.n1001 379.062
R5926 VDDH.t531 VDDH.n1005 379.062
R5927 VDDH.t323 VDDH.n1006 379.062
R5928 VDDH.t37 VDDH.n1065 379.062
R5929 VDDH.t40 VDDH.n1067 379.062
R5930 VDDH.t63 VDDH.n1024 379.062
R5931 VDDH.t61 VDDH.n1025 379.062
R5932 VDDH.t532 VDDH.n1011 379.062
R5933 VDDH.t533 VDDH.n1012 379.062
R5934 VDDH.t341 VDDH.n1016 379.062
R5935 VDDH.t357 VDDH.n1017 379.062
R5936 VDDH.t464 VDDH.n1084 379.062
R5937 VDDH.t576 VDDH.n1085 379.062
R5938 VDDH.t449 VDDH.n618 379.062
R5939 VDDH.t496 VDDH.n628 379.062
R5940 VDDH.t73 VDDH.n611 379.062
R5941 VDDH.t289 VDDH.n606 379.062
R5942 VDDH.t575 VDDH.t436 378.611
R5943 VDDH.t497 VDDH.t432 378.611
R5944 VDDH.t22 VDDH.t515 378.611
R5945 VDDH.t331 VDDH.t468 378.611
R5946 VDDH.t10 VDDH.t506 378.611
R5947 VDDH.t8 VDDH.t514 378.611
R5948 VDDH.t334 VDDH.t438 378.611
R5949 VDDH.t430 VDDH.t526 378.611
R5950 VDDH.n594 VDDH.n593 374.966
R5951 VDDH.n1044 VDDH.n1034 371.2
R5952 VDDH.n1075 VDDH.n1074 368.942
R5953 VDDH.n1082 VDDH.n1021 368.942
R5954 VDDH.n632 VDDH.n631 360.283
R5955 VDDH.n432 VDDH.n232 357.272
R5956 VDDH.n438 VDDH.n232 357.272
R5957 VDDH.n430 VDDH.n243 357.272
R5958 VDDH.n243 VDDH.n233 357.272
R5959 VDDH.n273 VDDH.n272 357.272
R5960 VDDH.n272 VDDH.n266 357.272
R5961 VDDH.n282 VDDH.n247 357.272
R5962 VDDH.n440 VDDH.n231 357.272
R5963 VDDH.n279 VDDH.n259 357.272
R5964 VDDH.n280 VDDH.n279 357.272
R5965 VDDH.n602 VDDH.n583 355.389
R5966 VDDH.n624 VDDH.n619 353.793
R5967 VDDH.n624 VDDH.n620 353.793
R5968 VDDH.n629 VDDH.n626 353.793
R5969 VDDH.n629 VDDH.n623 353.793
R5970 VDDH.n654 VDDH.n610 353.793
R5971 VDDH.n610 VDDH.n609 353.793
R5972 VDDH.n1056 VDDH.n1055 352.377
R5973 VDDH.n1083 VDDH.n1082 343.341
R5974 VDDH.n1093 VDDH.n1021 343.341
R5975 VDDH.n1096 VDDH.n1018 343.341
R5976 VDDH.n1098 VDDH.n1008 343.341
R5977 VDDH.n1114 VDDH.n1113 343.341
R5978 VDDH.n1010 VDDH.n999 343.341
R5979 VDDH.n1095 VDDH.n1094 339.954
R5980 VDDH.n1087 VDDH.n1015 339.954
R5981 VDDH.n686 VDDH.n685 339.954
R5982 VDDH.n625 VDDH.t395 332.812
R5983 VDDH.t440 VDDH.n625 332.812
R5984 VDDH.n630 VDDH.t442 332.812
R5985 VDDH.t494 VDDH.n630 332.812
R5986 VDDH.t71 VDDH.n615 332.812
R5987 VDDH.n615 VDDH.t398 332.812
R5988 VDDH.n1076 VDDH.n1026 332.8
R5989 VDDH.n1073 VDDH.n1028 332.8
R5990 VDDH.n1063 VDDH.n1062 332.8
R5991 VDDH.n1120 VDDH.n1003 332.8
R5992 VDDH.n69 VDDH.t369 330.12
R5993 VDDH.n71 VDDH.t390 330.12
R5994 VDDH.n74 VDDH.t411 330.12
R5995 VDDH.n56 VDDH.t394 330.12
R5996 VDDH.n699 VDDH.t393 330.12
R5997 VDDH.n700 VDDH.t412 330.12
R5998 VDDH.n710 VDDH.t367 330.12
R5999 VDDH.n709 VDDH.t410 330.12
R6000 VDDH.n708 VDDH.t413 330.12
R6001 VDDH.n707 VDDH.t391 330.12
R6002 VDDH.n705 VDDH.t366 330.12
R6003 VDDH.n704 VDDH.t370 330.12
R6004 VDDH.n281 VDDH.n280 325.272
R6005 VDDH.n280 VDDH.n257 325.272
R6006 VDDH.n266 VDDH.n257 325.272
R6007 VDDH.n267 VDDH.n266 325.272
R6008 VDDH.n267 VDDH.n233 325.272
R6009 VDDH.n437 VDDH.n233 325.272
R6010 VDDH.n438 VDDH.n437 325.272
R6011 VDDH.n439 VDDH.n438 325.272
R6012 VDDH.n730 VDDH.n66 321.882
R6013 VDDH.n720 VDDH.n60 321.882
R6014 VDDH.n84 VDDH.n64 321.882
R6015 VDDH.n62 VDDH.n58 321.882
R6016 VDDH.n957 VDDH.n956 321.882
R6017 VDDH.n948 VDDH.n947 321.882
R6018 VDDH.n17 VDDH.n16 321.882
R6019 VDDH.n927 VDDH.n28 321.882
R6020 VDDH.n931 VDDH.n28 321.882
R6021 VDDH.n932 VDDH.n931 321.882
R6022 VDDH.n932 VDDH.n26 321.882
R6023 VDDH.n936 VDDH.n26 321.882
R6024 VDDH.n902 VDDH.n36 321.882
R6025 VDDH.n906 VDDH.n36 321.882
R6026 VDDH.n907 VDDH.n906 321.882
R6027 VDDH.n907 VDDH.n34 321.882
R6028 VDDH.n911 VDDH.n34 321.882
R6029 VDDH.n869 VDDH.n48 321.882
R6030 VDDH.n48 VDDH.n45 321.882
R6031 VDDH.n890 VDDH.n45 321.882
R6032 VDDH.n890 VDDH.n46 321.882
R6033 VDDH.n881 VDDH.n46 321.882
R6034 VDDH.n851 VDDH.n54 321.882
R6035 VDDH.n851 VDDH.n53 321.882
R6036 VDDH.n856 VDDH.n53 321.882
R6037 VDDH.n856 VDDH.n50 321.882
R6038 VDDH.n865 VDDH.n50 321.882
R6039 VDDH.n739 VDDH.n738 321.882
R6040 VDDH.n740 VDDH.n739 321.882
R6041 VDDH.n826 VDDH.n740 321.882
R6042 VDDH.n826 VDDH.n825 321.882
R6043 VDDH.n825 VDDH.n813 321.882
R6044 VDDH.n794 VDDH.n750 321.882
R6045 VDDH.n794 VDDH.n749 321.882
R6046 VDDH.n799 VDDH.n749 321.882
R6047 VDDH.n799 VDDH.n746 321.882
R6048 VDDH.n808 VDDH.n746 321.882
R6049 VDDH.n768 VDDH.n757 321.882
R6050 VDDH.n772 VDDH.n757 321.882
R6051 VDDH.n773 VDDH.n772 321.882
R6052 VDDH.n773 VDDH.n755 321.882
R6053 VDDH.n778 VDDH.n755 321.882
R6054 VDDH.n981 VDDH.n4 321.882
R6055 VDDH.n1010 VDDH.n997 320
R6056 VDDH.n246 VDDH.n226 316.51
R6057 VDDH.n249 VDDH.n226 316.51
R6058 VDDH.n1086 VDDH.n1083 313.224
R6059 VDDH.n399 VDDH.n247 312.281
R6060 VDDH.n397 VDDH.n248 312.281
R6061 VDDH.n552 VDDH.n551 312.094
R6062 VDDH.n1018 VDDH.n1008 310.966
R6063 VDDH.n537 VDDH.n215 307.2
R6064 VDDH.n537 VDDH.n536 307.2
R6065 VDDH.n1098 VDDH.n1097 306.825
R6066 VDDH.n504 VDDH.n503 301.748
R6067 VDDH.n497 VDDH.n493 301.748
R6068 VDDH.n1097 VDDH.n1009 297.788
R6069 VDDH.n1105 VDDH.n1104 297.788
R6070 VDDH.n1131 VDDH.n1130 295.154
R6071 VDDH.n693 VDDH.n97 294.767
R6072 VDDH.n142 VDDH.n120 292.601
R6073 VDDH.n694 VDDH.n96 288.753
R6074 VDDH.n641 VDDH.n640 288
R6075 VDDH.n640 VDDH.n622 288
R6076 VDDH.n632 VDDH.n622 288
R6077 VDDH.n637 VDDH.n617 288
R6078 VDDH.n637 VDDH.n636 288
R6079 VDDH.n636 VDDH.n635 288
R6080 VDDH.n1123 VDDH.n1121 284.613
R6081 VDDH.n1114 VDDH.n999 284.613
R6082 VDDH.n1113 VDDH.n1009 283.106
R6083 VDDH.n486 VDDH.n485 281.976
R6084 VDDH.n485 VDDH.n471 281.976
R6085 VDDH.n514 VDDH.n513 281.976
R6086 VDDH.n513 VDDH.n461 281.976
R6087 VDDH.n1051 VDDH.t247 281.25
R6088 VDDH.n1074 VDDH.n1073 277.836
R6089 VDDH.n1094 VDDH.n1093 277.836
R6090 VDDH.n505 VDDH.n472 275.2
R6091 VDDH.n595 VDDH.n594 275.2
R6092 VDDH.n1064 VDDH.n1063 273.695
R6093 VDDH.n1131 VDDH.n997 272.565
R6094 VDDH.n1107 VDDH.n996 272.565
R6095 VDDH.n727 VDDH.n65 271.068
R6096 VDDH.n719 VDDH.n61 271.068
R6097 VDDH.n83 VDDH.n63 271.068
R6098 VDDH.n733 VDDH.n732 271.068
R6099 VDDH.n963 VDDH.n962 271.068
R6100 VDDH.n950 VDDH.n949 271.068
R6101 VDDH.n19 VDDH.n18 271.068
R6102 VDDH.n988 VDDH.n3 271.068
R6103 VDDH.n650 VDDH.n648 270.307
R6104 VDDH.n658 VDDH.n607 270.307
R6105 VDDH.n617 VDDH.n608 270.307
R6106 VDDH.n1096 VDDH.n1095 269.93
R6107 VDDH.n702 VDDH.t560 252.982
R6108 VDDH.n724 VDDH.t492 252.982
R6109 VDDH.n88 VDDH.t381 252.982
R6110 VDDH.n80 VDDH.t452 252.982
R6111 VDDH.n765 VDDH.t475 252.982
R6112 VDDH.n783 VDDH.t1 252.982
R6113 VDDH.n790 VDDH.t524 252.982
R6114 VDDH.n804 VDDH.t372 252.982
R6115 VDDH.n831 VDDH.t407 252.982
R6116 VDDH.n818 VDDH.t353 252.982
R6117 VDDH.n847 VDDH.t355 252.982
R6118 VDDH.n861 VDDH.t349 252.982
R6119 VDDH.n874 VDDH.t310 252.982
R6120 VDDH.n885 VDDH.t329 252.982
R6121 VDDH.n897 VDDH.t68 252.982
R6122 VDDH.n916 VDDH.t536 252.982
R6123 VDDH.n922 VDDH.t529 252.982
R6124 VDDH.n941 VDDH.t80 252.982
R6125 VDDH.n970 VDDH.t574 252.982
R6126 VDDH.n954 VDDH.t517 252.982
R6127 VDDH.n959 VDDH.t505 252.982
R6128 VDDH.n983 VDDH.t333 252.982
R6129 VDDH.n166 VDDH.n142 248.9
R6130 VDDH.n1076 VDDH.n1075 240.941
R6131 VDDH.n1045 VDDH.n1044 236.8
R6132 VDDH.n1056 VDDH.n1054 236.8
R6133 VDDH.n345 VDDH 236.048
R6134 VDDH.n644 VDDH.t409 235.939
R6135 VDDH.n631 VDDH.n607 232.66
R6136 VDDH.n100 VDDH.t17 227.737
R6137 VDDH.n148 VDDH.t392 226.81
R6138 VDDH.n1130 VDDH 225.882
R6139 VDDH.n529 VDDH.n528 224.754
R6140 VDDH.n578 VDDH.n177 224.754
R6141 VDDH.n344 VDDH.n177 224.754
R6142 VDDH.n528 VDDH.n197 224.754
R6143 VDDH.n588 VDDH.t69 216.383
R6144 VDDH.n1135 VDDH.t479 215.625
R6145 VDDH.n1135 VDDH.t477 215.625
R6146 VDDH.n1059 VDDH.t343 215.625
R6147 VDDH.n1059 VDDH.t415 215.625
R6148 VDDH.n1040 VDDH.t242 215.625
R6149 VDDH.t259 VDDH.n1040 215.625
R6150 VDDH.n1126 VDDH.t489 215.625
R6151 VDDH.n1126 VDDH.t487 215.625
R6152 VDDH.n1117 VDDH.t534 215.625
R6153 VDDH.n1117 VDDH.t324 215.625
R6154 VDDH.n1070 VDDH.t36 215.625
R6155 VDDH.n1070 VDDH.t41 215.625
R6156 VDDH.n1079 VDDH.t60 215.625
R6157 VDDH.n1079 VDDH.t465 215.625
R6158 VDDH.n1110 VDDH.t423 215.625
R6159 VDDH.n1110 VDDH.t420 215.625
R6160 VDDH.n1101 VDDH.t255 215.625
R6161 VDDH.n1101 VDDH.t518 215.625
R6162 VDDH.n1090 VDDH.t463 215.625
R6163 VDDH.n1090 VDDH.t577 215.625
R6164 VDDH.n591 VDDH.t419 209.843
R6165 VDDH.n648 VDDH.n616 207.812
R6166 VDDH.n391 VDDH.n289 206.352
R6167 VDDH.n391 VDDH.n390 206.352
R6168 VDDH.n393 VDDH.n248 205.361
R6169 VDDH.n553 VDDH.n552 205.177
R6170 VDDH.n1077 VDDH.n1076 202.918
R6171 VDDH.n1092 VDDH.n1083 202.918
R6172 VDDH.n602 VDDH.n601 201.412
R6173 VDDH.n291 VDDH.n290 200.282
R6174 VDDH.n291 VDDH.n213 200.282
R6175 VDDH.n670 VDDH.n110 200.282
R6176 VDDH.n162 VDDH.n119 200.282
R6177 VDDH.n2 VDDH.n1 200.111
R6178 VDDH.n7 VDDH.n6 200.111
R6179 VDDH.n952 VDDH.n945 200.111
R6180 VDDH.n972 VDDH.n12 200.111
R6181 VDDH.n920 VDDH.n919 200.111
R6182 VDDH.n895 VDDH.n40 200.111
R6183 VDDH.n43 VDDH.n42 200.111
R6184 VDDH.n845 VDDH.n844 200.111
R6185 VDDH.n830 VDDH.n743 200.111
R6186 VDDH.n788 VDDH.n787 200.111
R6187 VDDH.n763 VDDH.n761 200.111
R6188 VDDH.t562 VDDH.n598 199.565
R6189 VDDH.n598 VDDH.t246 199.565
R6190 VDDH.n645 VDDH.t405 193.75
R6191 VDDH.n768 VDDH.n767 191.167
R6192 VDDH.n974 VDDH.t436 189.305
R6193 VDDH.t432 VDDH.n974 189.305
R6194 VDDH.n975 VDDH.t22 189.305
R6195 VDDH.t468 VDDH.n975 189.305
R6196 VDDH.n976 VDDH.t10 189.305
R6197 VDDH.n976 VDDH.t8 189.305
R6198 VDDH.n979 VDDH.t438 189.305
R6199 VDDH.n979 VDDH.t430 189.305
R6200 VDDH.n964 VDDH.n957 185
R6201 VDDH.n965 VDDH.n956 185
R6202 VDDH.n956 VDDH.n8 185
R6203 VDDH.n951 VDDH.n948 185
R6204 VDDH.n947 VDDH.n946 185
R6205 VDDH.n947 VDDH.n9 185
R6206 VDDH.n17 VDDH.n14 185
R6207 VDDH.n16 VDDH.n15 185
R6208 VDDH.n16 VDDH.n10 185
R6209 VDDH.n779 VDDH.n778 185
R6210 VDDH.n778 VDDH.n777 185
R6211 VDDH.n780 VDDH.n755 185
R6212 VDDH.n775 VDDH.n755 185
R6213 VDDH.n773 VDDH.n754 185
R6214 VDDH.n774 VDDH.n773 185
R6215 VDDH.n772 VDDH.n758 185
R6216 VDDH.n772 VDDH.n771 185
R6217 VDDH.n759 VDDH.n757 185
R6218 VDDH.n770 VDDH.n757 185
R6219 VDDH.n769 VDDH.n768 185
R6220 VDDH.n808 VDDH.n807 185
R6221 VDDH.n809 VDDH.n808 185
R6222 VDDH.n747 VDDH.n746 185
R6223 VDDH.n746 VDDH.n745 185
R6224 VDDH.n800 VDDH.n799 185
R6225 VDDH.n799 VDDH.n798 185
R6226 VDDH.n749 VDDH.n748 185
R6227 VDDH.n796 VDDH.n749 185
R6228 VDDH.n794 VDDH.n793 185
R6229 VDDH.n795 VDDH.n794 185
R6230 VDDH.n751 VDDH.n750 185
R6231 VDDH.n776 VDDH.n750 185
R6232 VDDH.n814 VDDH.n813 185
R6233 VDDH.n823 VDDH.n813 185
R6234 VDDH.n825 VDDH.n821 185
R6235 VDDH.n825 VDDH.n824 185
R6236 VDDH.n826 VDDH.n741 185
R6237 VDDH.n827 VDDH.n826 185
R6238 VDDH.n834 VDDH.n740 185
R6239 VDDH.n812 VDDH.n740 185
R6240 VDDH.n835 VDDH.n739 185
R6241 VDDH.n811 VDDH.n739 185
R6242 VDDH.n836 VDDH.n738 185
R6243 VDDH.n810 VDDH.n738 185
R6244 VDDH.n865 VDDH.n864 185
R6245 VDDH.n866 VDDH.n865 185
R6246 VDDH.n51 VDDH.n50 185
R6247 VDDH.n50 VDDH.n49 185
R6248 VDDH.n857 VDDH.n856 185
R6249 VDDH.n856 VDDH.n855 185
R6250 VDDH.n53 VDDH.n52 185
R6251 VDDH.n853 VDDH.n53 185
R6252 VDDH.n851 VDDH.n850 185
R6253 VDDH.n852 VDDH.n851 185
R6254 VDDH.n55 VDDH.n54 185
R6255 VDDH.n822 VDDH.n54 185
R6256 VDDH.n882 VDDH.n881 185
R6257 VDDH.n881 VDDH.n880 185
R6258 VDDH.n878 VDDH.n46 185
R6259 VDDH.n879 VDDH.n46 185
R6260 VDDH.n890 VDDH.n889 185
R6261 VDDH.n891 VDDH.n890 185
R6262 VDDH.n877 VDDH.n45 185
R6263 VDDH.n45 VDDH.n44 185
R6264 VDDH.n48 VDDH.n47 185
R6265 VDDH.n867 VDDH.n48 185
R6266 VDDH.n870 VDDH.n869 185
R6267 VDDH.n869 VDDH.n868 185
R6268 VDDH.n912 VDDH.n911 185
R6269 VDDH.n911 VDDH.n910 185
R6270 VDDH.n913 VDDH.n34 185
R6271 VDDH.n909 VDDH.n34 185
R6272 VDDH.n907 VDDH.n33 185
R6273 VDDH.n908 VDDH.n907 185
R6274 VDDH.n906 VDDH.n37 185
R6275 VDDH.n906 VDDH.n905 185
R6276 VDDH.n38 VDDH.n36 185
R6277 VDDH.n904 VDDH.n36 185
R6278 VDDH.n902 VDDH.n901 185
R6279 VDDH.n903 VDDH.n902 185
R6280 VDDH.n937 VDDH.n936 185
R6281 VDDH.n936 VDDH.n935 185
R6282 VDDH.n938 VDDH.n26 185
R6283 VDDH.n934 VDDH.n26 185
R6284 VDDH.n932 VDDH.n25 185
R6285 VDDH.n933 VDDH.n932 185
R6286 VDDH.n931 VDDH.n29 185
R6287 VDDH.n931 VDDH.n930 185
R6288 VDDH.n30 VDDH.n28 185
R6289 VDDH.n929 VDDH.n28 185
R6290 VDDH.n927 VDDH.n926 185
R6291 VDDH.n928 VDDH.n927 185
R6292 VDDH.n986 VDDH.n981 185
R6293 VDDH.n981 VDDH.n980 185
R6294 VDDH.n987 VDDH.n4 185
R6295 VDDH.n58 VDDH.n57 185
R6296 VDDH.n76 VDDH.n62 185
R6297 VDDH.n731 VDDH.n62 185
R6298 VDDH.n85 VDDH.n84 185
R6299 VDDH.n75 VDDH.n64 185
R6300 VDDH.n731 VDDH.n64 185
R6301 VDDH.n721 VDDH.n720 185
R6302 VDDH.n72 VDDH.n60 185
R6303 VDDH.n731 VDDH.n60 185
R6304 VDDH.n728 VDDH.n66 185
R6305 VDDH.n730 VDDH.n729 185
R6306 VDDH.n731 VDDH.n730 185
R6307 VDDH.t16 VDDH.t338 179.685
R6308 VDDH.t338 VDDH.n144 175.309
R6309 VDDH.n496 VDDH.t545 174.853
R6310 VDDH.n474 VDDH.t547 174.853
R6311 VDDH.n1099 VDDH.n1096 173.929
R6312 VDDH.t425 VDDH.t417 168.685
R6313 VDDH.t418 VDDH.t368 168.685
R6314 VDDH.n1073 VDDH.n1072 166.024
R6315 VDDH.n1093 VDDH.n1092 166.024
R6316 VDDH.n1057 VDDH.n1056 163.766
R6317 VDDH.n1113 VDDH.n1112 160.754
R6318 VDDH.t368 VDDH.n59 158.225
R6319 VDDH.n493 VDDH.n473 155.107
R6320 VDDH.n504 VDDH.n473 155.107
R6321 VDDH.n599 VDDH.t502 154.424
R6322 VDDH.t563 VDDH.n599 154.424
R6323 VDDH.n590 VDDH.n585 152.471
R6324 VDDH.n694 VDDH.n693 152.471
R6325 VDDH.n593 VDDH.n590 152.095
R6326 VDDH.n1051 VDDH.t249 150
R6327 VDDH.n1130 VDDH.n994 148.707
R6328 VDDH.n731 VDDH.t380 144.494
R6329 VDDH.n360 VDDH.t199 139.454
R6330 VDDH.n350 VDDH.t169 139.454
R6331 VDDH.n351 VDDH.t217 139.454
R6332 VDDH.n365 VDDH.t196 139.454
R6333 VDDH.n343 VDDH.t150 139.454
R6334 VDDH.n365 VDDH.t172 139.454
R6335 VDDH.n343 VDDH.t110 139.454
R6336 VDDH.n557 VDDH.t126 139.454
R6337 VDDH.n211 VDDH.t92 139.454
R6338 VDDH.n557 VDDH.t88 139.454
R6339 VDDH.n211 VDDH.t205 139.454
R6340 VDDH.n316 VDDH.t153 139.454
R6341 VDDH.n315 VDDH.t187 139.454
R6342 VDDH.n562 VDDH.t133 139.454
R6343 VDDH.n209 VDDH.t95 139.454
R6344 VDDH.n320 VDDH.t193 139.454
R6345 VDDH.n338 VDDH.t156 139.454
R6346 VDDH.n302 VDDH.t98 139.454
R6347 VDDH.n304 VDDH.t202 139.454
R6348 VDDH.n303 VDDH.t102 139.454
R6349 VDDH.n448 VDDH.t178 139.454
R6350 VDDH.n451 VDDH.t106 139.454
R6351 VDDH.n402 VDDH.t144 139.454
R6352 VDDH.n401 VDDH.t190 139.454
R6353 VDDH.n407 VDDH.t84 139.454
R6354 VDDH.n406 VDDH.t123 139.454
R6355 VDDH.n222 VDDH.t181 139.454
R6356 VDDH.n221 VDDH.t220 139.454
R6357 VDDH.n218 VDDH.t175 139.454
R6358 VDDH.n217 VDDH.t214 139.454
R6359 VDDH.n545 VDDH.t120 139.454
R6360 VDDH.n544 VDDH.t159 139.454
R6361 VDDH.n541 VDDH.t117 139.454
R6362 VDDH.n540 VDDH.t147 139.454
R6363 VDDH.n313 VDDH.t232 139.454
R6364 VDDH.n523 VDDH.t226 139.454
R6365 VDDH.n524 VDDH.t223 139.454
R6366 VDDH.n522 VDDH.t140 139.454
R6367 VDDH.n521 VDDH.t136 139.454
R6368 VDDH.n563 VDDH.t162 139.454
R6369 VDDH.n105 VDDH.t235 139.454
R6370 VDDH.n107 VDDH.t211 139.454
R6371 VDDH.n664 VDDH.t166 139.454
R6372 VDDH.n680 VDDH.t208 139.454
R6373 VDDH.n114 VDDH.t113 139.454
R6374 VDDH.n134 VDDH.t229 139.454
R6375 VDDH.n136 VDDH.t129 139.454
R6376 VDDH.n129 VDDH.t184 139.454
R6377 VDDH.n1099 VDDH.n1098 137.036
R6378 VDDH.n316 VDDH.t154 135.662
R6379 VDDH.n315 VDDH.t189 135.662
R6380 VDDH.n304 VDDH.t203 135.662
R6381 VDDH.n303 VDDH.t105 135.662
R6382 VDDH.n402 VDDH.t145 135.662
R6383 VDDH.n401 VDDH.t192 135.662
R6384 VDDH.n407 VDDH.t86 135.662
R6385 VDDH.n406 VDDH.t125 135.662
R6386 VDDH.n222 VDDH.t182 135.662
R6387 VDDH.n221 VDDH.t222 135.662
R6388 VDDH.n218 VDDH.t176 135.662
R6389 VDDH.n217 VDDH.t216 135.662
R6390 VDDH.n545 VDDH.t121 135.662
R6391 VDDH.n544 VDDH.t161 135.662
R6392 VDDH.n541 VDDH.t118 135.662
R6393 VDDH.n540 VDDH.t149 135.662
R6394 VDDH.n662 VDDH.t168 135.362
R6395 VDDH.n372 VDDH.t206 135.312
R6396 VDDH.n372 VDDH.t93 135.312
R6397 VDDH.n250 VDDH.t100 135.312
R6398 VDDH.n312 VDDH.t234 135.312
R6399 VDDH.n564 VDDH.t135 135.312
R6400 VDDH.n556 VDDH.t91 135.312
R6401 VDDH.n556 VDDH.t128 135.312
R6402 VDDH.n342 VDDH.t111 135.312
R6403 VDDH.n342 VDDH.t151 135.312
R6404 VDDH.n366 VDDH.t174 135.312
R6405 VDDH.n366 VDDH.t198 135.312
R6406 VDDH.n349 VDDH.t170 135.312
R6407 VDDH.n104 VDDH.t237 135.312
R6408 VDDH.n104 VDDH.t236 135.312
R6409 VDDH.n106 VDDH.t213 135.312
R6410 VDDH.n106 VDDH.t212 135.312
R6411 VDDH.n113 VDDH.t115 135.312
R6412 VDDH.n113 VDDH.t116 135.312
R6413 VDDH.n681 VDDH.t210 135.312
R6414 VDDH.n133 VDDH.t231 135.312
R6415 VDDH.n133 VDDH.t230 135.312
R6416 VDDH.n135 VDDH.t131 135.312
R6417 VDDH.n135 VDDH.t132 135.312
R6418 VDDH.n130 VDDH.t185 135.312
R6419 VDDH.n665 VDDH.t167 135.312
R6420 VDDH.n351 VDDH.t219 135.127
R6421 VDDH.n351 VDDH.t218 135.127
R6422 VDDH.n451 VDDH.t109 135.127
R6423 VDDH.n451 VDDH.t108 135.127
R6424 VDDH.n523 VDDH.t228 135.127
R6425 VDDH.n523 VDDH.t227 135.127
R6426 VDDH.n524 VDDH.t225 135.127
R6427 VDDH.n524 VDDH.t224 135.127
R6428 VDDH.n522 VDDH.t143 135.127
R6429 VDDH.n522 VDDH.t142 135.127
R6430 VDDH.n521 VDDH.t139 135.127
R6431 VDDH.n521 VDDH.t138 135.127
R6432 VDDH.n563 VDDH.t165 135.127
R6433 VDDH.n563 VDDH.t164 135.127
R6434 VDDH.n449 VDDH.t180 135.026
R6435 VDDH.n174 VDDH.t179 135.026
R6436 VDDH.n352 VDDH.t508 134.712
R6437 VDDH.n352 VDDH.t201 134.712
R6438 VDDH.n362 VDDH.t200 134.712
R6439 VDDH.n362 VDDH.t171 134.712
R6440 VDDH.n363 VDDH.t197 134.712
R6441 VDDH.n363 VDDH.t152 134.712
R6442 VDDH.n210 VDDH.t90 134.712
R6443 VDDH.n210 VDDH.t207 134.712
R6444 VDDH.n314 VDDH.t233 134.712
R6445 VDDH.n314 VDDH.t195 134.712
R6446 VDDH.n317 VDDH.t188 134.712
R6447 VDDH.n317 VDDH.t155 134.712
R6448 VDDH.n560 VDDH.t134 134.712
R6449 VDDH.n560 VDDH.t97 134.712
R6450 VDDH.n559 VDDH.t127 134.712
R6451 VDDH.n559 VDDH.t94 134.712
R6452 VDDH.n321 VDDH.t194 134.712
R6453 VDDH.n321 VDDH.t555 134.712
R6454 VDDH.n323 VDDH.t51 134.712
R6455 VDDH.n323 VDDH.t278 134.712
R6456 VDDH.n325 VDDH.t306 134.712
R6457 VDDH.n325 VDDH.t53 134.712
R6458 VDDH.n327 VDDH.t264 134.712
R6459 VDDH.n327 VDDH.t303 134.712
R6460 VDDH.n329 VDDH.t551 134.712
R6461 VDDH.n329 VDDH.t294 134.712
R6462 VDDH.n307 VDDH.t280 134.712
R6463 VDDH.n307 VDDH.t158 134.712
R6464 VDDH.n341 VDDH.t173 134.712
R6465 VDDH.n341 VDDH.t112 134.712
R6466 VDDH.n340 VDDH.t157 134.712
R6467 VDDH.n340 VDDH.t101 134.712
R6468 VDDH.n305 VDDH.t104 134.712
R6469 VDDH.n305 VDDH.t204 134.712
R6470 VDDH.n308 VDDH.t292 134.712
R6471 VDDH.n308 VDDH.t265 134.712
R6472 VDDH.n309 VDDH.t313 134.712
R6473 VDDH.n309 VDDH.t276 134.712
R6474 VDDH.n310 VDDH.t281 134.712
R6475 VDDH.n310 VDDH.t317 134.712
R6476 VDDH.n311 VDDH.t556 134.712
R6477 VDDH.n311 VDDH.t261 134.712
R6478 VDDH.n331 VDDH.t304 134.712
R6479 VDDH.n331 VDDH.t557 134.712
R6480 VDDH.n403 VDDH.t191 134.712
R6481 VDDH.n403 VDDH.t146 134.712
R6482 VDDH.n408 VDDH.t124 134.712
R6483 VDDH.n408 VDDH.t87 134.712
R6484 VDDH.n219 VDDH.t215 134.712
R6485 VDDH.n219 VDDH.t177 134.712
R6486 VDDH.n223 VDDH.t221 134.712
R6487 VDDH.n223 VDDH.t183 134.712
R6488 VDDH.n542 VDDH.t148 134.712
R6489 VDDH.n542 VDDH.t119 134.712
R6490 VDDH.n546 VDDH.t160 134.712
R6491 VDDH.n546 VDDH.t122 134.712
R6492 VDDH.n191 VDDH.t296 134.712
R6493 VDDH.n191 VDDH.t569 134.712
R6494 VDDH.n202 VDDH.t282 134.712
R6495 VDDH.n202 VDDH.t507 134.712
R6496 VDDH.n203 VDDH.t239 134.712
R6497 VDDH.n203 VDDH.t283 134.712
R6498 VDDH.n204 VDDH.t43 134.712
R6499 VDDH.n204 VDDH.t295 134.712
R6500 VDDH.n194 VDDH.t267 134.712
R6501 VDDH.n194 VDDH.t362 134.712
R6502 VDDH.n192 VDDH.t565 134.712
R6503 VDDH.n192 VDDH.t385 134.712
R6504 VDDH.n355 VDDH.t513 134.712
R6505 VDDH.n355 VDDH.t384 134.712
R6506 VDDH.n354 VDDH.t383 134.712
R6507 VDDH.n354 VDDH.t571 134.712
R6508 VDDH.n353 VDDH.t358 134.712
R6509 VDDH.n353 VDDH.t47 134.712
R6510 VDDH.n201 VDDH.t96 134.712
R6511 VDDH.n201 VDDH.t269 134.712
R6512 VDDH.n373 VDDH.t568 134.712
R6513 VDDH.n373 VDDH.t359 134.712
R6514 VDDH.n374 VDDH.t364 134.712
R6515 VDDH.n374 VDDH.t386 134.712
R6516 VDDH.n376 VDDH.t316 134.712
R6517 VDDH.n376 VDDH.t512 134.712
R6518 VDDH.n377 VDDH.t299 134.712
R6519 VDDH.n377 VDDH.t567 134.712
R6520 VDDH.n379 VDDH.t361 134.712
R6521 VDDH.n379 VDDH.t290 134.712
R6522 VDDH.n380 VDDH.t387 134.712
R6523 VDDH.n380 VDDH.t314 134.712
R6524 VDDH.n382 VDDH.t509 134.712
R6525 VDDH.n382 VDDH.t270 134.712
R6526 VDDH.n383 VDDH.t564 134.712
R6527 VDDH.n383 VDDH.t360 134.712
R6528 VDDH.n385 VDDH.t553 134.712
R6529 VDDH.n385 VDDH.t511 134.712
R6530 VDDH.n386 VDDH.t55 134.712
R6531 VDDH.n386 VDDH.t566 134.712
R6532 VDDH.n292 VDDH.t274 134.712
R6533 VDDH.n292 VDDH.t302 134.712
R6534 VDDH.n293 VDDH.t554 134.712
R6535 VDDH.n293 VDDH.t552 134.712
R6536 VDDH.n294 VDDH.t49 134.712
R6537 VDDH.n294 VDDH.t263 134.712
R6538 VDDH.n295 VDDH.t510 134.712
R6539 VDDH.n295 VDDH.t305 134.712
R6540 VDDH.n296 VDDH.t45 134.712
R6541 VDDH.n296 VDDH.t388 134.712
R6542 VDDH.n297 VDDH.t572 134.712
R6543 VDDH.n297 VDDH.t298 134.712
R6544 VDDH.n298 VDDH.t315 134.712
R6545 VDDH.n298 VDDH.t363 134.712
R6546 VDDH.n299 VDDH.t570 134.712
R6547 VDDH.n299 VDDH.t389 134.712
R6548 VDDH.n300 VDDH.t293 134.712
R6549 VDDH.n300 VDDH.t318 134.712
R6550 VDDH.n301 VDDH.t319 134.712
R6551 VDDH.n301 VDDH.t300 134.712
R6552 VDDH.n115 VDDH.t209 134.712
R6553 VDDH.n115 VDDH.t580 134.712
R6554 VDDH.n116 VDDH.t582 134.712
R6555 VDDH.n116 VDDH.t57 134.712
R6556 VDDH.n117 VDDH.t347 134.712
R6557 VDDH.n117 VDDH.t583 134.712
R6558 VDDH.n127 VDDH.t346 134.712
R6559 VDDH.n127 VDDH.t186 134.712
R6560 VDDH.n124 VDDH.t271 134.712
R6561 VDDH.n124 VDDH.t581 134.712
R6562 VDDH.n126 VDDH.t584 134.712
R6563 VDDH.n126 VDDH.t272 134.712
R6564 VDDH.n147 VDDH.n146 129.44
R6565 VDDH.n635 VDDH.n607 127.624
R6566 VDDH.t538 VDDH.n144 125.675
R6567 VDDH.n1112 VDDH.n1010 123.859
R6568 VDDH.t33 VDDH.n415 117.921
R6569 VDDH.t31 VDDH.n413 117.921
R6570 VDDH VDDH.n1129 117.46
R6571 VDDH.t130 VDDH.t30 113.218
R6572 VDDH.t251 VDDH.t56 113.218
R6573 VDDH.t29 VDDH.t28 113.218
R6574 VDDH.t28 VDDH.t114 113.218
R6575 VDDH.n576 VDDH.t137 109.784
R6576 VDDH.n692 VDDH.n99 106.541
R6577 VDDH.n693 VDDH.n692 106.165
R6578 VDDH.t30 VDDH.n161 105.088
R6579 VDDH.n575 VDDH.n181 105.073
R6580 VDDH.n713 VDDH.t365 102.35
R6581 VDDH.n158 VDDH.n97 101.272
R6582 VDDH.t66 VDDH.t382 100.906
R6583 VDDH.t256 VDDH.t365 100.906
R6584 VDDH.n597 VDDH.t69 100.243
R6585 VDDH.n595 VDDH.n585 100.141
R6586 VDDH.n673 VDDH.t29 99.0655
R6587 VDDH.n150 VDDH.n97 96.9471
R6588 VDDH.t252 VDDH.t538 95.9301
R6589 VDDH.t392 VDDH.t257 95.9301
R6590 VDDH.n777 VDDH.n775 92.2149
R6591 VDDH.n809 VDDH.n745 92.2149
R6592 VDDH.n824 VDDH.n823 92.2149
R6593 VDDH.n866 VDDH.n49 92.2149
R6594 VDDH.n880 VDDH.n879 92.2149
R6595 VDDH.n910 VDDH.n909 92.2149
R6596 VDDH.n935 VDDH.n934 92.2149
R6597 VDDH.t474 VDDH.n769 89.3332
R6598 VDDH.n776 VDDH.t523 89.3332
R6599 VDDH.t406 VDDH.n810 89.3332
R6600 VDDH.n822 VDDH.t354 89.3332
R6601 VDDH.n868 VDDH.t309 89.3332
R6602 VDDH.t67 VDDH.n903 89.3332
R6603 VDDH.t528 VDDH.n928 89.3332
R6604 VDDH.n962 VDDH.n957 86.068
R6605 VDDH.n949 VDDH.n948 86.068
R6606 VDDH.n18 VDDH.n17 86.068
R6607 VDDH.n4 VDDH.n3 86.068
R6608 VDDH.n732 VDDH.n58 86.068
R6609 VDDH.n84 VDDH.n63 86.068
R6610 VDDH.n720 VDDH.n61 86.068
R6611 VDDH.n66 VDDH.n65 86.068
R6612 VDDH.n482 VDDH.t550 84.6474
R6613 VDDH.n484 VDDH.t546 84.6474
R6614 VDDH.n499 VDDH.t549 84.6474
R6615 VDDH.n501 VDDH.t548 84.6474
R6616 VDDH.n769 VDDH.t58 84.5303
R6617 VDDH.t459 VDDH.n776 84.5303
R6618 VDDH.n810 VDDH.t351 84.5303
R6619 VDDH.t38 VDDH.n822 84.5303
R6620 VDDH.n868 VDDH.t451 84.5303
R6621 VDDH.n903 VDDH.t537 84.5303
R6622 VDDH.n928 VDDH.t81 84.5303
R6623 VDDH.n145 VDDH.t417 84.3432
R6624 VDDH.n145 VDDH.t418 84.3432
R6625 VDDH.n777 VDDH.t503 82.6092
R6626 VDDH.t373 VDDH.n809 82.6092
R6627 VDDH.n823 VDDH.t561 82.6092
R6628 VDDH.t339 VDDH.n866 82.6092
R6629 VDDH.n880 VDDH.t374 82.6092
R6630 VDDH.n910 VDDH.t244 82.6092
R6631 VDDH.n935 VDDH.t521 82.6092
R6632 VDDH.t466 VDDH.n160 82.5045
R6633 VDDH.n165 VDDH.t467 82.5045
R6634 VDDH.n147 VDDH.t252 81.8009
R6635 VDDH.n601 VDDH.n585 80.1887
R6636 VDDH.n649 VDDH 77.9299
R6637 VDDH.t467 VDDH.t466 77.6867
R6638 VDDH.n258 VDDH.n247 74.7248
R6639 VDDH.n274 VDDH.n259 74.7248
R6640 VDDH.n273 VDDH.n244 74.7248
R6641 VDDH.n433 VDDH.n430 74.7248
R6642 VDDH.n432 VDDH.n431 74.7248
R6643 VDDH.n431 VDDH.n231 74.7248
R6644 VDDH VDDH.n258 73.2546
R6645 VDDH.n274 VDDH 73.2546
R6646 VDDH.n433 VDDH 73.2546
R6647 VDDH.n164 VDDH.t130 72.869
R6648 VDDH.t114 VDDH.n672 72.869
R6649 VDDH.n1044 VDDH.n1043 72.6593
R6650 VDDH.n599 VDDH.t419 72.653
R6651 VDDH.n599 VDDH.t562 72.653
R6652 VDDH.n1054 VDDH.n1033 72.2828
R6653 VDDH.n1048 VDDH.n1045 72.2828
R6654 VDDH.n1055 VDDH.n1003 72.2828
R6655 VDDH.n1043 VDDH.n1042 72.2828
R6656 VDDH.n1042 VDDH.n1028 72.2828
R6657 VDDH.n1038 VDDH.n1026 72.2828
R6658 VDDH.n1032 VDDH.n1029 72.2828
R6659 VDDH.n1062 VDDH.n1029 72.2828
R6660 VDDH.n1129 VDDH.n998 72.2828
R6661 VDDH.n1121 VDDH.n1002 72.2828
R6662 VDDH.n1114 VDDH.n1002 72.2828
R6663 VDDH.n1007 VDDH.n1004 72.2828
R6664 VDDH.n1008 VDDH.n1007 72.2828
R6665 VDDH.n1066 VDDH.n1064 72.2828
R6666 VDDH.n1066 VDDH.n1018 72.2828
R6667 VDDH.n1074 VDDH.n1027 72.2828
R6668 VDDH.n1027 VDDH.n1021 72.2828
R6669 VDDH.n1075 VDDH.n1022 72.2828
R6670 VDDH.n1082 VDDH.n1022 72.2828
R6671 VDDH.n1123 VDDH.n1122 72.2828
R6672 VDDH.n1122 VDDH.n999 72.2828
R6673 VDDH.n1106 VDDH.n997 72.2828
R6674 VDDH.n1107 VDDH.n1106 72.2828
R6675 VDDH.n1013 VDDH.n1009 72.2828
R6676 VDDH.n1105 VDDH.n1013 72.2828
R6677 VDDH.n1097 VDDH.n1014 72.2828
R6678 VDDH.n1104 VDDH.n1014 72.2828
R6679 VDDH.n1095 VDDH.n1019 72.2828
R6680 VDDH.n1019 VDDH.n1015 72.2828
R6681 VDDH.n1094 VDDH.n1020 72.2828
R6682 VDDH.n1087 VDDH.n1020 72.2828
R6683 VDDH.n1132 VDDH.n1131 72.2828
R6684 VDDH.n1132 VDDH.n996 72.2828
R6685 VDDH.n636 VDDH.n627 72.2828
R6686 VDDH.n627 VDDH.n622 72.2828
R6687 VDDH.n621 VDDH.n617 72.2828
R6688 VDDH.n641 VDDH.n621 72.2828
R6689 VDDH.n650 VDDH.n649 72.2828
R6690 VDDH.n613 VDDH.n612 72.2828
R6691 VDDH.n612 VDDH.n608 72.2828
R6692 VDDH.n659 VDDH.n658 72.2828
R6693 VDDH.t545 VDDH.n467 71.3334
R6694 VDDH.t547 VDDH.n467 71.3334
R6695 VDDH.n731 VDDH.n59 66.0363
R6696 VDDH.n489 VDDH.t345 64.1959
R6697 VDDH.n672 VDDH.n111 63.1385
R6698 VDDH.n771 VDDH.t4 59.5556
R6699 VDDH.n796 VDDH.t426 59.5556
R6700 VDDH.n812 VDDH.t24 59.5556
R6701 VDDH.n853 VDDH.t12 59.5556
R6702 VDDH.t2 VDDH.n44 59.5556
R6703 VDDH.n905 VDDH.t472 59.5556
R6704 VDDH.n930 VDDH.t20 59.5556
R6705 VDDH.n119 VDDH.n96 57.977
R6706 VDDH.t434 VDDH.n774 57.6345
R6707 VDDH.n798 VDDH.t470 57.6345
R6708 VDDH.n827 VDDH.t18 57.6345
R6709 VDDH.n855 VDDH.t6 57.6345
R6710 VDDH.n891 VDDH.t428 57.6345
R6711 VDDH.t26 VDDH.n908 57.6345
R6712 VDDH.t14 VDDH.n933 57.6345
R6713 VDDH.n160 VDDH.n149 55.8602
R6714 VDDH.n167 VDDH.n96 54.2123
R6715 VDDH.n171 VDDH.n130 52.8457
R6716 VDDH.n691 VDDH.n102 50.7802
R6717 VDDH.n103 VDDH.n102 50.7802
R6718 VDDH.n145 VDDH.t66 50.4534
R6719 VDDH VDDH.n429 50.2491
R6720 VDDH.n419 VDDH.t34 49.8991
R6721 VDDH.n411 VDDH.t32 49.8991
R6722 VDDH.n962 VDDH.n8 49.4675
R6723 VDDH.n949 VDDH.n9 49.4675
R6724 VDDH.n18 VDDH.n10 49.4675
R6725 VDDH.n980 VDDH.n3 49.4675
R6726 VDDH.n732 VDDH.n731 49.4675
R6727 VDDH.n731 VDDH.n63 49.4675
R6728 VDDH.n731 VDDH.n61 49.4675
R6729 VDDH.n731 VDDH.n65 49.4675
R6730 VDDH.n508 VDDH.n467 49.2055
R6731 VDDH.n459 VDDH.t402 48.2714
R6732 VDDH.n459 VDDH.t404 48.2714
R6733 VDDH.n454 VDDH.t527 48.2714
R6734 VDDH.n454 VDDH.t403 48.2714
R6735 VDDH.n417 VDDH.t33 48.1348
R6736 VDDH.n417 VDDH.t31 48.1348
R6737 VDDH.n567 VDDH.n566 47.9922
R6738 VDDH.n774 VDDH.n756 47.0682
R6739 VDDH.n798 VDDH.n797 47.0682
R6740 VDDH.n828 VDDH.n827 47.0682
R6741 VDDH.n855 VDDH.n854 47.0682
R6742 VDDH.n892 VDDH.n891 47.0682
R6743 VDDH.n908 VDDH.n35 47.0682
R6744 VDDH.n933 VDDH.n27 47.0682
R6745 VDDH.n165 VDDH.n164 46.3713
R6746 VDDH.n1047 VDDH.n1033 46.2505
R6747 VDDH.n1048 VDDH.n1046 46.2505
R6748 VDDH.n1055 VDDH.n1031 46.2505
R6749 VDDH.n1042 VDDH.n1041 46.2505
R6750 VDDH.n1039 VDDH.n1038 46.2505
R6751 VDDH.n1030 VDDH.n1029 46.2505
R6752 VDDH.n1001 VDDH.n998 46.2505
R6753 VDDH.n1006 VDDH.n1002 46.2505
R6754 VDDH.n1007 VDDH.n1005 46.2505
R6755 VDDH.n1067 VDDH.n1066 46.2505
R6756 VDDH.n1065 VDDH.n1027 46.2505
R6757 VDDH.n1025 VDDH.n1022 46.2505
R6758 VDDH.n1024 VDDH.n1023 46.2505
R6759 VDDH.n1122 VDDH.n1000 46.2505
R6760 VDDH.n1106 VDDH.n1012 46.2505
R6761 VDDH.n1013 VDDH.n1011 46.2505
R6762 VDDH.n1017 VDDH.n1014 46.2505
R6763 VDDH.n1019 VDDH.n1016 46.2505
R6764 VDDH.n1085 VDDH.n1020 46.2505
R6765 VDDH.n1086 VDDH.n1084 46.2505
R6766 VDDH.n1133 VDDH.n1132 46.2505
R6767 VDDH.n1138 VDDH.n995 46.2505
R6768 VDDH.n624 VDDH.n621 46.2505
R6769 VDDH.n625 VDDH.n624 46.2505
R6770 VDDH.n629 VDDH.n627 46.2505
R6771 VDDH.n630 VDDH.n629 46.2505
R6772 VDDH.n631 VDDH.n628 46.2505
R6773 VDDH.n618 VDDH.n616 46.2505
R6774 VDDH.n649 VDDH.n611 46.2505
R6775 VDDH.n612 VDDH.n610 46.2505
R6776 VDDH.n615 VDDH.n610 46.2505
R6777 VDDH.n659 VDDH.n606 46.2505
R6778 VDDH.t291 VDDH.t275 45.388
R6779 VDDH.t54 VDDH.t288 45.388
R6780 VDDH.n771 VDDH.n756 45.1471
R6781 VDDH.n797 VDDH.n796 45.1471
R6782 VDDH.n828 VDDH.n812 45.1471
R6783 VDDH.n854 VDDH.n853 45.1471
R6784 VDDH.n892 VDDH.n44 45.1471
R6785 VDDH.n905 VDDH.n35 45.1471
R6786 VDDH.n930 VDDH.n27 45.1471
R6787 VDDH.t246 VDDH.n597 45.0634
R6788 VDDH.t558 VDDH.t85 44.7845
R6789 VDDH.t238 VDDH.t559 43.3359
R6790 VDDH.n505 VDDH.n504 41.6919
R6791 VDDH.n493 VDDH.n492 41.6919
R6792 VDDH.n241 VDDH.t266 41.2839
R6793 VDDH.n277 VDDH.t46 40.801
R6794 VDDH.n1063 VDDH.n1004 37.2711
R6795 VDDH.n1121 VDDH.n1120 37.2711
R6796 VDDH.n729 VDDH.n728 36.1417
R6797 VDDH.n728 VDDH.n727 36.1417
R6798 VDDH.n721 VDDH.n72 36.1417
R6799 VDDH.n721 VDDH.n719 36.1417
R6800 VDDH.n85 VDDH.n75 36.1417
R6801 VDDH.n85 VDDH.n83 36.1417
R6802 VDDH.n965 VDDH.n964 36.1417
R6803 VDDH.n964 VDDH.n963 36.1417
R6804 VDDH.n951 VDDH.n946 36.1417
R6805 VDDH.n951 VDDH.n950 36.1417
R6806 VDDH.n15 VDDH.n14 36.1417
R6807 VDDH.n19 VDDH.n14 36.1417
R6808 VDDH.n926 VDDH.n30 36.1417
R6809 VDDH.n30 VDDH.n29 36.1417
R6810 VDDH.n29 VDDH.n25 36.1417
R6811 VDDH.n938 VDDH.n25 36.1417
R6812 VDDH.n938 VDDH.n937 36.1417
R6813 VDDH.n901 VDDH.n38 36.1417
R6814 VDDH.n38 VDDH.n37 36.1417
R6815 VDDH.n37 VDDH.n33 36.1417
R6816 VDDH.n913 VDDH.n33 36.1417
R6817 VDDH.n913 VDDH.n912 36.1417
R6818 VDDH.n870 VDDH.n47 36.1417
R6819 VDDH.n877 VDDH.n47 36.1417
R6820 VDDH.n889 VDDH.n877 36.1417
R6821 VDDH.n889 VDDH.n878 36.1417
R6822 VDDH.n882 VDDH.n878 36.1417
R6823 VDDH.n850 VDDH.n55 36.1417
R6824 VDDH.n850 VDDH.n52 36.1417
R6825 VDDH.n857 VDDH.n52 36.1417
R6826 VDDH.n857 VDDH.n51 36.1417
R6827 VDDH.n864 VDDH.n51 36.1417
R6828 VDDH.n836 VDDH.n835 36.1417
R6829 VDDH.n835 VDDH.n834 36.1417
R6830 VDDH.n834 VDDH.n741 36.1417
R6831 VDDH.n821 VDDH.n741 36.1417
R6832 VDDH.n821 VDDH.n814 36.1417
R6833 VDDH.n793 VDDH.n751 36.1417
R6834 VDDH.n793 VDDH.n748 36.1417
R6835 VDDH.n800 VDDH.n748 36.1417
R6836 VDDH.n800 VDDH.n747 36.1417
R6837 VDDH.n807 VDDH.n747 36.1417
R6838 VDDH.n759 VDDH.n758 36.1417
R6839 VDDH.n758 VDDH.n754 36.1417
R6840 VDDH.n780 VDDH.n754 36.1417
R6841 VDDH.n780 VDDH.n779 36.1417
R6842 VDDH.n988 VDDH.n987 36.1417
R6843 VDDH.n987 VDDH.n986 36.1417
R6844 VDDH.n76 VDDH.n57 36.1417
R6845 VDDH.n733 VDDH.n57 36.1417
R6846 VDDH.n146 VDDH.n145 35.5918
R6847 VDDH.n604 VDDH.n603 35.2755
R6848 VDDH.t262 VDDH.t454 35.1276
R6849 VDDH.n492 VDDH.n472 35.0123
R6850 VDDH.t48 VDDH.t541 34.6447
R6851 VDDH.t4 VDDH.n770 32.6598
R6852 VDDH.t426 VDDH.n795 32.6598
R6853 VDDH.t24 VDDH.n811 32.6598
R6854 VDDH.t12 VDDH.n852 32.6598
R6855 VDDH.n867 VDDH.t2 32.6598
R6856 VDDH.t472 VDDH.n904 32.6598
R6857 VDDH.t20 VDDH.n929 32.6598
R6858 VDDH.t0 VDDH.t434 31.6992
R6859 VDDH.t470 VDDH.t371 31.6992
R6860 VDDH.t352 VDDH.t18 31.6992
R6861 VDDH.t6 VDDH.t348 31.6992
R6862 VDDH.t328 VDDH.t428 31.6992
R6863 VDDH.t535 VDDH.t26 31.6992
R6864 VDDH.t79 VDDH.t14 31.6992
R6865 VDDH.n284 VDDH.t99 31.6269
R6866 VDDH.t245 VDDH.t455 31.1441
R6867 VDDH.n238 VDDH.t52 31.1441
R6868 VDDH.n601 VDDH.n600 30.8338
R6869 VDDH.t286 VDDH.t268 30.5405
R6870 VDDH.t336 VDDH.t287 29.092
R6871 VDDH.t277 VDDH.t325 29.092
R6872 VDDH.n534 VDDH.t107 28.9077
R6873 VDDH.t544 VDDH.t279 28.6091
R6874 VDDH.n1 VDDH.t439 27.6955
R6875 VDDH.n1 VDDH.t431 27.6955
R6876 VDDH.n6 VDDH.t11 27.6955
R6877 VDDH.n6 VDDH.t9 27.6955
R6878 VDDH.n945 VDDH.t23 27.6955
R6879 VDDH.n945 VDDH.t469 27.6955
R6880 VDDH.n12 VDDH.t437 27.6955
R6881 VDDH.n12 VDDH.t433 27.6955
R6882 VDDH.n919 VDDH.t21 27.6955
R6883 VDDH.n919 VDDH.t15 27.6955
R6884 VDDH.n40 VDDH.t473 27.6955
R6885 VDDH.n40 VDDH.t27 27.6955
R6886 VDDH.n42 VDDH.t3 27.6955
R6887 VDDH.n42 VDDH.t429 27.6955
R6888 VDDH.n844 VDDH.t13 27.6955
R6889 VDDH.n844 VDDH.t7 27.6955
R6890 VDDH.n743 VDDH.t25 27.6955
R6891 VDDH.n743 VDDH.t19 27.6955
R6892 VDDH.n787 VDDH.t427 27.6955
R6893 VDDH.n787 VDDH.t471 27.6955
R6894 VDDH.n761 VDDH.t5 27.6955
R6895 VDDH.n761 VDDH.t435 27.6955
R6896 VDDH.t52 VDDH.t335 26.4363
R6897 VDDH.n602 VDDH.n584 26.4291
R6898 VDDH.n599 VDDH.n584 26.4291
R6899 VDDH.t543 VDDH.t99 25.9535
R6900 VDDH.n596 VDDH.n595 23.1255
R6901 VDDH.n597 VDDH.n596 23.1255
R6902 VDDH.n159 VDDH.n158 23.1255
R6903 VDDH.n160 VDDH.n159 23.1255
R6904 VDDH.n692 VDDH.n98 23.1255
R6905 VDDH.n165 VDDH.n98 23.1255
R6906 VDDH.n429 VDDH.n244 23.0059
R6907 VDDH.n270 VDDH.t48 22.9357
R6908 VDDH.n270 VDDH.t262 22.4529
R6909 VDDH.n511 VDDH.t345 21.5134
R6910 VDDH.n511 VDDH.t401 21.5134
R6911 VDDH.t44 VDDH.t453 20.8836
R6912 VDDH.t301 VDDH.t320 20.4008
R6913 VDDH.t89 VDDH.n443 19.5719
R6914 VDDH.t103 VDDH.t543 19.4351
R6915 VDDH.n713 VDDH.n712 19.4051
R6916 VDDH.t335 VDDH.t42 18.9522
R6917 VDDH.n494 VDDH.n473 16.8187
R6918 VDDH.n494 VDDH.n467 16.8187
R6919 VDDH.n495 VDDH.n475 16.8187
R6920 VDDH.n495 VDDH.n467 16.8187
R6921 VDDH.n416 VDDH.n412 16.8187
R6922 VDDH.n417 VDDH.n416 16.8187
R6923 VDDH.n422 VDDH.n418 16.8187
R6924 VDDH.n418 VDDH.n417 16.8187
R6925 VDDH.n594 VDDH.n588 16.8187
R6926 VDDH.t46 VDDH.t544 16.7794
R6927 VDDH.t539 VDDH.n574 16.538
R6928 VDDH.t266 VDDH.t336 16.2966
R6929 VDDH.n763 VDDH.n762 16.2626
R6930 VDDH.n788 VDDH.n744 16.2626
R6931 VDDH.n830 VDDH.n829 16.2626
R6932 VDDH.n845 VDDH.n41 16.2626
R6933 VDDH.n893 VDDH.n43 16.2626
R6934 VDDH.n895 VDDH.n894 16.2626
R6935 VDDH.n920 VDDH.n11 16.2626
R6936 VDDH.n973 VDDH.n972 16.2626
R6937 VDDH.n952 VDDH.n5 16.2626
R6938 VDDH.n977 VDDH.n7 16.2626
R6939 VDDH.n978 VDDH.n2 16.2626
R6940 VDDH.n660 VDDH.n659 15.6337
R6941 VDDH.n262 VDDH.t542 15.5723
R6942 VDDH.t326 VDDH.n262 15.5723
R6943 VDDH.n276 VDDH.t453 15.5723
R6944 VDDH.t320 VDDH.n182 15.5723
R6945 VDDH.n435 VDDH.t327 15.5723
R6946 VDDH.n435 VDDH.t337 15.5723
R6947 VDDH.t325 VDDH.n237 15.5723
R6948 VDDH.n590 VDDH.n589 15.4172
R6949 VDDH.n762 VDDH.n756 15.4172
R6950 VDDH.n797 VDDH.n744 15.4172
R6951 VDDH.n829 VDDH.n828 15.4172
R6952 VDDH.n854 VDDH.n41 15.4172
R6953 VDDH.n893 VDDH.n892 15.4172
R6954 VDDH.n894 VDDH.n35 15.4172
R6955 VDDH.n27 VDDH.n11 15.4172
R6956 VDDH.n974 VDDH.n973 15.4172
R6957 VDDH.n975 VDDH.n5 15.4172
R6958 VDDH.n977 VDDH.n976 15.4172
R6959 VDDH.n979 VDDH.n978 15.4172
R6960 VDDH.n467 VDDH.t401 14.9909
R6961 VDDH.n589 VDDH.n587 14.8961
R6962 VDDH.n146 VDDH.t256 14.8631
R6963 VDDH.t50 VDDH.t286 14.848
R6964 VDDH.n574 VDDH.t540 14.6066
R6965 VDDH.n1139 VDDH.n1138 14.4353
R6966 VDDH.n238 VDDH.t238 14.2445
R6967 VDDH.n673 VDDH.t56 14.1526
R6968 VDDH.t257 VDDH.n147 14.1297
R6969 VDDH.n426 VDDH.n425 13.8332
R6970 VDDH.n442 VDDH.t85 12.7959
R6971 VDDH.t42 VDDH.t337 12.1924
R6972 VDDH.t542 VDDH.t103 11.7095
R6973 VDDH.n443 VDDH.n442 11.5888
R6974 VDDH.n289 VDDH.n288 11.563
R6975 VDDH.n288 VDDH.n287 11.563
R6976 VDDH.n290 VDDH.n188 11.563
R6977 VDDH.n534 VDDH.n188 11.563
R6978 VDDH.n445 VDDH.n213 11.563
R6979 VDDH.n534 VDDH.n445 11.563
R6980 VDDH.n390 VDDH.n187 11.563
R6981 VDDH.n287 VDDH.n187 11.563
R6982 VDDH.n593 VDDH.n592 11.563
R6983 VDDH.n671 VDDH.n670 11.563
R6984 VDDH.n672 VDDH.n671 11.563
R6985 VDDH.n163 VDDH.n162 11.563
R6986 VDDH.n164 VDDH.n163 11.563
R6987 VDDH.n152 VDDH.n94 11.4005
R6988 VDDH.n976 VDDH.n8 11.31
R6989 VDDH.n975 VDDH.n9 11.31
R6990 VDDH.n974 VDDH.n10 11.31
R6991 VDDH.n980 VDDH.n979 11.31
R6992 VDDH.n150 VDDH.n95 11.2946
R6993 VDDH.n676 VDDH.n675 11.2946
R6994 VDDH.n592 VDDH.n587 11.1723
R6995 VDDH.n151 VDDH.n149 10.9826
R6996 VDDH.t541 VDDH.t301 10.7438
R6997 VDDH.n992 VDDH.t285 10.5739
R6998 VDDH.n446 VDDH.n197 10.2783
R6999 VDDH.n531 VDDH.n446 10.2783
R7000 VDDH.n530 VDDH.n529 10.2783
R7001 VDDH.n531 VDDH.n530 10.2783
R7002 VDDH.n578 VDDH.n577 10.2783
R7003 VDDH.n577 VDDH.n576 10.2783
R7004 VDDH.n344 VDDH.n180 10.2783
R7005 VDDH.n576 VDDH.n180 10.2783
R7006 VDDH.n591 VDDH.n583 10.2783
R7007 VDDH.t454 VDDH.t44 10.261
R7008 VDDH.n716 VDDH.n715 9.73734
R7009 VDDH.n715 VDDH.n59 9.73734
R7010 VDDH.n714 VDDH.n90 9.73734
R7011 VDDH.n714 VDDH.n713 9.66826
R7012 VDDH.n983 VDDH.n982 9.3005
R7013 VDDH.n984 VDDH.n983 9.3005
R7014 VDDH.n986 VDDH.n985 9.3005
R7015 VDDH.n987 VDDH.n2 9.3005
R7016 VDDH.n989 VDDH.n988 9.3005
R7017 VDDH.n959 VDDH.n958 9.3005
R7018 VDDH.n960 VDDH.n959 9.3005
R7019 VDDH.n963 VDDH.n961 9.3005
R7020 VDDH.n964 VDDH.n7 9.3005
R7021 VDDH.n966 VDDH.n965 9.3005
R7022 VDDH.n954 VDDH.n953 9.3005
R7023 VDDH.n955 VDDH.n954 9.3005
R7024 VDDH.n950 VDDH.n944 9.3005
R7025 VDDH.n952 VDDH.n951 9.3005
R7026 VDDH.n946 VDDH.n21 9.3005
R7027 VDDH.n971 VDDH.n970 9.3005
R7028 VDDH.n970 VDDH.n969 9.3005
R7029 VDDH.n20 VDDH.n19 9.3005
R7030 VDDH.n972 VDDH.n14 9.3005
R7031 VDDH.n15 VDDH.n13 9.3005
R7032 VDDH.n941 VDDH.n940 9.3005
R7033 VDDH.n942 VDDH.n941 9.3005
R7034 VDDH.n923 VDDH.n922 9.3005
R7035 VDDH.n922 VDDH.n921 9.3005
R7036 VDDH.n937 VDDH.n23 9.3005
R7037 VDDH.n939 VDDH.n938 9.3005
R7038 VDDH.n25 VDDH.n24 9.3005
R7039 VDDH.n918 VDDH.n29 9.3005
R7040 VDDH.n924 VDDH.n30 9.3005
R7041 VDDH.n926 VDDH.n925 9.3005
R7042 VDDH.n916 VDDH.n915 9.3005
R7043 VDDH.n917 VDDH.n916 9.3005
R7044 VDDH.n898 VDDH.n897 9.3005
R7045 VDDH.n897 VDDH.n896 9.3005
R7046 VDDH.n912 VDDH.n31 9.3005
R7047 VDDH.n914 VDDH.n913 9.3005
R7048 VDDH.n33 VDDH.n32 9.3005
R7049 VDDH.n39 VDDH.n37 9.3005
R7050 VDDH.n899 VDDH.n38 9.3005
R7051 VDDH.n901 VDDH.n900 9.3005
R7052 VDDH.n886 VDDH.n885 9.3005
R7053 VDDH.n885 VDDH.n884 9.3005
R7054 VDDH.n874 VDDH.n873 9.3005
R7055 VDDH.n875 VDDH.n874 9.3005
R7056 VDDH.n883 VDDH.n882 9.3005
R7057 VDDH.n887 VDDH.n878 9.3005
R7058 VDDH.n889 VDDH.n888 9.3005
R7059 VDDH.n877 VDDH.n876 9.3005
R7060 VDDH.n872 VDDH.n47 9.3005
R7061 VDDH.n871 VDDH.n870 9.3005
R7062 VDDH.n861 VDDH.n860 9.3005
R7063 VDDH.n862 VDDH.n861 9.3005
R7064 VDDH.n848 VDDH.n847 9.3005
R7065 VDDH.n847 VDDH.n846 9.3005
R7066 VDDH.n864 VDDH.n863 9.3005
R7067 VDDH.n859 VDDH.n51 9.3005
R7068 VDDH.n858 VDDH.n857 9.3005
R7069 VDDH.n843 VDDH.n52 9.3005
R7070 VDDH.n850 VDDH.n849 9.3005
R7071 VDDH.n842 VDDH.n55 9.3005
R7072 VDDH.n819 VDDH.n818 9.3005
R7073 VDDH.n818 VDDH.n817 9.3005
R7074 VDDH.n831 VDDH.n742 9.3005
R7075 VDDH.n832 VDDH.n831 9.3005
R7076 VDDH.n816 VDDH.n814 9.3005
R7077 VDDH.n821 VDDH.n820 9.3005
R7078 VDDH.n815 VDDH.n741 9.3005
R7079 VDDH.n834 VDDH.n833 9.3005
R7080 VDDH.n835 VDDH.n737 9.3005
R7081 VDDH.n837 VDDH.n836 9.3005
R7082 VDDH.n804 VDDH.n803 9.3005
R7083 VDDH.n805 VDDH.n804 9.3005
R7084 VDDH.n791 VDDH.n790 9.3005
R7085 VDDH.n790 VDDH.n789 9.3005
R7086 VDDH.n807 VDDH.n806 9.3005
R7087 VDDH.n802 VDDH.n747 9.3005
R7088 VDDH.n801 VDDH.n800 9.3005
R7089 VDDH.n786 VDDH.n748 9.3005
R7090 VDDH.n793 VDDH.n792 9.3005
R7091 VDDH.n785 VDDH.n751 9.3005
R7092 VDDH.n783 VDDH.n782 9.3005
R7093 VDDH.n784 VDDH.n783 9.3005
R7094 VDDH.n766 VDDH.n765 9.3005
R7095 VDDH.n765 VDDH.n764 9.3005
R7096 VDDH.n779 VDDH.n752 9.3005
R7097 VDDH.n781 VDDH.n780 9.3005
R7098 VDDH.n754 VDDH.n753 9.3005
R7099 VDDH.n760 VDDH.n758 9.3005
R7100 VDDH.n81 VDDH.n80 9.3005
R7101 VDDH.n80 VDDH.n79 9.3005
R7102 VDDH.n89 VDDH.n88 9.3005
R7103 VDDH.n88 VDDH.n87 9.3005
R7104 VDDH.n725 VDDH.n724 9.3005
R7105 VDDH.n724 VDDH.n723 9.3005
R7106 VDDH.n703 VDDH.n702 9.3005
R7107 VDDH.n702 VDDH.n701 9.3005
R7108 VDDH.n83 VDDH.n82 9.3005
R7109 VDDH.n86 VDDH.n85 9.3005
R7110 VDDH.n75 VDDH.n73 9.3005
R7111 VDDH.n719 VDDH.n718 9.3005
R7112 VDDH.n722 VDDH.n721 9.3005
R7113 VDDH.n72 VDDH.n70 9.3005
R7114 VDDH.n727 VDDH.n726 9.3005
R7115 VDDH.n728 VDDH.n68 9.3005
R7116 VDDH.n729 VDDH.n67 9.3005
R7117 VDDH.n734 VDDH.n733 9.3005
R7118 VDDH.n78 VDDH.n57 9.3005
R7119 VDDH.n77 VDDH.n76 9.3005
R7120 VDDH.n575 VDDH.t273 9.29529
R7121 VDDH.n633 VDDH.n632 9.2505
R7122 VDDH.t495 VDDH.n633 9.2505
R7123 VDDH.n640 VDDH.n639 9.2505
R7124 VDDH.n639 VDDH.t441 9.2505
R7125 VDDH.n635 VDDH.n634 9.2505
R7126 VDDH.n634 VDDH.t495 9.2505
R7127 VDDH.n638 VDDH.n637 9.2505
R7128 VDDH.t441 VDDH.n638 9.2505
R7129 VDDH.n525 VDDH.n522 8.96925
R7130 VDDH.n525 VDDH.n524 8.96717
R7131 VDDH.t297 VDDH.n276 8.93316
R7132 VDDH.n472 VDDH.n464 8.81002
R7133 VDDH.n511 VDDH.n464 8.81002
R7134 VDDH.n485 VDDH.n465 8.81002
R7135 VDDH.n511 VDDH.n465 8.81002
R7136 VDDH.n513 VDDH.n512 8.81002
R7137 VDDH.n512 VDDH.n511 8.81002
R7138 VDDH.n510 VDDH.n456 8.81002
R7139 VDDH.n511 VDDH.n510 8.81002
R7140 VDDH.n451 VDDH.n450 8.55258
R7141 VDDH.n450 VDDH.n449 8.42133
R7142 VDDH.n503 VDDH.n474 8.40959
R7143 VDDH.n497 VDDH.n496 8.40959
R7144 VDDH.n161 VDDH.t251 8.13045
R7145 VDDH.t288 VDDH.t540 8.08818
R7146 VDDH.n439 VDDH.n230 7.70883
R7147 VDDH.n237 VDDH.n230 7.70883
R7148 VDDH.n437 VDDH.n436 7.70883
R7149 VDDH.n436 VDDH.n435 7.70883
R7150 VDDH.n268 VDDH.n267 7.70883
R7151 VDDH.n268 VDDH.n182 7.70883
R7152 VDDH.n263 VDDH.n257 7.70883
R7153 VDDH.n276 VDDH.n263 7.70883
R7154 VDDH.n281 VDDH.n256 7.70883
R7155 VDDH.n262 VDDH.n256 7.70883
R7156 VDDH.n431 VDDH.n229 7.70883
R7157 VDDH.n237 VDDH.n229 7.70883
R7158 VDDH.n434 VDDH.n433 7.70883
R7159 VDDH.n435 VDDH.n434 7.70883
R7160 VDDH.n264 VDDH.n244 7.70883
R7161 VDDH.n264 VDDH.n182 7.70883
R7162 VDDH.n275 VDDH.n274 7.70883
R7163 VDDH.n276 VDDH.n275 7.70883
R7164 VDDH.n258 VDDH.n255 7.70883
R7165 VDDH.n262 VDDH.n255 7.70883
R7166 VDDH.n536 VDDH.n535 7.70883
R7167 VDDH.n535 VDDH.n534 7.70883
R7168 VDDH.n286 VDDH.n249 7.70883
R7169 VDDH.n287 VDDH.n286 7.70883
R7170 VDDH.n254 VDDH.n246 7.70883
R7171 VDDH.n287 VDDH.n254 7.70883
R7172 VDDH.n533 VDDH.n215 7.70883
R7173 VDDH.n534 VDDH.n533 7.70883
R7174 VDDH.t275 VDDH.t245 7.60533
R7175 VDDH.t338 VDDH.n148 7.4369
R7176 VDDH.n685 VDDH.n111 7.11588
R7177 VDDH.n991 VDDH.n0 7.1155
R7178 VDDH.n272 VDDH.n271 6.85235
R7179 VDDH.n271 VDDH.n270 6.85235
R7180 VDDH.n243 VDDH.n242 6.85235
R7181 VDDH.n242 VDDH.n241 6.85235
R7182 VDDH.n283 VDDH.n282 6.85235
R7183 VDDH.n284 VDDH.n283 6.85235
R7184 VDDH.n239 VDDH.n232 6.85235
R7185 VDDH.n239 VDDH.n238 6.85235
R7186 VDDH.n441 VDDH.n440 6.85235
R7187 VDDH.n442 VDDH.n441 6.85235
R7188 VDDH.n279 VDDH.n278 6.85235
R7189 VDDH.n278 VDDH.n277 6.85235
R7190 VDDH.n143 VDDH.n93 6.85235
R7191 VDDH.n144 VDDH.n143 6.85235
R7192 VDDH.n167 VDDH.n166 6.85235
R7193 VDDH.n166 VDDH.n165 6.85235
R7194 VDDH.t455 VDDH.t297 6.63964
R7195 VDDH.n398 VDDH.n226 6.4005
R7196 VDDH.n392 VDDH.n391 6.4005
R7197 VDDH.n686 VDDH 6.4005
R7198 VDDH.n428 VDDH.n405 6.33487
R7199 VDDH.n428 VDDH.n427 6.33487
R7200 VDDH.n539 VDDH.n225 6.33487
R7201 VDDH.n548 VDDH.n539 6.33487
R7202 VDDH.t273 VDDH.t539 6.15679
R7203 VDDH.n767 VDDH.n759 6.13579
R7204 VDDH.n481 VDDH.n480 5.93473
R7205 VDDH.n1035 VDDH.n1034 5.78175
R7206 VDDH.n1040 VDDH.n1035 5.78175
R7207 VDDH.n1058 VDDH.n1057 5.78175
R7208 VDDH.n1059 VDDH.n1058 5.78175
R7209 VDDH.n1037 VDDH.n1036 5.78175
R7210 VDDH.n1040 VDDH.n1037 5.78175
R7211 VDDH.n1061 VDDH.n1060 5.78175
R7212 VDDH.n1060 VDDH.n1059 5.78175
R7213 VDDH.n1078 VDDH.n1077 5.78175
R7214 VDDH.n1079 VDDH.n1078 5.78175
R7215 VDDH.n1072 VDDH.n1071 5.78175
R7216 VDDH.n1071 VDDH.n1070 5.78175
R7217 VDDH.n1119 VDDH.n1118 5.78175
R7218 VDDH.n1118 VDDH.n1117 5.78175
R7219 VDDH.n1125 VDDH.n1124 5.78175
R7220 VDDH.n1126 VDDH.n1125 5.78175
R7221 VDDH.n1081 VDDH.n1080 5.78175
R7222 VDDH.n1080 VDDH.n1079 5.78175
R7223 VDDH.n1069 VDDH.n1068 5.78175
R7224 VDDH.n1070 VDDH.n1069 5.78175
R7225 VDDH.n1116 VDDH.n1115 5.78175
R7226 VDDH.n1117 VDDH.n1116 5.78175
R7227 VDDH.n1128 VDDH.n1127 5.78175
R7228 VDDH.n1127 VDDH.n1126 5.78175
R7229 VDDH.n1092 VDDH.n1091 5.78175
R7230 VDDH.n1091 VDDH.n1090 5.78175
R7231 VDDH.n1100 VDDH.n1099 5.78175
R7232 VDDH.n1101 VDDH.n1100 5.78175
R7233 VDDH.n1112 VDDH.n1111 5.78175
R7234 VDDH.n1111 VDDH.n1110 5.78175
R7235 VDDH.n1134 VDDH.n994 5.78175
R7236 VDDH.n1135 VDDH.n1134 5.78175
R7237 VDDH.n1089 VDDH.n1088 5.78175
R7238 VDDH.n1090 VDDH.n1089 5.78175
R7239 VDDH.n1103 VDDH.n1102 5.78175
R7240 VDDH.n1102 VDDH.n1101 5.78175
R7241 VDDH.n1109 VDDH.n1108 5.78175
R7242 VDDH.n1110 VDDH.n1109 5.78175
R7243 VDDH.n1137 VDDH.n1136 5.78175
R7244 VDDH.n1136 VDDH.n1135 5.78175
R7245 VDDH.n151 VDDH.n150 5.78175
R7246 VDDH.n415 VDDH.n414 5.60656
R7247 VDDH.n423 VDDH.n413 5.60656
R7248 VDDH.n509 VDDH.n466 5.28621
R7249 VDDH.n509 VDDH.n508 5.28621
R7250 VDDH.n515 VDDH.n457 5.28621
R7251 VDDH.n489 VDDH.n457 5.28621
R7252 VDDH.n534 VDDH.n531 5.17455
R7253 VDDH.n655 VDDH.n605 5.13939
R7254 VDDH.t75 VDDH.n655 5.13939
R7255 VDDH.n653 VDDH.n614 5.13939
R7256 VDDH.n653 VDDH.t500 5.13939
R7257 VDDH.n657 VDDH.n656 5.13939
R7258 VDDH.n656 VDDH.t75 5.13939
R7259 VDDH.n652 VDDH.n651 5.13939
R7260 VDDH.t500 VDDH.n652 5.13939
R7261 VDDH.n399 VDDH.n246 5.04292
R7262 VDDH.n393 VDDH.n289 5.04292
R7263 VDDH.n397 VDDH.n249 5.04292
R7264 VDDH.n390 VDDH.n189 5.04292
R7265 VDDH.n149 VDDH.t16 4.99224
R7266 VDDH.n529 VDDH.n520 4.89462
R7267 VDDH.n579 VDDH.n578 4.89462
R7268 VDDH.n345 VDDH.n344 4.89462
R7269 VDDH.n568 VDDH.n197 4.89462
R7270 VDDH.n551 VDDH.n215 4.89462
R7271 VDDH.n536 VDDH.n227 4.89462
R7272 VDDH.n290 VDDH.n190 4.89462
R7273 VDDH.n553 VDDH.n213 4.89462
R7274 VDDH.n670 VDDH.n669 4.89462
R7275 VDDH.n158 VDDH.n157 4.89462
R7276 VDDH.n162 VDDH.n123 4.89462
R7277 VDDH.n668 VDDH.n122 4.74409
R7278 VDDH.n122 VDDH.t56 4.74409
R7279 VDDH.n491 VDDH.n490 4.6255
R7280 VDDH.n490 VDDH.n489 4.6255
R7281 VDDH.n507 VDDH.n506 4.6255
R7282 VDDH.n508 VDDH.n507 4.6255
R7283 VDDH.n488 VDDH.n458 4.6255
R7284 VDDH.n489 VDDH.n488 4.6255
R7285 VDDH.n470 VDDH.n468 4.6255
R7286 VDDH.n508 VDDH.n468 4.6255
R7287 VDDH.n661 VDDH.n660 4.61883
R7288 VDDH.n277 VDDH.t291 4.58754
R7289 VDDH.n643 VDDH.n642 4.40526
R7290 VDDH.n644 VDDH.n643 4.40526
R7291 VDDH.n647 VDDH.n646 4.40526
R7292 VDDH.n646 VDDH.n645 4.40526
R7293 VDDH.n675 VDDH.n674 4.40526
R7294 VDDH.n674 VDDH.n673 4.40526
R7295 VDDH.n698 VDDH.n91 4.12585
R7296 VDDH.n241 VDDH.t54 4.10469
R7297 VDDH.n991 VDDH.n990 3.91654
R7298 VDDH.n967 VDDH 3.7711
R7299 VDDH VDDH.n968 3.7711
R7300 VDDH.n943 VDDH 3.7711
R7301 VDDH VDDH.n22 3.7711
R7302 VDDH.n839 VDDH 3.7711
R7303 VDDH.n840 VDDH 3.7711
R7304 VDDH VDDH.n841 3.7711
R7305 VDDH.n838 VDDH 3.7711
R7306 VDDH VDDH.n736 3.7711
R7307 VDDH.n990 VDDH 3.7711
R7308 VDDH.n993 VDDH.n991 3.41321
R7309 VDDH.n138 VDDH.n92 3.38392
R7310 VDDH.n170 VDDH.n132 3.36612
R7311 VDDH.n687 VDDH.n109 3.36414
R7312 VDDH.n161 VDDH.n109 3.36414
R7313 VDDH.n1050 VDDH.n1049 3.13609
R7314 VDDH.n1051 VDDH.n1050 3.13609
R7315 VDDH.n1053 VDDH.n1052 3.13609
R7316 VDDH.n1052 VDDH.n1051 3.13609
R7317 VDDH.n132 VDDH.n131 3.1255
R7318 VDDH.n141 VDDH.n140 2.93701
R7319 VDDH.n148 VDDH.n141 2.93701
R7320 VDDH.n696 VDDH.n94 2.93701
R7321 VDDH.n148 VDDH.n94 2.93701
R7322 VDDH.n770 VDDH.t474 2.8822
R7323 VDDH.n775 VDDH.t0 2.8822
R7324 VDDH.n795 VDDH.t523 2.8822
R7325 VDDH.t371 VDDH.n745 2.8822
R7326 VDDH.n811 VDDH.t406 2.8822
R7327 VDDH.n824 VDDH.t352 2.8822
R7328 VDDH.n852 VDDH.t354 2.8822
R7329 VDDH.t348 VDDH.n49 2.8822
R7330 VDDH.t309 VDDH.n867 2.8822
R7331 VDDH.n879 VDDH.t328 2.8822
R7332 VDDH.n904 VDDH.t67 2.8822
R7333 VDDH.n909 VDDH.t535 2.8822
R7334 VDDH.n929 VDDH.t528 2.8822
R7335 VDDH.n934 VDDH.t79 2.8822
R7336 VDDH.n1139 VDDH.n993 2.55404
R7337 VDDH.t279 VDDH.t326 2.53544
R7338 VDDH.n421 VDDH.n420 2.44894
R7339 VDDH.n688 VDDH.n108 2.39269
R7340 VDDH VDDH.n1139 2.33717
R7341 VDDH.n696 VDDH.n695 2.25932
R7342 VDDH.n993 VDDH.n992 2.23833
R7343 VDDH.t287 VDDH.t327 2.0526
R7344 VDDH.t559 VDDH.t277 2.0526
R7345 VDDH.n424 VDDH.n411 2.04581
R7346 VDDH.n420 VDDH.n419 2.04581
R7347 VDDH.n684 VDDH.n108 1.99425
R7348 VDDH.n425 VDDH.n424 1.78175
R7349 VDDH.n603 VDDH.n602 1.75795
R7350 VDDH.n690 VDDH.n103 1.66612
R7351 VDDH.n767 VDDH.n766 1.60272
R7352 VDDH.n645 VDDH.n644 1.563
R7353 VDDH.n101 VDDH.n100 1.48331
R7354 VDDH.n735 VDDH 1.47967
R7355 VDDH.n259 VDDH 1.47077
R7356 VDDH VDDH.n273 1.47077
R7357 VDDH.n430 VDDH 1.47077
R7358 VDDH VDDH.n432 1.47077
R7359 VDDH.n131 VDDH.n91 1.4624
R7360 VDDH.n502 VDDH.n501 1.45988
R7361 VDDH.n499 VDDH.n498 1.45988
R7362 VDDH.n516 VDDH.n199 1.43637
R7363 VDDH.n460 VDDH.n199 1.40704
R7364 VDDH.n517 VDDH.n516 1.388
R7365 VDDH.n178 VDDH.n176 1.3811
R7366 VDDH.n181 VDDH.n178 1.3811
R7367 VDDH.n569 VDDH.n196 1.3811
R7368 VDDH.n196 VDDH.n181 1.3811
R7369 VDDH.n429 VDDH.n185 1.3811
R7370 VDDH.n574 VDDH.n185 1.3811
R7371 VDDH.n214 VDDH.n186 1.3811
R7372 VDDH.n574 VDDH.n186 1.3811
R7373 VDDH.n573 VDDH.n572 1.3811
R7374 VDDH.n574 VDDH.n573 1.3811
R7375 VDDH.n684 VDDH.n683 1.3755
R7376 VDDH.n538 VDDH.n184 1.37087
R7377 VDDH.n574 VDDH.n184 1.37087
R7378 VDDH.n389 VDDH.n183 1.37087
R7379 VDDH.n574 VDDH.n183 1.37087
R7380 VDDH.n527 VDDH.n526 1.36079
R7381 VDDH.n526 VDDH.n181 1.36079
R7382 VDDH.n480 VDDH.n460 1.32758
R7383 VDDH.n549 VDDH.n216 1.29217
R7384 VDDH.n550 VDDH.n212 1.29217
R7385 VDDH.n550 VDDH.n549 1.29217
R7386 VDDH.n519 VDDH.n198 1.24425
R7387 VDDH.n567 VDDH.n198 1.24425
R7388 VDDH.n498 VDDH 1.238
R7389 VDDH.n138 VDDH.n102 1.19112
R7390 VDDH.n692 VDDH.n691 1.163
R7391 VDDH.n157 VDDH.n103 1.163
R7392 VDDH.n426 VDDH.n216 1.15755
R7393 VDDH.n139 VDDH.n138 1.14843
R7394 VDDH.n517 VDDH.n453 1.14581
R7395 VDDH.n689 VDDH.n688 1.13331
R7396 VDDH.n102 VDDH.n101 1.08019
R7397 VDDH.n582 VDDH.n173 1.01113
R7398 VDDH.n679 VDDH.n678 0.985808
R7399 VDDH.n324 VDDH.n322 0.947451
R7400 VDDH.n337 VDDH.n336 0.947451
R7401 VDDH.n128 VDDH.n125 0.947451
R7402 VDDH.n476 VDDH.n173 0.922375
R7403 VDDH.n326 VDDH.n324 0.91925
R7404 VDDH.n328 VDDH.n326 0.91925
R7405 VDDH.n330 VDDH.n328 0.91925
R7406 VDDH.n336 VDDH.n335 0.91925
R7407 VDDH.n335 VDDH.n334 0.91925
R7408 VDDH.n334 VDDH.n333 0.91925
R7409 VDDH.n333 VDDH.n332 0.91925
R7410 VDDH.n332 VDDH.n330 0.91925
R7411 VDDH.n378 VDDH.n375 0.91925
R7412 VDDH.n381 VDDH.n378 0.91925
R7413 VDDH.n384 VDDH.n381 0.91925
R7414 VDDH.n387 VDDH.n384 0.91925
R7415 VDDH.n371 VDDH.n370 0.91925
R7416 VDDH.n370 VDDH.n369 0.91925
R7417 VDDH.n369 VDDH.n368 0.91925
R7418 VDDH.n368 VDDH.n367 0.91925
R7419 VDDH.n172 VDDH.n0 0.914875
R7420 VDDH.n677 VDDH.n118 0.873938
R7421 VDDH.n477 VDDH.n476 0.863521
R7422 VDDH.n736 VDDH.n735 0.8605
R7423 VDDH.n555 VDDH.n554 0.837038
R7424 VDDH.n554 VDDH.n212 0.837038
R7425 VDDH.n565 VDDH.n200 0.837038
R7426 VDDH.n555 VDDH.n200 0.837038
R7427 VDDH.n662 VDDH.n112 0.816125
R7428 VDDH.n682 VDDH.n112 0.816125
R7429 VDDH.n483 VDDH.n473 0.7755
R7430 VDDH.n500 VDDH.n475 0.7755
R7431 VDDH.n422 VDDH.n421 0.7755
R7432 VDDH.n412 VDDH.n410 0.7755
R7433 VDDH.n477 VDDH.n453 0.761438
R7434 VDDH.n667 VDDH.n666 0.753625
R7435 VDDH.n405 VDDH.n400 0.737359
R7436 VDDH.n237 VDDH.t50 0.724769
R7437 VDDH.n425 VDDH.n410 0.667688
R7438 VDDH.n523 VDDH.n198 0.63175
R7439 VDDH.n100 VDDH.n92 0.6255
R7440 VDDH.n480 VDDH.n479 0.623
R7441 VDDH.n200 VDDH.n190 0.6205
R7442 VDDH.n554 VDDH.n553 0.6205
R7443 VDDH.n394 VDDH.n393 0.6205
R7444 VDDH.n347 VDDH.n189 0.6205
R7445 VDDH.n669 VDDH.n112 0.6205
R7446 VDDH.n169 VDDH.n123 0.6205
R7447 VDDH.n838 VDDH.n736 0.61925
R7448 VDDH.n841 VDDH.n838 0.61925
R7449 VDDH.n841 VDDH.n840 0.61925
R7450 VDDH.n840 VDDH.n839 0.61925
R7451 VDDH.n839 VDDH.n22 0.61925
R7452 VDDH.n943 VDDH.n22 0.61925
R7453 VDDH.n968 VDDH.n943 0.61925
R7454 VDDH.n968 VDDH.n967 0.61925
R7455 VDDH.n690 VDDH.n689 0.61925
R7456 VDDH.n735 VDDH 0.617892
R7457 VDDH.t268 VDDH.t558 0.604058
R7458 VDDH.n479 VDDH 0.6015
R7459 VDDH.n518 VDDH.n452 0.58175
R7460 VDDH.n549 VDDH.n548 0.577063
R7461 VDDH.n661 VDDH.n172 0.571125
R7462 VDDH.n521 VDDH.n175 0.56925
R7463 VDDH.n967 VDDH 0.56425
R7464 VDDH.t163 VDDH.t89 0.562896
R7465 VDDH.n520 VDDH.n519 0.547559
R7466 VDDH.n568 VDDH.n567 0.547559
R7467 VDDH.n346 VDDH.n345 0.547559
R7468 VDDH.n580 VDDH.n579 0.547559
R7469 VDDH.n427 VDDH.n426 0.545851
R7470 VDDH.n502 VDDH.n481 0.54401
R7471 VDDH.n666 VDDH.n665 0.534794
R7472 VDDH.n375 VDDH.n372 0.528735
R7473 VDDH.n367 VDDH.n366 0.528735
R7474 VDDH.n712 VDDH.n711 0.517167
R7475 VDDH.n706 VDDH.n90 0.517167
R7476 VDDH.n717 VDDH.n716 0.517167
R7477 VDDH.n245 VDDH.n225 0.516125
R7478 VDDH.n137 VDDH.n118 0.516125
R7479 VDDH.n358 VDDH.n357 0.51137
R7480 VDDH.n357 VDDH.n356 0.51137
R7481 VDDH.n356 VDDH.n193 0.51137
R7482 VDDH.n571 VDDH.n193 0.51137
R7483 VDDH.n205 VDDH.n195 0.51137
R7484 VDDH.n206 VDDH.n205 0.51137
R7485 VDDH.n207 VDDH.n206 0.51137
R7486 VDDH.n359 VDDH.n358 0.495392
R7487 VDDH.n208 VDDH.n207 0.495392
R7488 VDDH.n570 VDDH.n195 0.494386
R7489 VDDH.n460 VDDH.n459 0.49364
R7490 VDDH.n455 VDDH.n454 0.49364
R7491 VDDH.n131 VDDH.n0 0.475677
R7492 VDDH.n663 VDDH.n661 0.475145
R7493 VDDH.n388 VDDH.n371 0.459875
R7494 VDDH.n388 VDDH.n387 0.459875
R7495 VDDH.n513 VDDH.n460 0.443357
R7496 VDDH.n456 VDDH.n455 0.443357
R7497 VDDH.n581 VDDH.n174 0.440083
R7498 VDDH.n503 VDDH.n502 0.423227
R7499 VDDH.n498 VDDH.n497 0.423227
R7500 VDDH.n691 VDDH.n690 0.40675
R7501 VDDH.n551 VDDH.n550 0.404848
R7502 VDDH.n227 VDDH.n216 0.404848
R7503 VDDH.n400 VDDH.n399 0.404848
R7504 VDDH.n397 VDDH.n396 0.404848
R7505 VDDH.n500 VDDH.n499 0.403625
R7506 VDDH.n501 VDDH.n500 0.403625
R7507 VDDH.n484 VDDH.n483 0.403625
R7508 VDDH.n483 VDDH.n482 0.403625
R7509 VDDH.n421 VDDH.n411 0.403625
R7510 VDDH.n419 VDDH.n410 0.403625
R7511 VDDH.n685 VDDH.n684 0.3725
R7512 VDDH.t137 VDDH.t141 0.362819
R7513 VDDH.t457 VDDH.t83 0.362819
R7514 VDDH.t82 VDDH.t456 0.362819
R7515 VDDH.n93 VDDH.n91 0.358192
R7516 VDDH.n168 VDDH.n167 0.358192
R7517 VDDH.n341 VDDH.n340 0.346537
R7518 VDDH.n560 VDDH.n559 0.346537
R7519 VDDH.n314 VDDH.n210 0.346537
R7520 VDDH.n363 VDDH.n362 0.346537
R7521 VDDH.n101 VDDH.n95 0.3005
R7522 VDDH.n170 VDDH.n169 0.300179
R7523 VDDH.n424 VDDH.n423 0.291125
R7524 VDDH.n420 VDDH.n414 0.291125
R7525 VDDH.n318 VDDH.n315 0.288543
R7526 VDDH.n318 VDDH.n316 0.288543
R7527 VDDH.n306 VDDH.n303 0.288543
R7528 VDDH.n306 VDDH.n304 0.288543
R7529 VDDH.n404 VDDH.n401 0.288543
R7530 VDDH.n404 VDDH.n402 0.288543
R7531 VDDH.n409 VDDH.n406 0.288543
R7532 VDDH.n409 VDDH.n407 0.288543
R7533 VDDH.n224 VDDH.n221 0.288543
R7534 VDDH.n224 VDDH.n222 0.288543
R7535 VDDH.n220 VDDH.n217 0.288543
R7536 VDDH.n220 VDDH.n218 0.288543
R7537 VDDH.n547 VDDH.n544 0.288543
R7538 VDDH.n547 VDDH.n545 0.288543
R7539 VDDH.n543 VDDH.n540 0.288543
R7540 VDDH.n543 VDDH.n541 0.288543
R7541 VDDH.n566 VDDH.n565 0.285826
R7542 VDDH.n450 VDDH.n173 0.284771
R7543 VDDH.n582 VDDH.n581 0.283341
R7544 VDDH.n476 VDDH.n452 0.275396
R7545 VDDH.n479 VDDH.n466 0.274029
R7546 VDDH.n516 VDDH.n515 0.274029
R7547 VDDH.n519 VDDH.n518 0.273417
R7548 VDDH.n566 VDDH.n199 0.273356
R7549 VDDH.n324 VDDH.n323 0.255835
R7550 VDDH.n326 VDDH.n325 0.255835
R7551 VDDH.n328 VDDH.n327 0.255835
R7552 VDDH.n330 VDDH.n329 0.255835
R7553 VDDH.n336 VDDH.n308 0.255835
R7554 VDDH.n335 VDDH.n309 0.255835
R7555 VDDH.n334 VDDH.n310 0.255835
R7556 VDDH.n333 VDDH.n311 0.255835
R7557 VDDH.n332 VDDH.n331 0.255835
R7558 VDDH.n375 VDDH.n373 0.255835
R7559 VDDH.n375 VDDH.n374 0.255835
R7560 VDDH.n378 VDDH.n376 0.255835
R7561 VDDH.n378 VDDH.n377 0.255835
R7562 VDDH.n381 VDDH.n379 0.255835
R7563 VDDH.n381 VDDH.n380 0.255835
R7564 VDDH.n384 VDDH.n382 0.255835
R7565 VDDH.n384 VDDH.n383 0.255835
R7566 VDDH.n387 VDDH.n385 0.255835
R7567 VDDH.n387 VDDH.n386 0.255835
R7568 VDDH.n371 VDDH.n292 0.255835
R7569 VDDH.n371 VDDH.n293 0.255835
R7570 VDDH.n370 VDDH.n294 0.255835
R7571 VDDH.n370 VDDH.n295 0.255835
R7572 VDDH.n369 VDDH.n296 0.255835
R7573 VDDH.n369 VDDH.n297 0.255835
R7574 VDDH.n368 VDDH.n298 0.255835
R7575 VDDH.n368 VDDH.n299 0.255835
R7576 VDDH.n367 VDDH.n300 0.255835
R7577 VDDH.n367 VDDH.n301 0.255835
R7578 VDDH.n678 VDDH.n116 0.255835
R7579 VDDH.n118 VDDH.n117 0.255835
R7580 VDDH.n125 VDDH.n124 0.255835
R7581 VDDH.n666 VDDH.n126 0.255835
R7582 VDDH.n172 VDDH.n171 0.251034
R7583 VDDH.n452 VDDH.n451 0.2505
R7584 VDDH.n683 VDDH.n682 0.241125
R7585 VDDH.n668 VDDH.n667 0.238962
R7586 VDDH.n339 VDDH.n306 0.232207
R7587 VDDH.n319 VDDH.n318 0.232207
R7588 VDDH.n322 VDDH.n321 0.227634
R7589 VDDH.n340 VDDH.n339 0.227634
R7590 VDDH.n337 VDDH.n307 0.227634
R7591 VDDH.n319 VDDH.n314 0.227634
R7592 VDDH.n128 VDDH.n127 0.227634
R7593 VDDH.n677 VDDH.n676 0.227329
R7594 VDDH.n171 VDDH.n170 0.226462
R7595 VDDH.n571 VDDH.n191 0.225348
R7596 VDDH.n207 VDDH.n202 0.225348
R7597 VDDH.n206 VDDH.n203 0.225348
R7598 VDDH.n205 VDDH.n204 0.225348
R7599 VDDH.n195 VDDH.n194 0.225348
R7600 VDDH.n193 VDDH.n192 0.225348
R7601 VDDH.n356 VDDH.n355 0.225348
R7602 VDDH.n357 VDDH.n354 0.225348
R7603 VDDH.n358 VDDH.n353 0.225348
R7604 VDDH.n598 VDDH.n587 0.224528
R7605 VDDH VDDH.n484 0.222375
R7606 VDDH.n396 VDDH.n395 0.221734
R7607 VDDH.n396 VDDH.n245 0.221734
R7608 VDDH.n400 VDDH.n245 0.221734
R7609 VDDH.n700 VDDH.n699 0.218612
R7610 VDDH.n710 VDDH.n709 0.218612
R7611 VDDH.n708 VDDH.n707 0.218612
R7612 VDDH.n705 VDDH.n704 0.218612
R7613 VDDH.n169 VDDH.n168 0.214709
R7614 VDDH.n482 VDDH.n481 0.20675
R7615 VDDH.n698 VDDH.n697 0.205663
R7616 VDDH.n405 VDDH.n404 0.204006
R7617 VDDH.n427 VDDH.n409 0.204006
R7618 VDDH.n225 VDDH.n220 0.204006
R7619 VDDH.n225 VDDH.n224 0.204006
R7620 VDDH.n548 VDDH.n543 0.204006
R7621 VDDH.n548 VDDH.n547 0.204006
R7622 VDDH.n604 VDDH.n582 0.198625
R7623 VDDH VDDH.n13 0.195324
R7624 VDDH VDDH.n21 0.195324
R7625 VDDH VDDH.n966 0.195324
R7626 VDDH VDDH.n989 0.195324
R7627 VDDH.n312 VDDH.n212 0.192606
R7628 VDDH.n699 VDDH.n698 0.190551
R7629 VDDH.n556 VDDH.n555 0.186547
R7630 VDDH.n306 VDDH.n305 0.186476
R7631 VDDH.n404 VDDH.n403 0.186476
R7632 VDDH.n409 VDDH.n408 0.186476
R7633 VDDH.n220 VDDH.n219 0.186476
R7634 VDDH.n224 VDDH.n223 0.186476
R7635 VDDH.n543 VDDH.n542 0.186476
R7636 VDDH.n547 VDDH.n546 0.186476
R7637 VDDH.n318 VDDH.n317 0.186476
R7638 VDDH.n137 VDDH.n136 0.185122
R7639 VDDH.n348 VDDH.n346 0.182662
R7640 VDDH.n688 VDDH.n687 0.172722
R7641 VDDH.n359 VDDH.n352 0.168945
R7642 VDDH.n364 VDDH.n341 0.168945
R7643 VDDH.n208 VDDH.n201 0.168945
R7644 VDDH.n561 VDDH.n560 0.168945
R7645 VDDH.n559 VDDH.n558 0.168945
R7646 VDDH.n558 VDDH.n210 0.168945
R7647 VDDH.n362 VDDH.n361 0.168945
R7648 VDDH.n364 VDDH.n363 0.168945
R7649 VDDH.n679 VDDH.n115 0.168945
R7650 VDDH.n689 VDDH.n105 0.168674
R7651 VDDH.n108 VDDH.n107 0.168674
R7652 VDDH.n680 VDDH.n114 0.168674
R7653 VDDH.n581 VDDH.n580 0.166549
R7654 VDDH.n580 VDDH.n175 0.166549
R7655 VDDH.n346 VDDH.n175 0.166549
R7656 VDDH.n667 VDDH.n125 0.166125
R7657 VDDH.n348 VDDH.n347 0.161065
R7658 VDDH.n682 VDDH.n681 0.159794
R7659 VDDH.n680 VDDH.n679 0.153097
R7660 VDDH.n140 VDDH.n132 0.152959
R7661 VDDH.n697 VDDH.n696 0.152959
R7662 VDDH.n518 VDDH 0.151176
R7663 VDDH.n347 VDDH.n251 0.147467
R7664 VDDH.n394 VDDH.n251 0.147467
R7665 VDDH.n395 VDDH.n394 0.147467
R7666 VDDH.n709 VDDH 0.145908
R7667 VDDH.n704 VDDH 0.145908
R7668 VDDH.n395 VDDH.n250 0.131669
R7669 VDDH.n711 VDDH.n700 0.129327
R7670 VDDH.n707 VDDH.n706 0.129327
R7671 VDDH.n342 VDDH.n251 0.12561
R7672 VDDH.n785 VDDH 0.1255
R7673 VDDH VDDH.n837 0.1255
R7674 VDDH.n842 VDDH 0.1255
R7675 VDDH.n871 VDDH 0.1255
R7676 VDDH.n900 VDDH 0.1255
R7677 VDDH.n925 VDDH 0.1255
R7678 VDDH.n287 VDDH.n284 0.121212
R7679 VDDH.n575 VDDH.n182 0.121212
R7680 VDDH.t107 VDDH.t163 0.112979
R7681 VDDH VDDH.n517 0.112662
R7682 VDDH.n660 VDDH.n604 0.111125
R7683 VDDH VDDH.n708 0.108918
R7684 VDDH.n302 VDDH.n250 0.105208
R7685 VDDH.n313 VDDH.n312 0.105208
R7686 VDDH.n681 VDDH.n680 0.105208
R7687 VDDH.n130 VDDH.n129 0.105208
R7688 VDDH.n665 VDDH.n664 0.105208
R7689 VDDH.n558 VDDH.n211 0.10357
R7690 VDDH.n558 VDDH.n557 0.10357
R7691 VDDH.n364 VDDH.n343 0.10357
R7692 VDDH.n365 VDDH.n364 0.10357
R7693 VDDH.n209 VDDH.n208 0.0915853
R7694 VDDH.n561 VDDH.n209 0.0915853
R7695 VDDH.n562 VDDH.n561 0.0915853
R7696 VDDH.n361 VDDH.n360 0.0915853
R7697 VDDH.n360 VDDH.n359 0.0915853
R7698 VDDH.n711 VDDH.n710 0.0897857
R7699 VDDH.n706 VDDH.n705 0.0897857
R7700 VDDH.n565 VDDH.n564 0.087051
R7701 VDDH.n322 VDDH.n320 0.086539
R7702 VDDH.n320 VDDH.n319 0.086539
R7703 VDDH.n339 VDDH.n302 0.086539
R7704 VDDH.n339 VDDH.n338 0.086539
R7705 VDDH.n338 VDDH.n337 0.086539
R7706 VDDH.n319 VDDH.n313 0.086539
R7707 VDDH.n129 VDDH.n128 0.086539
R7708 VDDH.n168 VDDH.n139 0.0865043
R7709 VDDH.n139 VDDH.n137 0.078625
R7710 VDDH.n429 VDDH.n428 0.0731563
R7711 VDDH.n332 VDDH.n214 0.0731563
R7712 VDDH.n539 VDDH.n538 0.0731563
R7713 VDDH.n572 VDDH.n571 0.0731563
R7714 VDDH.n389 VDDH.n388 0.0731563
R7715 VDDH.n450 VDDH.n176 0.072593
R7716 VDDH.n527 VDDH.n525 0.072593
R7717 VDDH.n570 VDDH.n569 0.072593
R7718 VDDH.n372 VDDH.n211 0.0712237
R7719 VDDH.n557 VDDH.n556 0.0712237
R7720 VDDH.n343 VDDH.n342 0.0712237
R7721 VDDH.n366 VDDH.n365 0.0712237
R7722 VDDH.n361 VDDH.n351 0.0707519
R7723 VDDH.n350 VDDH.n349 0.063
R7724 VDDH.n603 VDDH 0.0609167
R7725 VDDH.n564 VDDH.n563 0.0605775
R7726 VDDH.n349 VDDH.n348 0.0605565
R7727 VDDH.n448 VDDH.n174 0.0575652
R7728 VDDH.n449 VDDH.n448 0.0575652
R7729 VDDH.n990 VDDH 0.0555
R7730 VDDH.n781 VDDH.n753 0.047375
R7731 VDDH.n792 VDDH.n785 0.047375
R7732 VDDH.n802 VDDH.n801 0.047375
R7733 VDDH.n837 VDDH.n737 0.047375
R7734 VDDH.n820 VDDH.n815 0.047375
R7735 VDDH.n849 VDDH.n842 0.047375
R7736 VDDH.n859 VDDH.n858 0.047375
R7737 VDDH.n872 VDDH.n871 0.047375
R7738 VDDH.n888 VDDH.n887 0.047375
R7739 VDDH.n900 VDDH.n899 0.047375
R7740 VDDH.n914 VDDH.n32 0.047375
R7741 VDDH.n925 VDDH.n924 0.047375
R7742 VDDH.n939 VDDH.n24 0.047375
R7743 VDDH.n972 VDDH.n13 0.047375
R7744 VDDH.n952 VDDH.n21 0.047375
R7745 VDDH.n966 VDDH.n7 0.047375
R7746 VDDH.n989 VDDH.n2 0.047375
R7747 VDDH.n678 VDDH.n677 0.0458125
R7748 VDDH.n664 VDDH.n663 0.0386493
R7749 VDDH.n137 VDDH.n134 0.0379178
R7750 VDDH VDDH.n725 0.0363146
R7751 VDDH VDDH.n81 0.0338567
R7752 VDDH.n766 VDDH.n760 0.0322383
R7753 VDDH.n782 VDDH.n752 0.0322383
R7754 VDDH.n791 VDDH.n786 0.0322383
R7755 VDDH.n806 VDDH.n803 0.0322383
R7756 VDDH.n833 VDDH.n742 0.0322383
R7757 VDDH.n819 VDDH.n816 0.0322383
R7758 VDDH.n848 VDDH.n843 0.0322383
R7759 VDDH.n863 VDDH.n860 0.0322383
R7760 VDDH.n876 VDDH.n873 0.0322383
R7761 VDDH.n886 VDDH.n883 0.0322383
R7762 VDDH.n898 VDDH.n39 0.0322383
R7763 VDDH.n915 VDDH.n31 0.0322383
R7764 VDDH.n923 VDDH.n918 0.0322383
R7765 VDDH.n940 VDDH.n23 0.0322383
R7766 VDDH.n971 VDDH.n20 0.0322383
R7767 VDDH.n953 VDDH.n944 0.0322383
R7768 VDDH.n961 VDDH.n958 0.0322383
R7769 VDDH.n985 VDDH.n982 0.0322383
R7770 VDDH.n718 VDDH.n71 0.0282388
R7771 VDDH.n82 VDDH.n74 0.0282388
R7772 VDDH.n734 VDDH.n56 0.0282388
R7773 VDDH.n683 VDDH 0.0270625
R7774 VDDH VDDH.n717 0.0268343
R7775 VDDH.n726 VDDH.n69 0.0257809
R7776 VDDH VDDH.n753 0.0239375
R7777 VDDH.n801 VDDH 0.0239375
R7778 VDDH.n815 VDDH 0.0239375
R7779 VDDH.n858 VDDH 0.0239375
R7780 VDDH.n888 VDDH 0.0239375
R7781 VDDH VDDH.n32 0.0239375
R7782 VDDH VDDH.n24 0.0239375
R7783 VDDH.n701 VDDH.n67 0.023323
R7784 VDDH.n723 VDDH.n70 0.023323
R7785 VDDH.n87 VDDH.n73 0.023323
R7786 VDDH.n79 VDDH.n77 0.023323
R7787 VDDH.n351 VDDH.n350 0.0213333
R7788 VDDH.n969 VDDH 0.0205195
R7789 VDDH VDDH.n955 0.0205195
R7790 VDDH.n960 VDDH 0.0205195
R7791 VDDH.n984 VDDH 0.0205195
R7792 VDDH.n764 VDDH.n763 0.0200312
R7793 VDDH.n789 VDDH.n788 0.0200312
R7794 VDDH.n832 VDDH.n830 0.0200312
R7795 VDDH.n846 VDDH.n845 0.0200312
R7796 VDDH.n875 VDDH.n43 0.0200312
R7797 VDDH.n896 VDDH.n895 0.0200312
R7798 VDDH.n921 VDDH.n920 0.0200312
R7799 VDDH.n663 VDDH.n662 0.017691
R7800 VDDH.n571 VDDH.n570 0.0174837
R7801 VDDH.n726 VDDH 0.0173539
R7802 VDDH.n718 VDDH 0.0173539
R7803 VDDH.n82 VDDH 0.0173539
R7804 VDDH VDDH.n734 0.0173539
R7805 VDDH VDDH.n703 0.0161716
R7806 VDDH.n782 VDDH.n781 0.0156367
R7807 VDDH VDDH.n784 0.0156367
R7808 VDDH.n792 VDDH.n791 0.0156367
R7809 VDDH.n803 VDDH.n802 0.0156367
R7810 VDDH.n805 VDDH 0.0156367
R7811 VDDH.n742 VDDH.n737 0.0156367
R7812 VDDH.n820 VDDH.n819 0.0156367
R7813 VDDH.n817 VDDH 0.0156367
R7814 VDDH.n849 VDDH.n848 0.0156367
R7815 VDDH.n860 VDDH.n859 0.0156367
R7816 VDDH.n862 VDDH 0.0156367
R7817 VDDH.n873 VDDH.n872 0.0156367
R7818 VDDH.n887 VDDH.n886 0.0156367
R7819 VDDH.n884 VDDH 0.0156367
R7820 VDDH.n899 VDDH.n898 0.0156367
R7821 VDDH.n915 VDDH.n914 0.0156367
R7822 VDDH VDDH.n917 0.0156367
R7823 VDDH.n924 VDDH.n923 0.0156367
R7824 VDDH.n940 VDDH.n939 0.0156367
R7825 VDDH VDDH.n942 0.0156367
R7826 VDDH.n972 VDDH.n971 0.0156367
R7827 VDDH.n953 VDDH.n952 0.0156367
R7828 VDDH.n958 VDDH.n7 0.0156367
R7829 VDDH.n982 VDDH.n2 0.0156367
R7830 VDDH.n478 VDDH.n477 0.013
R7831 VDDH.n701 VDDH.n68 0.0113848
R7832 VDDH.n723 VDDH.n722 0.0113848
R7833 VDDH.n87 VDDH.n86 0.0113848
R7834 VDDH.n79 VDDH.n78 0.0113848
R7835 VDDH.n105 VDDH.n104 0.00995724
R7836 VDDH.n107 VDDH.n106 0.00995724
R7837 VDDH.n114 VDDH.n113 0.00995724
R7838 VDDH.n134 VDDH.n133 0.00995724
R7839 VDDH.n136 VDDH.n135 0.00995724
R7840 VDDH.n69 VDDH.n68 0.00892697
R7841 VDDH.n455 VDDH.n453 0.00812195
R7842 VDDH.n717 VDDH.n89 0.00752247
R7843 VDDH VDDH.n478 0.007
R7844 VDDH.n722 VDDH.n71 0.0064691
R7845 VDDH.n86 VDDH.n74 0.0064691
R7846 VDDH.n78 VDDH.n56 0.0064691
R7847 VDDH.n697 VDDH.n92 0.00457609
R7848 VDDH.n478 VDDH 0.0045625
R7849 VDDH.n764 VDDH.n760 0.00391797
R7850 VDDH.n784 VDDH.n752 0.00391797
R7851 VDDH.n789 VDDH.n786 0.00391797
R7852 VDDH.n806 VDDH.n805 0.00391797
R7853 VDDH.n833 VDDH.n832 0.00391797
R7854 VDDH.n817 VDDH.n816 0.00391797
R7855 VDDH.n846 VDDH.n843 0.00391797
R7856 VDDH.n863 VDDH.n862 0.00391797
R7857 VDDH.n876 VDDH.n875 0.00391797
R7858 VDDH.n884 VDDH.n883 0.00391797
R7859 VDDH.n896 VDDH.n39 0.00391797
R7860 VDDH.n917 VDDH.n31 0.00391797
R7861 VDDH.n921 VDDH.n918 0.00391797
R7862 VDDH.n942 VDDH.n23 0.00391797
R7863 VDDH.n969 VDDH.n20 0.00391797
R7864 VDDH.n955 VDDH.n944 0.00391797
R7865 VDDH.n961 VDDH.n960 0.00391797
R7866 VDDH.n985 VDDH.n984 0.00391797
R7867 VDDH.n703 VDDH.n67 0.00295787
R7868 VDDH.n725 VDDH.n70 0.00295787
R7869 VDDH.n89 VDDH.n73 0.00295787
R7870 VDDH.n81 VDDH.n77 0.00295787
R7871 VDDH.n563 VDDH.n562 0.00292248
R7872 VDDH.n524 VDDH.n523 0.00258333
R7873 VDDH.n522 VDDH.n521 0.00258333
R7874 VDDH.n763 VDDH 0.000988281
R7875 VDDH.n788 VDDH 0.000988281
R7876 VDDH.n830 VDDH 0.000988281
R7877 VDDH.n845 VDDH 0.000988281
R7878 VDDH VDDH.n43 0.000988281
R7879 VDDH.n895 VDDH 0.000988281
R7880 VDDH.n920 VDDH 0.000988281
R7881 a_23629_18133.n0 a_23629_18133.t5 241.998
R7882 a_23629_18133.n2 a_23629_18133.t1 239.899
R7883 a_23629_18133.n2 a_23629_18133.t4 239.264
R7884 a_23629_18133.n1 a_23629_18133.t2 239.065
R7885 a_23629_18133.n0 a_23629_18133.t3 239.065
R7886 a_23629_18133.t0 a_23629_18133.n3 239.065
R7887 a_23629_18133.n1 a_23629_18133.n0 2.93383
R7888 a_23629_18133.n3 a_23629_18133.n1 2.93383
R7889 a_23629_18133.n3 a_23629_18133.n2 2.7755
R7890 a_21927_20174.t0 a_21927_20174.n1 251.352
R7891 a_21927_20174.n0 a_21927_20174.t3 248.684
R7892 a_21927_20174.n1 a_21927_20174.t2 241.264
R7893 a_21927_20174.n0 a_21927_20174.t1 239.282
R7894 a_21927_20174.n1 a_21927_20174.n0 2.66925
R7895 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2.n0 238.046
R7896 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2.t2 10.7009
R7897 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2.t1 10.5739
R7898 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.n0 240.27
R7899 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.t1 10.6692
R7900 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.t2 10.5285
R7901 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t5 222.043
R7902 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t3 222.043
R7903 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n27 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t1 140.061
R7904 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n28 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t0 139.566
R7905 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t12 126.178
R7906 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t28 124.9
R7907 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t21 124.9
R7908 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t22 124.9
R7909 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t9 124.9
R7910 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t16 124.9
R7911 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t26 124.9
R7912 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t10 124.9
R7913 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t19 124.9
R7914 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t27 124.9
R7915 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t14 124.9
R7916 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t20 124.9
R7917 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t7 124.9
R7918 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t15 124.9
R7919 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t25 124.9
R7920 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t8 124.9
R7921 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t6 124.9
R7922 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t13 124.9
R7923 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t23 124.9
R7924 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t24 124.9
R7925 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t17 124.9
R7926 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t18 124.9
R7927 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t4 108.754
R7928 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n25 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t2 108.365
R7929 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t11 20.8855
R7930 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 9.08711
R7931 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n25 7.91883
R7932 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n27 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n26 5.02291
R7933 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n21 3.41379
R7934 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n28 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n27 3.40258
R7935 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n19 1.27824
R7936 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n17 1.27824
R7937 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n15 1.27824
R7938 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n13 1.27824
R7939 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n11 1.27824
R7940 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n9 1.27824
R7941 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n7 1.27824
R7942 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n5 1.27824
R7943 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n3 1.27824
R7944 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n1 1.27824
R7945 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R7946 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n18 0.391454
R7947 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R7948 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n16 0.391454
R7949 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R7950 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n14 0.391454
R7951 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R7952 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n12 0.391454
R7953 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R7954 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n10 0.391454
R7955 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R7956 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n8 0.391454
R7957 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R7958 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n6 0.391454
R7959 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R7960 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n4 0.391454
R7961 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R7962 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n2 0.391454
R7963 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R7964 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n0 0.391454
R7965 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n25 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n24 0.310917
R7966 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n22 0.270394
R7967 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n20 0.266454
R7968 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n23 0.224458
R7969 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n28 0.063
R7970 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.0498421
R7971 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t1 227.856
R7972 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R7973 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t3 140.163
R7974 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t2 114.031
R7975 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t0 83.3993
R7976 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t4 81.5883
R7977 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R7978 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R7979 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R7980 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R7981 a_44234_9966.t0 a_44234_9966.t1 114.052
R7982 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t11 241.862
R7983 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t10 222.089
R7984 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t20 221.974
R7985 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t14 221.974
R7986 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t6 221.913
R7987 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t4 221.913
R7988 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t19 221.913
R7989 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t0 221.913
R7990 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t18 221.911
R7991 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t8 221.911
R7992 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t3 221.851
R7993 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t7 221.851
R7994 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t21 221.851
R7995 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t13 221.851
R7996 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t12 221.851
R7997 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t16 221.851
R7998 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t5 221.851
R7999 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t17 221.851
R8000 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t1 221.851
R8001 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t9 221.851
R8002 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t2 221.851
R8003 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t15 221.851
R8004 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t77 111.398
R8005 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n84 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t61 111.398
R8006 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t53 111.398
R8007 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t28 111.398
R8008 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t76 110.615
R8009 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t56 110.615
R8010 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t35 110.615
R8011 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n47 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t81 110.615
R8012 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t59 110.615
R8013 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t37 110.615
R8014 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t36 110.615
R8015 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t74 110.615
R8016 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t48 110.615
R8017 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t42 110.615
R8018 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t66 110.615
R8019 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t64 110.615
R8020 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t44 110.615
R8021 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t24 110.615
R8022 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t23 110.615
R8023 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n84 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t60 110.615
R8024 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n85 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t38 110.615
R8025 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n86 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t78 110.615
R8026 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n87 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t62 110.615
R8027 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n88 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t41 110.615
R8028 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n89 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t22 110.615
R8029 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n90 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t80 110.615
R8030 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n91 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t58 110.615
R8031 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n83 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t32 110.615
R8032 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n82 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t27 110.615
R8033 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n81 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t49 110.615
R8034 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n80 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t47 110.615
R8035 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n79 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t29 110.615
R8036 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t67 110.615
R8037 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n77 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t65 110.615
R8038 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t33 110.615
R8039 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t69 110.615
R8040 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t54 110.615
R8041 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t34 110.615
R8042 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t72 110.615
R8043 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t70 110.615
R8044 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t51 110.615
R8045 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t26 110.615
R8046 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t75 110.615
R8047 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t40 110.615
R8048 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t39 110.615
R8049 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n74 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t79 110.615
R8050 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n75 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t57 110.615
R8051 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t63 110.615
R8052 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t43 110.615
R8053 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t30 110.615
R8054 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t68 110.615
R8055 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t46 110.615
R8056 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t45 110.615
R8057 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t25 110.615
R8058 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n55 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t55 110.615
R8059 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n56 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t50 110.615
R8060 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t73 110.615
R8061 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n58 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t71 110.615
R8062 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t52 110.615
R8063 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t31 110.615
R8064 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 8.31322
R8065 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n15 5.697
R8066 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n20 5.697
R8067 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n3 5.697
R8068 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n0 5.6845
R8069 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n4 5.55802
R8070 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n6 5.55802
R8071 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n8 5.55802
R8072 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n10 5.55802
R8073 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n23 5.55802
R8074 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n21 5.55802
R8075 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n16 5.55802
R8076 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n18 5.55802
R8077 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n12 5.43008
R8078 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n75 5.35189
R8079 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n61 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n60 5.35189
R8080 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n77 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n76 4.88189
R8081 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n29 4.56856
R8082 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n52 3.72383
R8083 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n53 3.4105
R8084 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n27 3.4105
R8085 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n93 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n92 3.4105
R8086 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n25 3.4105
R8087 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n7 2.888
R8088 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n24 1.57967
R8089 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n19 1.30883
R8090 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n28 1.30883
R8091 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n1 1.07342
R8092 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n13 1.07342
R8093 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n77 0.783833
R8094 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n79 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n78 0.783833
R8095 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n80 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n79 0.783833
R8096 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n81 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n80 0.783833
R8097 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n82 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n81 0.783833
R8098 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n83 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n82 0.783833
R8099 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n91 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n90 0.783833
R8100 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n90 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n89 0.783833
R8101 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n89 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n88 0.783833
R8102 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n88 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n87 0.783833
R8103 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n87 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n86 0.783833
R8104 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n86 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n85 0.783833
R8105 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n85 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n84 0.783833
R8106 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n75 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n74 0.783833
R8107 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n74 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n73 0.783833
R8108 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n72 0.783833
R8109 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n71 0.783833
R8110 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n70 0.783833
R8111 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n67 0.783833
R8112 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n66 0.783833
R8113 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n65 0.783833
R8114 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n64 0.783833
R8115 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n63 0.783833
R8116 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n62 0.783833
R8117 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n59 0.783833
R8118 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n58 0.783833
R8119 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n58 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n57 0.783833
R8120 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n56 0.783833
R8121 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n56 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n55 0.783833
R8122 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n35 0.783833
R8123 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n34 0.783833
R8124 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n33 0.783833
R8125 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n32 0.783833
R8126 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n31 0.783833
R8127 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n30 0.783833
R8128 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n37 0.783833
R8129 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n38 0.783833
R8130 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n39 0.783833
R8131 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n40 0.783833
R8132 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n41 0.783833
R8133 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n42 0.783833
R8134 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n50 0.783833
R8135 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n49 0.783833
R8136 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n48 0.783833
R8137 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n47 0.783833
R8138 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n47 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n46 0.783833
R8139 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n45 0.783833
R8140 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n44 0.783833
R8141 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n92 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n91 0.527583
R8142 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n68 0.527583
R8143 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n36 0.527583
R8144 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n51 0.527583
R8145 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n61 0.390742
R8146 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n27 0.390742
R8147 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n61 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n29 0.313833
R8148 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n93 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n27 0.313833
R8149 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n92 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n83 0.25675
R8150 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n69 0.25675
R8151 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n55 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n54 0.25675
R8152 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n43 0.25675
R8153 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n16 0.246333
R8154 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n21 0.246333
R8155 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n8 0.246333
R8156 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n4 0.246333
R8157 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n93 0.174258
R8158 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n5 0.123417
R8159 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n9 0.123417
R8160 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n22 0.123417
R8161 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n17 0.123417
R8162 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n26 0.0916515
R8163 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n2 0.0604849
R8164 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n14 0.0604849
R8165 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n11 0.013
R8166 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t4 228.174
R8167 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t30 228.174
R8168 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t2 228.174
R8169 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t3 228.174
R8170 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t1 226.853
R8171 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t5 226.853
R8172 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t27 226.853
R8173 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t7 226.853
R8174 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t24 226.853
R8175 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t28 226.853
R8176 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t26 226.853
R8177 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t6 226.853
R8178 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t25 226.853
R8179 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t29 226.853
R8180 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t31 226.853
R8181 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t0 226.853
R8182 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t21 221.911
R8183 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t10 221.911
R8184 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t23 221.911
R8185 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t9 221.911
R8186 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t22 221.911
R8187 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t18 221.911
R8188 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t14 221.911
R8189 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t15 221.911
R8190 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t11 221.911
R8191 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t12 221.911
R8192 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t8 221.911
R8193 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t17 221.911
R8194 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t13 221.911
R8195 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t19 221.911
R8196 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t16 221.911
R8197 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t20 221.911
R8198 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n22 7.63383
R8199 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n15 7.63383
R8200 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n18 7.63383
R8201 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n27 7.49842
R8202 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n6 5.05408
R8203 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n23 4.5005
R8204 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n25 4.5005
R8205 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n16 4.5005
R8206 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n19 4.5005
R8207 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n21 4.30208
R8208 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n28 3.4105
R8209 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n13 3.4105
R8210 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n24 3.13383
R8211 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n0 1.813
R8212 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n2 1.813
R8213 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n4 1.813
R8214 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n7 1.813
R8215 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n10 1.813
R8216 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n17 1.70258
R8217 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n20 1.43175
R8218 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n1 1.32133
R8219 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n8 1.32133
R8220 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n11 1.32133
R8221 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n9 1.04217
R8222 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n3 0.796333
R8223 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n12 0.771333
R8224 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n5 0.5255
R8225 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n14 0.279652
R8226 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n29 0.236924
R8227 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n26 0.135917
R8228 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t4 739.082
R8229 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t15 241.536
R8230 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t9 230.155
R8231 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t17 230.155
R8232 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t18 230.155
R8233 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t12 230.155
R8234 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t10 230.155
R8235 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t8 230.155
R8236 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n26 203.922
R8237 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 181.496
R8238 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t5 169.237
R8239 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t16 157.856
R8240 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t11 157.856
R8241 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t6 157.856
R8242 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t13 157.856
R8243 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t7 157.856
R8244 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t14 157.856
R8245 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 154.867
R8246 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 153.911
R8247 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 153.338
R8248 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 152
R8249 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 152
R8250 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 152
R8251 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 101.49
R8252 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t2 26.5955
R8253 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t0 26.5955
R8254 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 25.9222
R8255 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t3 24.9236
R8256 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t1 24.9236
R8257 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 21.542
R8258 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 21.248
R8259 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 19.5688
R8260 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 19.3054
R8261 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 18.6011
R8262 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 18.542
R8263 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y 13.0565
R8264 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[0] 12.2693
R8265 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 12.2559
R8266 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 11.1817
R8267 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 11.0199
R8268 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y 10.7525
R8269 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y 6.6565
R8270 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 5.10675
R8271 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 5.04292
R8272 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 4.3525
R8273 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x2.A 3.05722
R8274 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x1.B 2.5605
R8275 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 2.5605
R8276 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.A 2.48408
R8277 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.A 2.10199
R8278 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.A 2.10199
R8279 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x2.A 2.10199
R8280 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y 1.93989
R8281 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x3.A 1.52886
R8282 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 1.40284
R8283 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 1.23683
R8284 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 0.926281
R8285 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 0.842297
R8286 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[6] 0.119641
R8287 a_44234_17252.t0 a_44234_17252.t1 114.052
R8288 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t21 154.608
R8289 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t43 142.488
R8290 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t25 142.488
R8291 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t49 142.488
R8292 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t36 142.488
R8293 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t72 142.488
R8294 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n47 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t53 142.488
R8295 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n74 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t77 142.488
R8296 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t62 142.488
R8297 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t64 141.704
R8298 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t24 141.704
R8299 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t101 141.704
R8300 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t65 141.704
R8301 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t87 141.704
R8302 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t98 141.704
R8303 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t42 141.704
R8304 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t70 141.704
R8305 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t99 141.704
R8306 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t50 141.704
R8307 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t46 141.704
R8308 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t82 141.704
R8309 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t30 141.704
R8310 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t81 141.704
R8311 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t80 141.704
R8312 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t22 141.704
R8313 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t66 141.704
R8314 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t89 141.704
R8315 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t67 141.704
R8316 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t34 141.704
R8317 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t29 141.704
R8318 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t69 141.704
R8319 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t94 141.704
R8320 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t26 141.704
R8321 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t44 141.704
R8322 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t75 141.704
R8323 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t28 141.704
R8324 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t59 141.704
R8325 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t54 141.704
R8326 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t90 141.704
R8327 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t39 141.704
R8328 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t88 141.704
R8329 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t85 141.704
R8330 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t33 141.704
R8331 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t71 141.704
R8332 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t96 141.704
R8333 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t83 141.704
R8334 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n55 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t52 141.704
R8335 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n56 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t48 141.704
R8336 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t84 141.704
R8337 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n58 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t32 141.704
R8338 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t45 141.704
R8339 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t68 141.704
R8340 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n61 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t93 141.704
R8341 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t47 141.704
R8342 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t76 141.704
R8343 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t74 141.704
R8344 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t27 141.704
R8345 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t57 141.704
R8346 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t23 141.704
R8347 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t100 141.704
R8348 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t51 141.704
R8349 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t86 141.704
R8350 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n47 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t37 141.704
R8351 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n74 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t91 141.704
R8352 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n75 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t61 141.704
R8353 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t58 141.704
R8354 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n77 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t92 141.704
R8355 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t40 141.704
R8356 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n79 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t55 141.704
R8357 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n80 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t73 141.704
R8358 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n81 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t97 141.704
R8359 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n82 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t56 141.704
R8360 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n83 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t79 141.704
R8361 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n84 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t78 141.704
R8362 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t38 141.704
R8363 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t63 141.704
R8364 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t35 141.704
R8365 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t31 141.704
R8366 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t60 141.704
R8367 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t95 141.704
R8368 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t41 141.704
R8369 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t17 134.811
R8370 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n87 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t4 134.712
R8371 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n89 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t16 134.712
R8372 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n89 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t13 134.712
R8373 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n90 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t14 134.712
R8374 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n90 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t1 134.712
R8375 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n92 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t8 134.712
R8376 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n92 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t2 134.712
R8377 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t3 134.712
R8378 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t15 134.712
R8379 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t10 134.712
R8380 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t18 134.712
R8381 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t9 134.712
R8382 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t5 134.712
R8383 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t20 134.712
R8384 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t19 134.712
R8385 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n97 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t7 134.712
R8386 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n97 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t6 134.712
R8387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n99 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t12 134.712
R8388 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n99 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t11 134.712
R8389 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n87 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t0 134.712
R8390 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n102 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n101 9.92246
R8391 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n101 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n2 9.18808
R8392 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n91 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n89 7.7474
R8393 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n3 7.7474
R8394 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n101 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n100 5.72717
R8395 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n95 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n94 5.30474
R8396 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n91 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n90 4.61407
R8397 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n93 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n92 4.61407
R8398 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n1 4.61407
R8399 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n4 4.61407
R8400 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n6 4.61407
R8401 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n98 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n97 4.61407
R8402 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n100 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n99 4.61407
R8403 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n88 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n87 4.61407
R8404 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n26 4.07135
R8405 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n86 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n85 3.4105
R8406 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n65 3.4105
R8407 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n45 3.4105
R8408 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n96 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n95 3.4105
R8409 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n100 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n98 3.13383
R8410 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n5 3.13383
R8411 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n88 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n2 3.13383
R8412 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n93 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n91 3.13383
R8413 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n98 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n96 2.73592
R8414 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n94 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n93 1.96508
R8415 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n102 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n0 1.87758
R8416 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n94 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n88 1.16925
R8417 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n8 0.783833
R8418 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n9 0.783833
R8419 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n10 0.783833
R8420 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n11 0.783833
R8421 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n12 0.783833
R8422 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n13 0.783833
R8423 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n24 0.783833
R8424 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n23 0.783833
R8425 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n22 0.783833
R8426 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n21 0.783833
R8427 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n20 0.783833
R8428 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n19 0.783833
R8429 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n18 0.783833
R8430 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n17 0.783833
R8431 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n16 0.783833
R8432 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n15 0.783833
R8433 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n27 0.783833
R8434 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n28 0.783833
R8435 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n29 0.783833
R8436 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n30 0.783833
R8437 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n31 0.783833
R8438 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n32 0.783833
R8439 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n43 0.783833
R8440 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n42 0.783833
R8441 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n41 0.783833
R8442 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n40 0.783833
R8443 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n39 0.783833
R8444 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n38 0.783833
R8445 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n37 0.783833
R8446 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n36 0.783833
R8447 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n35 0.783833
R8448 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n34 0.783833
R8449 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n47 0.783833
R8450 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n48 0.783833
R8451 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n49 0.783833
R8452 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n50 0.783833
R8453 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n51 0.783833
R8454 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n52 0.783833
R8455 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n63 0.783833
R8456 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n62 0.783833
R8457 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n61 0.783833
R8458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n61 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n60 0.783833
R8459 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n59 0.783833
R8460 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n58 0.783833
R8461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n58 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n57 0.783833
R8462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n56 0.783833
R8463 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n56 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n55 0.783833
R8464 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n55 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n54 0.783833
R8465 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n67 0.783833
R8466 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n68 0.783833
R8467 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n69 0.783833
R8468 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n70 0.783833
R8469 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n71 0.783833
R8470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n72 0.783833
R8471 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n84 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n83 0.783833
R8472 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n83 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n82 0.783833
R8473 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n82 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n81 0.783833
R8474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n81 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n80 0.783833
R8475 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n80 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n79 0.783833
R8476 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n79 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n78 0.783833
R8477 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n77 0.783833
R8478 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n77 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n76 0.783833
R8479 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n75 0.783833
R8480 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n75 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n74 0.783833
R8481 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n14 0.777583
R8482 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n33 0.777583
R8483 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n53 0.777583
R8484 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n85 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n73 0.777583
R8485 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n86 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n66 0.661348
R8486 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n96 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n7 0.398417
R8487 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n95 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n86 0.328076
R8488 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n46 0.140076
R8489 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n102 0.0755
R8490 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n25 0.00675
R8491 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n44 0.00675
R8492 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n64 0.00675
R8493 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n85 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n84 0.00675
R8494 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t35 141.215
R8495 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t28 141.215
R8496 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t24 141.215
R8497 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t25 141.215
R8498 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t26 139.879
R8499 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t27 139.879
R8500 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t33 139.879
R8501 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t38 139.879
R8502 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t36 139.879
R8503 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t30 139.879
R8504 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t31 139.879
R8505 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t37 139.879
R8506 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t23 139.879
R8507 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t22 139.879
R8508 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t39 139.879
R8509 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t29 139.879
R8510 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t34 139.879
R8511 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t20 139.879
R8512 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t32 139.879
R8513 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t21 139.879
R8514 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t7 134.738
R8515 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t14 134.738
R8516 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t9 134.738
R8517 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t8 134.738
R8518 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t1 134.738
R8519 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t6 134.738
R8520 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t0 134.738
R8521 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t2 134.738
R8522 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t18 134.738
R8523 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t11 134.738
R8524 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t12 134.738
R8525 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t13 134.738
R8526 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t5 134.738
R8527 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t3 134.738
R8528 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t4 134.738
R8529 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t16 134.738
R8530 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t17 134.738
R8531 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t15 134.738
R8532 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t10 134.738
R8533 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n37 134.738
R8534 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n24 7.63383
R8535 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n29 7.63383
R8536 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n36 7.63383
R8537 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n0 7.63383
R8538 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n13 5.55541
R8539 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n33 4.52426
R8540 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n25 4.5005
R8541 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n27 4.5005
R8542 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n30 4.5005
R8543 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n35 4.5005
R8544 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n3 4.5005
R8545 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n1 4.5005
R8546 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n22 3.4105
R8547 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n32 3.4105
R8548 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n26 3.13383
R8549 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n2 3.13383
R8550 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n31 3.00675
R8551 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n14 1.79633
R8552 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n19 1.79633
R8553 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n17 1.79633
R8554 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n5 1.79633
R8555 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n7 1.79633
R8556 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n11 1.79633
R8557 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n9 1.79633
R8558 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n34 1.69425
R8559 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n4 1.44008
R8560 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n15 1.338
R8561 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n20 1.338
R8562 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n18 1.338
R8563 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n6 1.338
R8564 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n10 1.338
R8565 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n16 1.0255
R8566 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n8 0.796333
R8567 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n21 0.771333
R8568 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n12 0.542167
R8569 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n23 0.3765
R8570 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n28 0.127583
R8571 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t8 752.088
R8572 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t7 212.081
R8573 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t6 212.081
R8574 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 203.922
R8575 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 186.001
R8576 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t5 139.78
R8577 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t4 139.78
R8578 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 101.49
R8579 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 61.346
R8580 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t0 26.5955
R8581 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t1 26.5955
R8582 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t2 24.9236
R8583 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t3 24.9236
R8584 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y 13.5685
R8585 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y 10.7525
R8586 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 9.64425
R8587 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 9.30224
R8588 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y 6.6565
R8589 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 5.04292
R8590 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 3.8405
R8591 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.A 3.0725
R8592 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 2.5605
R8593 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y 1.93989
R8594 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t4 761.467
R8595 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 203.923
R8596 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 101.49
R8597 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t3 26.5955
R8598 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t2 26.5955
R8599 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t1 24.9236
R8600 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t0 24.9236
R8601 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 13.0565
R8602 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 10.7525
R8603 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y 6.6565
R8604 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y 5.04292
R8605 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y 4.3525
R8606 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y 2.5605
R8607 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 1.93989
R8608 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t0 274.793
R8609 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t6 230.576
R8610 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t5 230.155
R8611 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t7 229.369
R8612 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n9 205.28
R8613 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t8 158.275
R8614 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n0 157.927
R8615 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t9 157.856
R8616 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t4 157.07
R8617 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n5 153.067
R8618 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n1 152
R8619 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t2 133.124
R8620 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n10 67.4857
R8621 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n8 36.3299
R8622 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t1 26.5955
R8623 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t3 26.5955
R8624 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n4 24.8988
R8625 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n3 13.8092
R8626 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n2 12.5635
R8627 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n7 10.6878
R8628 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n6 9.3005
R8629 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 7.11161
R8630 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 5.67507
R8631 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 5.6005
R8632 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 2.13383
R8633 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.602583
R8634 a_45023_21964.t0 a_45023_21964.t1 49.8467
R8635 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t14 141.399
R8636 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t13 141.399
R8637 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t8 141.399
R8638 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t11 141.399
R8639 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t9 140.061
R8640 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t15 140.061
R8641 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t10 140.061
R8642 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t12 140.061
R8643 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t3 134.732
R8644 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t1 134.732
R8645 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t5 134.732
R8646 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t2 134.732
R8647 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t4 134.712
R8648 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t0 134.712
R8649 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t6 134.712
R8650 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n13 134.712
R8651 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n12 8.29542
R8652 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n2 6.98292
R8653 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n1 6.72342
R8654 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n0 5.41092
R8655 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n3 3.89759
R8656 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n6 3.55008
R8657 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n9 3.4105
R8658 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n11 3.4105
R8659 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n4 3.12133
R8660 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n8 1.80883
R8661 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n10 1.6925
R8662 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n7 1.55467
R8663 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n5 0.242167
R8664 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t13 241.536
R8665 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t10 241.536
R8666 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t9 230.155
R8667 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t18 230.155
R8668 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t15 229.369
R8669 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t5 228.649
R8670 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t11 212.081
R8671 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t8 212.081
R8672 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n0 203.923
R8673 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n3 186.001
R8674 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t17 169.237
R8675 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t6 169.237
R8676 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n5 157.927
R8677 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t19 157.856
R8678 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t4 157.856
R8679 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t7 157.07
R8680 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t12 156.35
R8681 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n11 154.934
R8682 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n13 154.744
R8683 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n15 154.744
R8684 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n8 153.338
R8685 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n6 152
R8686 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t16 139.78
R8687 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t14 139.78
R8688 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n20 101.49
R8689 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n2 61.346
R8690 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t2 26.5955
R8691 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t3 26.5955
R8692 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t0 24.9236
R8693 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t1 24.9236
R8694 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 24.013
R8695 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 21.1432
R8696 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 19.8144
R8697 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n7 19.6746
R8698 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n16 18.2347
R8699 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n9 18.2231
R8700 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 17.3957
R8701 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n19 13.5685
R8702 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n17 12.788
R8703 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n1 10.7525
R8704 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n18 9.64425
R8705 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n4 9.30224
R8706 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 6.6565
R8707 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 5.04292
R8708 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 3.8405
R8709 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 3.0725
R8710 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 3.05722
R8711 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 2.5605
R8712 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n14 2.37941
R8713 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 2.13383
R8714 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n21 1.93989
R8715 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n12 1.08448
R8716 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n10 1.05323
R8717 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.186047
R8718 a_43167_4358.t0 a_43167_4358.t1 49.8467
R8719 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 272.038
R8720 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t0 258.846
R8721 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t4 228.463
R8722 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n0 224.776
R8723 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t3 157.07
R8724 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n1 152
R8725 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n2 30.3559
R8726 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t1 26.5955
R8727 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t2 26.5955
R8728 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 4.20621
R8729 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n4 3.03935
R8730 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 2.30266
R8731 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n3 2.25932
R8732 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 1.50638
R8733 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n5 0.921363
R8734 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t30 141.399
R8735 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t31 141.399
R8736 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t36 141.399
R8737 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t35 141.399
R8738 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t37 140.061
R8739 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t29 140.061
R8740 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t25 140.061
R8741 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t39 140.061
R8742 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t38 140.061
R8743 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t27 140.061
R8744 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t26 140.061
R8745 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t32 140.061
R8746 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t33 140.061
R8747 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t34 140.061
R8748 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t21 140.061
R8749 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t28 140.061
R8750 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t22 140.061
R8751 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t20 140.061
R8752 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t24 140.061
R8753 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t23 140.061
R8754 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t0 134.738
R8755 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t1 134.738
R8756 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t15 134.738
R8757 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t13 134.738
R8758 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t14 134.738
R8759 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t7 134.738
R8760 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t8 134.738
R8761 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t6 134.738
R8762 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t18 134.738
R8763 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t9 134.738
R8764 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t5 134.738
R8765 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t4 134.738
R8766 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t16 134.738
R8767 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t2 134.738
R8768 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t12 134.738
R8769 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t17 134.738
R8770 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t10 134.738
R8771 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t11 134.738
R8772 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t3 134.738
R8773 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n37 134.738
R8774 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n24 7.63383
R8775 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n27 7.63383
R8776 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n0 7.63383
R8777 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n36 7.63383
R8778 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n13 5.68074
R8779 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n33 4.64959
R8780 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n25 4.5005
R8781 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n30 4.5005
R8782 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n28 4.5005
R8783 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n1 4.5005
R8784 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n3 4.5005
R8785 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n35 4.5005
R8786 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n22 3.4105
R8787 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n32 3.4105
R8788 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n29 3.13383
R8789 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n2 3.13383
R8790 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n34 2.74425
R8791 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n26 1.95675
R8792 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n14 1.79633
R8793 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n16 1.79633
R8794 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n20 1.79633
R8795 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n18 1.79633
R8796 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n5 1.79633
R8797 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n10 1.79633
R8798 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n8 1.79633
R8799 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n15 1.338
R8800 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n19 1.338
R8801 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n6 1.338
R8802 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n11 1.338
R8803 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n9 1.338
R8804 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n7 1.288
R8805 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n31 1.17758
R8806 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n17 1.05883
R8807 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n12 0.508833
R8808 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n4 0.390083
R8809 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n21 0.279667
R8810 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n23 0.251167
R8811 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t15 738.899
R8812 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t11 241.536
R8813 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t14 232.214
R8814 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t10 232.214
R8815 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t13 229.369
R8816 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t16 229.369
R8817 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t19 229.369
R8818 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t20 212.081
R8819 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t12 212.081
R8820 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 203.923
R8821 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 186.001
R8822 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t17 169.237
R8823 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t18 159.915
R8824 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t7 159.915
R8825 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t6 157.07
R8826 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t8 157.07
R8827 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t5 157.07
R8828 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 155.88
R8829 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 154.065
R8830 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 152.712
R8831 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 152.475
R8832 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 152
R8833 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 152
R8834 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t9 139.78
R8835 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t4 139.78
R8836 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 101.49
R8837 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 61.346
R8838 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t2 26.5955
R8839 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t3 26.5955
R8840 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t0 24.9236
R8841 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t1 24.9236
R8842 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 23.417
R8843 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 21.961
R8844 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 20.0025
R8845 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 18.2158
R8846 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 15.6884
R8847 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 13.5685
R8848 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 12.4213
R8849 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[0] 11.8734
R8850 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 10.9817
R8851 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 10.7525
R8852 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 10.2234
R8853 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 9.77342
R8854 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 9.64425
R8855 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 9.30224
R8856 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x2.C 6.98232
R8857 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y 6.6565
R8858 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x1.B 5.92643
R8859 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.B 5.45235
R8860 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.B 5.21532
R8861 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y 5.04292
R8862 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 4.91925
R8863 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y 3.8405
R8864 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.A 3.0725
R8865 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.A 2.68437
R8866 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y 2.5605
R8867 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 2.30909
R8868 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 1.93989
R8869 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 1.42823
R8870 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.A 0.970197
R8871 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 0.623547
R8872 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[6] 0.451672
R8873 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t2 674.658
R8874 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t0 10.7661
R8875 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t1 10.7361
R8876 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.n0 4.09773
R8877 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t0 673.34
R8878 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t2 10.7207
R8879 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t1 10.6931
R8880 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.n0 3.42321
R8881 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t8 754.659
R8882 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t5 212.081
R8883 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t4 212.081
R8884 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 203.922
R8885 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 186.001
R8886 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t7 139.78
R8887 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t6 139.78
R8888 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 101.49
R8889 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 61.346
R8890 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t3 26.5955
R8891 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t0 26.5955
R8892 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t1 24.9236
R8893 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t2 24.9236
R8894 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y 13.5685
R8895 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y 10.7525
R8896 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 9.64425
R8897 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 9.30224
R8898 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y 6.6565
R8899 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 5.04292
R8900 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 3.8405
R8901 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.A 3.0725
R8902 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 2.5605
R8903 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y 1.93989
R8904 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t4 762.88
R8905 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 203.923
R8906 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 101.49
R8907 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t3 26.5955
R8908 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t2 26.5955
R8909 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t1 24.9236
R8910 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t0 24.9236
R8911 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 13.0565
R8912 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 10.7525
R8913 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y 6.6565
R8914 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y 5.04292
R8915 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y 4.3525
R8916 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y 2.5605
R8917 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 1.93989
R8918 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n1 863.124
R8919 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n0 585
R8920 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t0 495.469
R8921 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t4 223.218
R8922 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t5 217.042
R8923 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t2 216.63
R8924 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t3 208.054
R8925 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t1 141.189
R8926 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t0 140.738
R8927 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n5 30.8338
R8928 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.b[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n7 29.688
R8929 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUT 14.3755
R8930 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 11.6369
R8931 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n6 10.8443
R8932 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 10.1408
R8933 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n8 8.53383
R8934 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n3 7.94225
R8935 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n5 top_DAC_0/top_final_switch_0.b[0] 7.89425
R8936 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 6.14988
R8937 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 5.81868
R8938 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.b[0] 4.71204
R8939 top_DAC_0/top_final_switch_0.b[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n4 3.59409
R8940 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 2.16154
R8941 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n2 0.665435
R8942 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUT top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.b[0] 0.19425
R8943 top_DAC_0/top_rseg_n_dcell_0.VH2.n0 top_DAC_0/top_rseg_n_dcell_0.VH2.t4 244.607
R8944 top_DAC_0/top_rseg_n_dcell_0.VH2.n1 top_DAC_0/top_rseg_n_dcell_0.VH2.t6 239.264
R8945 top_DAC_0/top_rseg_n_dcell_0.VH2.n3 top_DAC_0/top_rseg_n_dcell_0.VH2.t7 234.764
R8946 top_DAC_0/top_rseg_n_dcell_0.VH2.n0 top_DAC_0/top_rseg_n_dcell_0.VH2.t3 234.399
R8947 top_DAC_0/top_rseg_n_dcell_0.VH2.n4 top_DAC_0/top_rseg_n_dcell_0.VH2.t2 234.293
R8948 top_DAC_0/top_rseg_n_dcell_0.VH2.n6 top_DAC_0/top_rseg_n_dcell_0.VH2.t1 233.657
R8949 top_DAC_0/top_rseg_n_dcell_0.VH2.n4 top_DAC_0/top_rseg_n_dcell_0.VH2.t5 233.657
R8950 top_DAC_0/top_rseg_n_dcell_0.VH2.n5 top_DAC_0/top_rseg_n_dcell_0.VH2.t0 233.657
R8951 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.VH2.n3 30.4838
R8952 top_DAC_0/top_rseg_n_dcell_0.VH2.n1 top_DAC_0/top_rseg_n_dcell_0.VH2.n0 6.0755
R8953 top_DAC_0/top_rseg_n_dcell_0.VH2.n3 top_DAC_0/top_rseg_n_dcell_0.VH2.n2 4.5005
R8954 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.VH2.n1 1.09842
R8955 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.VH2.n6 1.00675
R8956 top_DAC_0/top_rseg_n_dcell_0.VH2.n6 top_DAC_0/top_rseg_n_dcell_0.VH2.n5 0.63637
R8957 top_DAC_0/top_rseg_n_dcell_0.VH2.n5 top_DAC_0/top_rseg_n_dcell_0.VH2.n4 0.63637
R8958 top_DAC_0/top_rseg_n_dcell_0.VH2.n2 top_DAC_0/top_rseg_n_dcell_0.VH2 0.110917
R8959 top_DAC_0/top_rseg_n_dcell_0.VH2.n2 top_DAC_0/top_rseg_n_dcell_0.VH2 0.063
R8960 a_14615_13536.t0 a_14615_13536.n0 439.543
R8961 a_14615_13536.n0 a_14615_13536.t2 39.3576
R8962 a_14615_13536.n0 a_14615_13536.t1 39.3576
R8963 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n1 863.124
R8964 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n0 585
R8965 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t0 495.469
R8966 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t10 217.555
R8967 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t8 216.893
R8968 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t6 216.893
R8969 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t13 216.893
R8970 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t3 215.142
R8971 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t11 213.218
R8972 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t12 213.218
R8973 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t7 212.554
R8974 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t2 212.393
R8975 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t5 208.054
R8976 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n14 152
R8977 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t1 141.189
R8978 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t0 140.738
R8979 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t9 114.031
R8980 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t4 81.5883
R8981 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n9 29.0755
R8982 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n13 22.0693
R8983 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 16.7132
R8984 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 14.6338
R8985 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 13.7979
R8986 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 13.1884
R8987 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 11.6369
R8988 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n12 11.3942
R8989 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n8 11.3755
R8990 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 10.1408
R8991 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n3 7.94225
R8992 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 6.14988
R8993 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n7 4.5005
R8994 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n11 4.5005
R8995 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n4 4.23159
R8996 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 2.16154
R8997 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 2.16154
R8998 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n15 1.16414
R8999 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n2 0.665435
R9000 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n5 0.663962
R9001 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n6 0.663962
R9002 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n16 0.582318
R9003 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n10 0.445212
R9004 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.28175
R9005 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.21925
R9006 a_19946_8950.t0 a_19946_8950.n0 671.561
R9007 a_19946_8950.n0 a_19946_8950.t2 671.109
R9008 a_19946_8950.n0 a_19946_8950.t1 665.524
R9009 a_20656_10031.n0 a_20656_10031.t1 667.841
R9010 a_20656_10031.n0 a_20656_10031.t2 667.491
R9011 a_20656_10031.t0 a_20656_10031.n0 665.484
R9012 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t0 227.856
R9013 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R9014 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t2 140.163
R9015 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t4 114.031
R9016 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t1 83.3993
R9017 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t3 81.5883
R9018 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R9019 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R9020 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R9021 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R9022 a_43724_9372.t0 a_43724_9372.t1 55.3905
R9023 a_43698_8776.t0 a_43698_8776.n0 228.04
R9024 a_43698_8776.n0 a_43698_8776.t2 145.648
R9025 a_43698_8776.n0 a_43698_8776.t1 83.2159
R9026 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t1 334.771
R9027 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t2 213.218
R9028 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t6 212.989
R9029 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t4 212.554
R9030 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t3 212.554
R9031 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t7 208.054
R9032 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t5 131.306
R9033 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t8 126.278
R9034 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t9 125.566
R9035 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t0 87.8231
R9036 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n3 56.8068
R9037 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n7 5.12863
R9038 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n5 4.68383
R9039 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n2 4.5005
R9040 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n0 0.663962
R9041 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n1 0.663962
R9042 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n4 0.608192
R9043 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.228865
R9044 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n6 0.177583
R9045 a_22193_18133.n0 a_22193_18133.t4 244.489
R9046 a_22193_18133.n2 a_22193_18133.t1 242.548
R9047 a_22193_18133.n0 a_22193_18133.t2 239.614
R9048 a_22193_18133.n1 a_22193_18133.t3 239.614
R9049 a_22193_18133.t0 a_22193_18133.n2 239.614
R9050 a_22193_18133.n2 a_22193_18133.n1 2.93383
R9051 a_22193_18133.n1 a_22193_18133.n0 2.93383
R9052 a_23307_20174.n1 a_23307_20174.t3 249.702
R9053 a_23307_20174.n0 a_23307_20174.t2 248.171
R9054 a_23307_20174.n0 a_23307_20174.t1 240.933
R9055 a_23307_20174.t0 a_23307_20174.n2 240.933
R9056 a_23307_20174.n1 a_23307_20174.t4 239.614
R9057 a_23307_20174.n2 a_23307_20174.n1 0.898417
R9058 a_23307_20174.n2 a_23307_20174.n0 0.633833
R9059 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n1 863.124
R9060 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n0 585
R9061 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t0 495.469
R9062 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t5 217.555
R9063 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t2 216.893
R9064 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t4 216.893
R9065 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t3 216.893
R9066 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t7 212.393
R9067 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n9 152
R9068 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t1 141.189
R9069 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t0 140.738
R9070 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t6 114.031
R9071 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n8 93.4484
R9072 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t8 81.5883
R9073 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 16.7132
R9074 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 13.7979
R9075 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 13.1884
R9076 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 11.6369
R9077 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 10.1408
R9078 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n3 7.94225
R9079 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 6.14988
R9080 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n7 4.5005
R9081 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 2.16154
R9082 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 2.16154
R9083 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n10 1.16414
R9084 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n2 0.665435
R9085 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n4 0.663962
R9086 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n6 0.663962
R9087 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n5 0.663962
R9088 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n11 0.582318
R9089 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.202423
R9090 a_14790_18696.t0 a_14790_18696.n0 670.26
R9091 a_14790_18696.n0 a_14790_18696.t1 667.083
R9092 a_14790_18696.n0 a_14790_18696.t2 665.481
R9093 a_14948_18696.t0 a_14948_18696.n0 671.708
R9094 a_14948_18696.n0 a_14948_18696.t1 667.766
R9095 a_14948_18696.n0 a_14948_18696.t2 666.221
R9096 VOUT.n0 VOUT.t84 170.625
R9097 VOUT.n23 VOUT.t83 170.625
R9098 VOUT.n22 VOUT.t51 170.625
R9099 VOUT.n21 VOUT.t86 170.625
R9100 VOUT.n2 VOUT.t56 170.625
R9101 VOUT.n13 VOUT.t71 170.625
R9102 VOUT.n12 VOUT.t70 170.625
R9103 VOUT.n11 VOUT.t79 170.625
R9104 VOUT.n4 VOUT.t85 170.625
R9105 VOUT.n5 VOUT.t52 170.625
R9106 VOUT.n27 VOUT.t69 170.625
R9107 VOUT.n26 VOUT.t54 170.625
R9108 VOUT.n1 VOUT.t80 170.625
R9109 VOUT.n18 VOUT.t59 170.625
R9110 VOUT.n17 VOUT.t57 170.625
R9111 VOUT.n16 VOUT.t63 170.625
R9112 VOUT.n3 VOUT.t72 170.625
R9113 VOUT.n8 VOUT.t61 170.625
R9114 VOUT.n7 VOUT.t76 170.625
R9115 VOUT.n6 VOUT.t67 170.625
R9116 VOUT.n105 VOUT.t78 120.255
R9117 VOUT.n104 VOUT.t77 120.255
R9118 VOUT.n79 VOUT.t87 120.255
R9119 VOUT.n96 VOUT.t82 120.255
R9120 VOUT.n95 VOUT.t50 120.255
R9121 VOUT.n94 VOUT.t66 120.255
R9122 VOUT.n81 VOUT.t65 120.255
R9123 VOUT.n86 VOUT.t74 120.255
R9124 VOUT.n85 VOUT.t81 120.255
R9125 VOUT.n84 VOUT.t48 120.255
R9126 VOUT.n78 VOUT.t64 120.255
R9127 VOUT.n101 VOUT.t49 120.255
R9128 VOUT.n100 VOUT.t75 120.255
R9129 VOUT.n99 VOUT.t55 120.255
R9130 VOUT.n80 VOUT.t53 120.255
R9131 VOUT.n91 VOUT.t60 120.255
R9132 VOUT.n90 VOUT.t68 120.255
R9133 VOUT.n89 VOUT.t58 120.255
R9134 VOUT.n82 VOUT.t73 120.255
R9135 VOUT.n83 VOUT.t62 120.255
R9136 VOUT.n30 VOUT.n29 75.2042
R9137 VOUT.n30 VOUT.n28 75.1988
R9138 VOUT.n33 VOUT.n31 66.6872
R9139 VOUT.n33 VOUT.n32 66.6872
R9140 VOUT.n31 VOUT.t45 16.5305
R9141 VOUT.n31 VOUT.t44 16.5305
R9142 VOUT.n32 VOUT.t47 16.5305
R9143 VOUT.n32 VOUT.t46 16.5305
R9144 VOUT.n6 VOUT.n5 14.1588
R9145 VOUT.n84 VOUT.n83 12.4588
R9146 VOUT.n25 VOUT.n24 12.4088
R9147 VOUT.n20 VOUT.n19 12.4088
R9148 VOUT.n15 VOUT.n14 12.4088
R9149 VOUT.n10 VOUT.n9 12.4088
R9150 VOUT.n103 VOUT.n102 10.7088
R9151 VOUT.n98 VOUT.n97 10.7088
R9152 VOUT.n93 VOUT.n92 10.7088
R9153 VOUT.n88 VOUT.n87 10.7088
R9154 VOUT.n77 VOUT.n0 9.62342
R9155 VOUT.n28 VOUT.t38 9.23217
R9156 VOUT.n28 VOUT.t41 9.23217
R9157 VOUT.n29 VOUT.t40 9.23217
R9158 VOUT.n29 VOUT.t39 9.23217
R9159 VOUT.n73 VOUT.n72 9.02001
R9160 VOUT VOUT.n30 8.64633
R9161 VOUT.n106 VOUT.n78 7.38592
R9162 VOUT.n106 VOUT.n105 6.21508
R9163 VOUT.n76 VOUT.n75 6.10613
R9164 VOUT.n73 VOUT.n33 5.72967
R9165 VOUT.n77 VOUT.n76 4.5005
R9166 VOUT.n40 VOUT.n36 3.90596
R9167 VOUT.n72 VOUT.n71 3.4105
R9168 VOUT.n68 VOUT.n67 3.4105
R9169 VOUT.n64 VOUT.n63 3.4105
R9170 VOUT.n60 VOUT.n59 3.4105
R9171 VOUT.n56 VOUT.n55 3.4105
R9172 VOUT.n52 VOUT.n51 3.4105
R9173 VOUT.n48 VOUT.n47 3.4105
R9174 VOUT.n44 VOUT.n43 3.4105
R9175 VOUT.n40 VOUT.n39 3.4105
R9176 VOUT.n74 VOUT.n73 2.75779
R9177 VOUT.n87 VOUT.n85 1.91925
R9178 VOUT.n93 VOUT.n81 1.91925
R9179 VOUT.n97 VOUT.n95 1.91925
R9180 VOUT.n103 VOUT.n79 1.91925
R9181 VOUT.n10 VOUT.n4 1.91925
R9182 VOUT.n14 VOUT.n12 1.91925
R9183 VOUT.n20 VOUT.n2 1.91925
R9184 VOUT.n24 VOUT.n22 1.91925
R9185 VOUT.n83 VOUT.n82 1.613
R9186 VOUT.n90 VOUT.n89 1.613
R9187 VOUT.n91 VOUT.n80 1.613
R9188 VOUT.n100 VOUT.n99 1.613
R9189 VOUT.n101 VOUT.n78 1.613
R9190 VOUT.n7 VOUT.n6 1.613
R9191 VOUT.n8 VOUT.n3 1.613
R9192 VOUT.n17 VOUT.n16 1.613
R9193 VOUT.n18 VOUT.n1 1.613
R9194 VOUT.n27 VOUT.n26 1.613
R9195 VOUT.n88 VOUT.n82 1.38175
R9196 VOUT.n92 VOUT.n90 1.38175
R9197 VOUT.n98 VOUT.n80 1.38175
R9198 VOUT.n102 VOUT.n100 1.38175
R9199 VOUT.n9 VOUT.n7 1.38175
R9200 VOUT.n15 VOUT.n3 1.38175
R9201 VOUT.n19 VOUT.n17 1.38175
R9202 VOUT.n25 VOUT.n1 1.38175
R9203 VOUT.n76 VOUT.n27 1.17758
R9204 VOUT.n87 VOUT.n86 1.14425
R9205 VOUT.n94 VOUT.n93 1.14425
R9206 VOUT.n97 VOUT.n96 1.14425
R9207 VOUT.n104 VOUT.n103 1.14425
R9208 VOUT.n11 VOUT.n10 1.14425
R9209 VOUT.n14 VOUT.n13 1.14425
R9210 VOUT.n21 VOUT.n20 1.14425
R9211 VOUT.n24 VOUT.n23 1.14425
R9212 VOUT.n34 VOUT.t17 1.082
R9213 VOUT.n37 VOUT.t11 1.082
R9214 VOUT.n41 VOUT.t3 1.082
R9215 VOUT.n45 VOUT.t0 1.082
R9216 VOUT.n49 VOUT.t8 1.082
R9217 VOUT.n53 VOUT.t19 1.082
R9218 VOUT.n57 VOUT.t22 1.082
R9219 VOUT.n61 VOUT.t30 1.082
R9220 VOUT.n65 VOUT.t33 1.082
R9221 VOUT.n69 VOUT.t36 1.082
R9222 VOUT.n56 VOUT.n52 0.991417
R9223 VOUT.n36 VOUT.t16 0.90575
R9224 VOUT.n39 VOUT.t9 0.90575
R9225 VOUT.n43 VOUT.t1 0.90575
R9226 VOUT.n47 VOUT.t42 0.90575
R9227 VOUT.n51 VOUT.t7 0.90575
R9228 VOUT.n55 VOUT.t20 0.90575
R9229 VOUT.n59 VOUT.t23 0.90575
R9230 VOUT.n63 VOUT.t31 0.90575
R9231 VOUT.n67 VOUT.t34 0.90575
R9232 VOUT.n71 VOUT.t37 0.90575
R9233 VOUT VOUT.n77 0.871333
R9234 VOUT VOUT.n106 0.846333
R9235 VOUT.n75 VOUT.n74 0.7505
R9236 VOUT.n34 VOUT.t4 0.7295
R9237 VOUT.n35 VOUT.t43 0.7295
R9238 VOUT.n37 VOUT.t6 0.7295
R9239 VOUT.n38 VOUT.t2 0.7295
R9240 VOUT.n41 VOUT.t10 0.7295
R9241 VOUT.n42 VOUT.t5 0.7295
R9242 VOUT.n45 VOUT.t15 0.7295
R9243 VOUT.n46 VOUT.t13 0.7295
R9244 VOUT.n49 VOUT.t14 0.7295
R9245 VOUT.n50 VOUT.t12 0.7295
R9246 VOUT.n53 VOUT.t32 0.7295
R9247 VOUT.n54 VOUT.t26 0.7295
R9248 VOUT.n57 VOUT.t35 0.7295
R9249 VOUT.n58 VOUT.t28 0.7295
R9250 VOUT.n61 VOUT.t25 0.7295
R9251 VOUT.n62 VOUT.t18 0.7295
R9252 VOUT.n65 VOUT.t27 0.7295
R9253 VOUT.n66 VOUT.t21 0.7295
R9254 VOUT.n69 VOUT.t29 0.7295
R9255 VOUT.n70 VOUT.t24 0.7295
R9256 VOUT.n89 VOUT.n88 0.60675
R9257 VOUT.n92 VOUT.n91 0.60675
R9258 VOUT.n99 VOUT.n98 0.60675
R9259 VOUT.n102 VOUT.n101 0.60675
R9260 VOUT.n9 VOUT.n8 0.60675
R9261 VOUT.n16 VOUT.n15 0.60675
R9262 VOUT.n19 VOUT.n18 0.60675
R9263 VOUT.n26 VOUT.n25 0.60675
R9264 VOUT.n75 VOUT 0.557646
R9265 VOUT.n85 VOUT.n84 0.538
R9266 VOUT.n86 VOUT.n81 0.538
R9267 VOUT.n95 VOUT.n94 0.538
R9268 VOUT.n96 VOUT.n79 0.538
R9269 VOUT.n105 VOUT.n104 0.538
R9270 VOUT.n5 VOUT.n4 0.538
R9271 VOUT.n12 VOUT.n11 0.538
R9272 VOUT.n13 VOUT.n2 0.538
R9273 VOUT.n22 VOUT.n21 0.538
R9274 VOUT.n23 VOUT.n0 0.538
R9275 VOUT.n44 VOUT.n40 0.495958
R9276 VOUT.n48 VOUT.n44 0.495958
R9277 VOUT.n52 VOUT.n48 0.495958
R9278 VOUT.n60 VOUT.n56 0.495958
R9279 VOUT.n64 VOUT.n60 0.495958
R9280 VOUT.n68 VOUT.n64 0.495958
R9281 VOUT.n72 VOUT.n68 0.495958
R9282 VOUT.n35 VOUT.n34 0.353
R9283 VOUT.n38 VOUT.n37 0.353
R9284 VOUT.n42 VOUT.n41 0.353
R9285 VOUT.n46 VOUT.n45 0.353
R9286 VOUT.n50 VOUT.n49 0.353
R9287 VOUT.n54 VOUT.n53 0.353
R9288 VOUT.n58 VOUT.n57 0.353
R9289 VOUT.n62 VOUT.n61 0.353
R9290 VOUT.n66 VOUT.n65 0.353
R9291 VOUT.n70 VOUT.n69 0.353
R9292 VOUT.n36 VOUT.n35 0.17675
R9293 VOUT.n39 VOUT.n38 0.17675
R9294 VOUT.n43 VOUT.n42 0.17675
R9295 VOUT.n47 VOUT.n46 0.17675
R9296 VOUT.n51 VOUT.n50 0.17675
R9297 VOUT.n55 VOUT.n54 0.17675
R9298 VOUT.n59 VOUT.n58 0.17675
R9299 VOUT.n63 VOUT.n62 0.17675
R9300 VOUT.n67 VOUT.n66 0.17675
R9301 VOUT.n71 VOUT.n70 0.17675
R9302 VOUT.n74 VOUT 0.0838333
R9303 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t8 241.536
R9304 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t6 241.536
R9305 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t13 230.363
R9306 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t16 230.155
R9307 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t17 230.155
R9308 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t11 229.369
R9309 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t5 229.369
R9310 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n0 203.923
R9311 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n7 181.496
R9312 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t14 169.237
R9313 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t10 169.237
R9314 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n5 159.37
R9315 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t15 158.064
R9316 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n17 157.927
R9317 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t12 157.856
R9318 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t4 157.856
R9319 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t7 157.07
R9320 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t9 157.07
R9321 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n11 156.655
R9322 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n2 153.529
R9323 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n18 152
R9324 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n14 152
R9325 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n23 101.49
R9326 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n21 44.3335
R9327 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n6 40.9264
R9328 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n12 29.3297
R9329 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t2 26.5955
R9330 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t3 26.5955
R9331 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t1 24.9236
R9332 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t0 24.9236
R9333 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n15 18.1923
R9334 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n20 16.335
R9335 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n3 16.0286
R9336 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 13.1418
R9337 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n22 13.0565
R9338 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n1 10.7525
R9339 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n8 9.3005
R9340 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n19 7.9365
R9341 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 6.6565
R9342 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n9 6.5302
R9343 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 5.04292
R9344 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 4.3525
R9345 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 3.49141
R9346 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.86617
R9347 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.5605
R9348 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.5605
R9349 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.3045
R9350 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.10199
R9351 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.03686
R9352 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n24 1.93989
R9353 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n10 1.39698
R9354 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n16 1.06105
R9355 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n13 0.988781
R9356 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n4 0.852062
R9357 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.338391
R9358 a_43167_3162.t0 a_43167_3162.t1 49.8467
R9359 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 272.038
R9360 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t1 258.846
R9361 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t4 228.463
R9362 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n5 224.775
R9363 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t3 157.07
R9364 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n0 153.28
R9365 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t2 26.5955
R9366 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t0 26.5955
R9367 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n1 21.3673
R9368 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n4 3.76521
R9369 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n3 3.03935
R9370 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 2.92621
R9371 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n2 1.56597
R9372 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.921363
R9373 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n2 0.737191
R9374 DIN2.n1 DIN2.t0 212.081
R9375 DIN2.n0 DIN2.t3 212.081
R9376 DIN2.n2 DIN2.n1 183.185
R9377 DIN2.n1 DIN2.t2 139.78
R9378 DIN2.n0 DIN2.t1 139.78
R9379 DIN2.n1 DIN2.n0 61.346
R9380 DIN2 DIN2.n2 14.2776
R9381 DIN2.n2 DIN2 5.8885
R9382 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t62 214.787
R9383 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t82 214.787
R9384 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t4 214.011
R9385 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t24 214.011
R9386 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n61 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t60 142.488
R9387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t18 142.488
R9388 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t83 142.488
R9389 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t14 142.488
R9390 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t77 142.488
R9391 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t26 142.488
R9392 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t10 142.488
R9393 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n75 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t79 141.704
R9394 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t12 141.704
R9395 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n77 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t59 141.704
R9396 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t55 141.704
R9397 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n79 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t15 141.704
R9398 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n80 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t40 141.704
R9399 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n81 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t51 141.704
R9400 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n82 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t72 141.704
R9401 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t22 141.704
R9402 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t54 141.704
R9403 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t87 141.704
R9404 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t85 141.704
R9405 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t38 141.704
R9406 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t63 141.704
R9407 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t36 141.704
R9408 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t33 141.704
R9409 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t58 141.704
R9410 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t17 141.704
R9411 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n61 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t41 141.704
R9412 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t31 141.704
R9413 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t81 141.704
R9414 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t78 141.704
R9415 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n55 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t32 141.704
R9416 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n56 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t57 141.704
R9417 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t73 141.704
R9418 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n58 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t13 141.704
R9419 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t39 141.704
R9420 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t75 141.704
R9421 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t23 141.704
R9422 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t21 141.704
R9423 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n47 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t52 141.704
R9424 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t86 141.704
R9425 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t50 141.704
R9426 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t48 141.704
R9427 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t80 141.704
R9428 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t35 141.704
R9429 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t61 141.704
R9430 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t27 141.704
R9431 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t76 141.704
R9432 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t71 141.704
R9433 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t28 141.704
R9434 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t53 141.704
R9435 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t69 141.704
R9436 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t11 141.704
R9437 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t37 141.704
R9438 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t70 141.704
R9439 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t20 141.704
R9440 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t19 141.704
R9441 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t49 141.704
R9442 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t84 141.704
R9443 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t46 141.704
R9444 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t45 141.704
R9445 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t74 141.704
R9446 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t29 141.704
R9447 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t56 141.704
R9448 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t42 141.704
R9449 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t9 141.704
R9450 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t7 141.704
R9451 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t43 141.704
R9452 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t67 141.704
R9453 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t5 141.704
R9454 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t25 141.704
R9455 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t47 141.704
R9456 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t6 141.704
R9457 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t34 141.704
R9458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t30 141.704
R9459 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t66 141.704
R9460 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t16 141.704
R9461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t65 141.704
R9462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t64 141.704
R9463 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t8 141.704
R9464 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t44 141.704
R9465 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t68 141.704
R9466 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n86 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n85 119.186
R9467 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n0 119.186
R9468 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n85 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t1 15.3866
R9469 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n85 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t3 15.3866
R9470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t2 15.3866
R9471 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t0 15.3866
R9472 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n86 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n1 10.5922
R9473 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n73 7.95883
R9474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n74 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 6.74425
R9475 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n87 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n84 6.37582
R9476 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n87 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n86 5.23592
R9477 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n87 5.17342
R9478 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n20 4.22517
R9479 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n75 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n74 4.13592
R9480 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n39 3.4105
R9481 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n59 3.4105
R9482 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n84 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n83 3.4105
R9483 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n74 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n72 0.973417
R9484 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n84 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n60 0.815167
R9485 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n61 0.783833
R9486 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n62 0.783833
R9487 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n63 0.783833
R9488 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n64 0.783833
R9489 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n65 0.783833
R9490 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n66 0.783833
R9491 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n67 0.783833
R9492 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n68 0.783833
R9493 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n69 0.783833
R9494 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n70 0.783833
R9495 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n82 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n81 0.783833
R9496 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n81 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n80 0.783833
R9497 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n80 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n79 0.783833
R9498 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n79 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n78 0.783833
R9499 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n77 0.783833
R9500 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n77 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n76 0.783833
R9501 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n75 0.783833
R9502 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n41 0.783833
R9503 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n42 0.783833
R9504 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n43 0.783833
R9505 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n44 0.783833
R9506 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n45 0.783833
R9507 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n47 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n46 0.783833
R9508 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n47 0.783833
R9509 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n48 0.783833
R9510 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n49 0.783833
R9511 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n50 0.783833
R9512 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n58 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n57 0.783833
R9513 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n56 0.783833
R9514 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n56 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n55 0.783833
R9515 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n55 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n54 0.783833
R9516 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n53 0.783833
R9517 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n52 0.783833
R9518 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n21 0.783833
R9519 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n22 0.783833
R9520 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n23 0.783833
R9521 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n24 0.783833
R9522 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n25 0.783833
R9523 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n26 0.783833
R9524 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n27 0.783833
R9525 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n28 0.783833
R9526 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n29 0.783833
R9527 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n30 0.783833
R9528 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n37 0.783833
R9529 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n36 0.783833
R9530 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n35 0.783833
R9531 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n34 0.783833
R9532 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n33 0.783833
R9533 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n32 0.783833
R9534 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n2 0.783833
R9535 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n3 0.783833
R9536 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n4 0.783833
R9537 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n5 0.783833
R9538 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n6 0.783833
R9539 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n7 0.783833
R9540 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n8 0.783833
R9541 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n9 0.783833
R9542 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n10 0.783833
R9543 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n11 0.783833
R9544 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n18 0.783833
R9545 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n17 0.783833
R9546 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n16 0.783833
R9547 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n15 0.783833
R9548 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n14 0.783833
R9549 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n13 0.783833
R9550 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n83 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n82 0.777583
R9551 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n58 0.777583
R9552 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n38 0.777583
R9553 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n19 0.777583
R9554 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n40 0.39003
R9555 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n1 0.063
R9556 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n83 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n71 0.00675
R9557 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n51 0.00675
R9558 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n31 0.00675
R9559 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n12 0.00675
R9560 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t9 168.994
R9561 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t7 168.994
R9562 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t6 168.375
R9563 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t8 168.375
R9564 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t2 69.6757
R9565 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t0 60.3003
R9566 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t4 59.8829
R9567 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t1 59.4176
R9568 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t5 49.8882
R9569 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t3 49.6789
R9570 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n0 12.9172
R9571 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n5 10.0151
R9572 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n7 6.413
R9573 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n1 5.5094
R9574 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n2 2.75326
R9575 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n4 1.48383
R9576 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n3 1.47967
R9577 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n6 0.8255
R9578 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21.t2 246.63
R9579 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21.t1 10.6701
R9580 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21.t0 10.5739
R9581 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21.n0 2.78018
R9582 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.t2 246.501
R9583 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.t1 10.5309
R9584 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.t0 10.5295
R9585 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.n0 2.14784
R9586 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t0 672.309
R9587 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t1 10.791
R9588 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t2 10.6937
R9589 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.n0 1.35575
R9590 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t1 672.655
R9591 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t0 10.7134
R9592 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t2 10.6712
R9593 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.n0 2.05317
R9594 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t1 334.788
R9595 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t8 213.218
R9596 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t6 212.982
R9597 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t5 212.554
R9598 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t3 212.554
R9599 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t9 208.054
R9600 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t7 126.27
R9601 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t4 125.558
R9602 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t2 121.127
R9603 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t0 87.8063
R9604 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n3 60.0689
R9605 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n6 5.73592
R9606 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n7 5.388
R9607 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n2 4.5005
R9608 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n0 0.663962
R9609 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n1 0.663962
R9610 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n4 0.322615
R9611 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.236077
R9612 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n5 0.177583
R9613 a_43240_20580.t0 a_43240_20580.t1 65.941
R9614 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t1 334.822
R9615 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t8 213.218
R9616 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t5 213.218
R9617 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t4 212.554
R9618 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t9 212.554
R9619 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t6 208.054
R9620 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t7 126.27
R9621 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t2 125.558
R9622 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t3 125.558
R9623 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t0 87.8063
R9624 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n3 63.3651
R9625 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n6 5.73592
R9626 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n7 5.66196
R9627 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n2 4.5005
R9628 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n5 0.713
R9629 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n1 0.663962
R9630 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.457231
R9631 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n0 0.207231
R9632 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n4 0.197295
R9633 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t1 334.788
R9634 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t8 213.218
R9635 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t14 213.218
R9636 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t12 212.554
R9637 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t19 212.554
R9638 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t9 212.554
R9639 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t20 212.554
R9640 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t3 212.554
R9641 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t11 212.554
R9642 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t21 212.554
R9643 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t13 212.554
R9644 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t17 212.554
R9645 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t2 212.554
R9646 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t15 212.554
R9647 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t5 212.554
R9648 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t4 212.554
R9649 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t18 212.554
R9650 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t6 212.554
R9651 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t16 126.27
R9652 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t7 125.558
R9653 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t10 121.127
R9654 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t0 87.8063
R9655 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n15 81.7495
R9656 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n18 5.73592
R9657 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n19 5.388
R9658 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n13 0.663962
R9659 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n12 0.663962
R9660 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n11 0.663962
R9661 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n10 0.663962
R9662 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n9 0.663962
R9663 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n8 0.663962
R9664 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n7 0.663962
R9665 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n0 0.663962
R9666 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n1 0.663962
R9667 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n3 0.663962
R9668 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n4 0.663962
R9669 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n5 0.663962
R9670 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n6 0.518014
R9671 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n2 0.442808
R9672 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n16 0.322615
R9673 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.221654
R9674 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n17 0.177583
R9675 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n14 0.133398
R9676 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.n0 238.819
R9677 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.t2 10.758
R9678 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.t1 10.7137
R9679 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t6 228.413
R9680 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t37 228.413
R9681 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t4 228.413
R9682 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t0 228.413
R9683 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t39 227.093
R9684 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t11 227.093
R9685 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t10 227.093
R9686 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t34 227.093
R9687 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t36 227.093
R9688 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t8 227.093
R9689 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t1 227.093
R9690 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t9 227.093
R9691 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t2 227.093
R9692 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t33 227.093
R9693 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t7 224.073
R9694 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t35 224.073
R9695 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t27 221.974
R9696 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t20 221.974
R9697 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t15 221.911
R9698 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t14 221.911
R9699 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t23 221.911
R9700 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t17 221.911
R9701 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t28 221.911
R9702 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t21 221.911
R9703 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t30 221.911
R9704 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t32 221.911
R9705 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t18 221.911
R9706 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t26 221.911
R9707 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t24 221.911
R9708 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t25 221.911
R9709 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t22 221.911
R9710 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t13 221.911
R9711 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t3 221.851
R9712 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t38 221.851
R9713 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t5 221.851
R9714 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t12 221.851
R9715 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t16 221.851
R9716 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t19 221.851
R9717 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t31 221.851
R9718 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t29 221.851
R9719 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n33 7.90675
R9720 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n28 7.90675
R9721 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n21 7.90675
R9722 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n24 7.90675
R9723 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n3 5.2428
R9724 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n10 5.2428
R9725 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n8 5.17941
R9726 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n34 4.77342
R9727 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n29 4.77342
R9728 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n25 4.77342
R9729 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n22 4.77342
R9730 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n27 4.55274
R9731 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n36 3.4105
R9732 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n17 3.4105
R9733 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n35 3.00675
R9734 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n11 1.813
R9735 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n14 1.813
R9736 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n0 1.813
R9737 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n6 1.813
R9738 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n4 1.813
R9739 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n2 1.70775
R9740 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n9 1.70775
R9741 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n23 1.69425
R9742 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n31 1.65556
R9743 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n19 1.65556
R9744 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n26 1.44008
R9745 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n12 1.32133
R9746 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n15 1.32133
R9747 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n5 1.32133
R9748 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n13 1.03383
R9749 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n1 0.788
R9750 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n16 0.779667
R9751 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n7 0.533833
R9752 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n18 0.216985
R9753 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n30 0.127583
R9754 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n37 0.111591
R9755 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n32 0.0619583
R9756 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n20 0.0619583
R9757 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t18 93.2073
R9758 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t17 83.2414
R9759 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t9 83.2414
R9760 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t6 83.2414
R9761 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t14 83.2414
R9762 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t22 83.2414
R9763 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t11 83.2221
R9764 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t5 83.2221
R9765 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t15 83.2221
R9766 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t23 83.2221
R9767 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n6 66.665
R9768 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n5 66.665
R9769 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n4 66.665
R9770 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n3 66.665
R9771 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n2 66.665
R9772 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t2 55.7445
R9773 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t3 55.4987
R9774 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t0 50.8843
R9775 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t1 49.6518
R9776 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n25 25.8797
R9777 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t19 16.5305
R9778 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t16 16.5305
R9779 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t8 16.5305
R9780 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t10 16.5305
R9781 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t4 16.5305
R9782 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t7 16.5305
R9783 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t13 16.5305
R9784 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t12 16.5305
R9785 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t21 16.5305
R9786 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t20 16.5305
R9787 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n10 9.98569
R9788 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n14 9.98569
R9789 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n18 9.98569
R9790 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n22 9.98569
R9791 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n0 7.99425
R9792 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n1 7.27133
R9793 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n26 6.8255
R9794 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n9 6.00467
R9795 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n13 6.00467
R9796 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n17 6.00467
R9797 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n21 6.00467
R9798 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n8 4.5005
R9799 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n12 4.5005
R9800 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n16 4.5005
R9801 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n20 4.5005
R9802 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n24 4.5005
R9803 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n7 1.06361
R9804 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n11 1.06361
R9805 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n15 1.06361
R9806 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n19 1.06361
R9807 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n23 1.06361
R9808 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.04425
R9809 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.04425
R9810 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.04425
R9811 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.04425
R9812 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.04425
R9813 a_6923_9707.n0 a_6923_9707.t4 221.913
R9814 a_6923_9707.n14 a_6923_9707.t2 221.913
R9815 a_6923_9707.n0 a_6923_9707.t1 221.911
R9816 a_6923_9707.n14 a_6923_9707.t16 221.911
R9817 a_6923_9707.n32 a_6923_9707.t7 221.851
R9818 a_6923_9707.n2 a_6923_9707.t5 221.851
R9819 a_6923_9707.n3 a_6923_9707.t15 221.851
R9820 a_6923_9707.n29 a_6923_9707.t8 221.851
R9821 a_6923_9707.n28 a_6923_9707.t18 221.851
R9822 a_6923_9707.n16 a_6923_9707.t10 221.851
R9823 a_6923_9707.n17 a_6923_9707.t6 221.851
R9824 a_6923_9707.n20 a_6923_9707.t9 221.851
R9825 a_6923_9707.n21 a_6923_9707.t17 221.851
R9826 a_6923_9707.n23 a_6923_9707.t19 221.851
R9827 a_6923_9707.n13 a_6923_9707.t3 221.851
R9828 a_6923_9707.t0 a_6923_9707.n33 221.851
R9829 a_6923_9707.n8 a_6923_9707.n7 71.3963
R9830 a_6923_9707.n8 a_6923_9707.n6 71.3963
R9831 a_6923_9707.n11 a_6923_9707.n10 71.3963
R9832 a_6923_9707.n11 a_6923_9707.n9 71.3963
R9833 a_6923_9707.n7 a_6923_9707.t20 16.5305
R9834 a_6923_9707.n7 a_6923_9707.t13 16.5305
R9835 a_6923_9707.n6 a_6923_9707.t12 16.5305
R9836 a_6923_9707.n6 a_6923_9707.t23 16.5305
R9837 a_6923_9707.n10 a_6923_9707.t14 16.5305
R9838 a_6923_9707.n10 a_6923_9707.t21 16.5305
R9839 a_6923_9707.n9 a_6923_9707.t22 16.5305
R9840 a_6923_9707.n9 a_6923_9707.t11 16.5305
R9841 a_6923_9707.n27 a_6923_9707.n26 6.69433
R9842 a_6923_9707.n15 a_6923_9707.n14 5.57739
R9843 a_6923_9707.n1 a_6923_9707.n0 5.57739
R9844 a_6923_9707.n25 a_6923_9707.n13 5.49597
R9845 a_6923_9707.n4 a_6923_9707.n3 5.31889
R9846 a_6923_9707.n2 a_6923_9707.n1 5.31889
R9847 a_6923_9707.n33 a_6923_9707.n5 5.31889
R9848 a_6923_9707.n28 a_6923_9707.n27 5.31889
R9849 a_6923_9707.n30 a_6923_9707.n29 5.31889
R9850 a_6923_9707.n16 a_6923_9707.n15 5.31889
R9851 a_6923_9707.n18 a_6923_9707.n17 5.31889
R9852 a_6923_9707.n20 a_6923_9707.n19 5.31889
R9853 a_6923_9707.n22 a_6923_9707.n21 5.31889
R9854 a_6923_9707.n24 a_6923_9707.n23 5.31889
R9855 a_6923_9707.n32 a_6923_9707.n31 5.31889
R9856 a_6923_9707.n26 a_6923_9707.n12 4.0215
R9857 a_6923_9707.n26 a_6923_9707.n25 3.4105
R9858 a_6923_9707.n24 a_6923_9707.n22 2.888
R9859 a_6923_9707.n19 a_6923_9707.n18 2.888
R9860 a_6923_9707.n31 a_6923_9707.n30 2.888
R9861 a_6923_9707.n5 a_6923_9707.n4 2.888
R9862 a_6923_9707.n12 a_6923_9707.n8 0.3505
R9863 a_6923_9707.n12 a_6923_9707.n11 0.3505
R9864 a_6923_9707.n22 a_6923_9707.n19 0.246333
R9865 a_6923_9707.n18 a_6923_9707.n15 0.246333
R9866 a_6923_9707.n30 a_6923_9707.n27 0.246333
R9867 a_6923_9707.n31 a_6923_9707.n5 0.246333
R9868 a_6923_9707.n4 a_6923_9707.n1 0.246333
R9869 a_6923_9707.n3 a_6923_9707.n2 0.123417
R9870 a_6923_9707.n29 a_6923_9707.n28 0.123417
R9871 a_6923_9707.n17 a_6923_9707.n16 0.123417
R9872 a_6923_9707.n21 a_6923_9707.n20 0.123417
R9873 a_6923_9707.n23 a_6923_9707.n13 0.123417
R9874 a_6923_9707.n33 a_6923_9707.n32 0.123417
R9875 a_6923_9707.n25 a_6923_9707.n24 0.06925
R9876 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t0 232.294
R9877 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t1 222.117
R9878 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t11 139.66
R9879 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t4 139.454
R9880 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t2 139.454
R9881 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n25 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t17 139.206
R9882 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t13 139.206
R9883 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t9 139.206
R9884 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t7 139.206
R9885 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t27 139.206
R9886 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t24 139.206
R9887 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t21 139.206
R9888 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t18 139.206
R9889 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t16 139.206
R9890 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t10 139.206
R9891 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t8 139.206
R9892 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t28 139.206
R9893 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t25 139.206
R9894 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t22 139.206
R9895 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t14 139.206
R9896 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t12 139.206
R9897 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t26 139.206
R9898 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t6 139.206
R9899 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t20 139.206
R9900 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t19 139.206
R9901 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t15 139.206
R9902 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t5 135.197
R9903 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t3 134.625
R9904 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t23 17.157
R9905 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n27 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n26 13.2737
R9906 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n27 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n4 6.81925
R9907 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n2 4.5005
R9908 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n27 4.44425
R9909 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n3 1.10467
R9910 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n24 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R9911 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n23 0.804667
R9912 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R9913 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n21 0.804667
R9914 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R9915 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n19 0.804667
R9916 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R9917 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n17 0.804667
R9918 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R9919 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n15 0.804667
R9920 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R9921 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n13 0.804667
R9922 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R9923 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n11 0.804667
R9924 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R9925 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n9 0.804667
R9926 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R9927 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n7 0.804667
R9928 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R9929 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n5 0.804667
R9930 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n0 0.701587
R9931 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n25 0.660917
R9932 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n1 0.51454
R9933 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n25 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n24 0.454667
R9934 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n22 0.454667
R9935 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n20 0.454667
R9936 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n18 0.454667
R9937 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n16 0.454667
R9938 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n14 0.454667
R9939 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n12 0.454667
R9940 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n10 0.454667
R9941 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n8 0.454667
R9942 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n6 0.454667
R9943 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.01925
R9944 a_43724_8936.t0 a_43724_8936.t1 55.3905
R9945 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n1 863.124
R9946 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n0 585
R9947 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t0 495.469
R9948 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t4 217.555
R9949 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t2 216.893
R9950 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t6 212.393
R9951 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n7 152
R9952 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t1 141.189
R9953 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t0 140.738
R9954 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t3 114.031
R9955 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t5 81.5883
R9956 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n6 76.1359
R9957 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 16.7132
R9958 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 13.7979
R9959 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 13.1884
R9960 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 11.6369
R9961 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 10.1408
R9962 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n3 7.94225
R9963 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 6.14988
R9964 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n5 4.5005
R9965 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 2.16154
R9966 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 2.16154
R9967 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n8 1.16414
R9968 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n2 0.665435
R9969 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n4 0.663962
R9970 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n9 0.582318
R9971 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.272135
R9972 a_15618_18696.t0 a_15618_18696.n0 671.716
R9973 a_15618_18696.n0 a_15618_18696.t1 667.361
R9974 a_15618_18696.n0 a_15618_18696.t2 666.032
R9975 a_18284_18696.n0 a_18284_18696.t2 672.731
R9976 a_18284_18696.n0 a_18284_18696.t1 671.336
R9977 a_18284_18696.t0 a_18284_18696.n0 660.739
R9978 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34.n0 237.841
R9979 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34.t2 10.7808
R9980 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34.t1 10.6951
R9981 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33.n0 237.419
R9982 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33.t2 10.6247
R9983 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33.t1 10.5285
R9984 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t1 334.771
R9985 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t3 213.218
R9986 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t20 213.218
R9987 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t12 213.218
R9988 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t4 212.899
R9989 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t10 212.554
R9990 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t7 212.554
R9991 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t15 212.554
R9992 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t2 212.554
R9993 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t22 212.554
R9994 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t5 212.554
R9995 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t19 212.554
R9996 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t17 212.554
R9997 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t21 212.554
R9998 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t11 212.554
R9999 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t8 212.554
R10000 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t13 208.054
R10001 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t14 208.054
R10002 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t16 208.054
R10003 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n22 152
R10004 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t24 131.306
R10005 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t18 126.278
R10006 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t23 125.566
R10007 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t6 114.031
R10008 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t0 87.8231
R10009 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t9 81.5883
R10010 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n21 34.7422
R10011 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n4 31.4317
R10012 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n20 28.8753
R10013 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 14.6403
R10014 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n23 11.4706
R10015 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n3 5.12863
R10016 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 4.82021
R10017 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n1 4.68383
R10018 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n11 4.5005
R10019 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n18 4.5005
R10020 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 4.48881
R10021 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n19 2.63367
R10022 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n24 1.01821
R10023 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.7755
R10024 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n5 0.663962
R10025 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n6 0.663962
R10026 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n7 0.663962
R10027 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n8 0.663962
R10028 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n9 0.663962
R10029 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n10 0.663962
R10030 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n17 0.663962
R10031 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n16 0.663962
R10032 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n15 0.663962
R10033 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n14 0.663962
R10034 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n13 0.663962
R10035 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n0 0.608192
R10036 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n12 0.34425
R10037 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.269731
R10038 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n2 0.177583
R10039 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28.t0 249.328
R10040 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28.t1 10.5296
R10041 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28.t2 10.5285
R10042 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28.n0 2.13671
R10043 a_31042_7686.n2 a_31042_7686.t2 246.612
R10044 a_31042_7686.n0 a_31042_7686.t4 242.863
R10045 a_31042_7686.n0 a_31042_7686.t1 239.639
R10046 a_31042_7686.n1 a_31042_7686.t3 239.326
R10047 a_31042_7686.t0 a_31042_7686.n2 239.326
R10048 a_31042_7686.n2 a_31042_7686.n1 6.788
R10049 a_31042_7686.n1 a_31042_7686.n0 3.04425
R10050 a_36888_19786.t0 a_36888_19786.n4 239.399
R10051 a_36888_19786.n4 a_36888_19786.t1 227.651
R10052 a_36888_19786.n0 a_36888_19786.t5 222.332
R10053 a_36888_19786.n2 a_36888_19786.t3 222.332
R10054 a_36888_19786.n1 a_36888_19786.t7 111.007
R10055 a_36888_19786.n3 a_36888_19786.t6 111.007
R10056 a_36888_19786.n0 a_36888_19786.t4 108.365
R10057 a_36888_19786.n2 a_36888_19786.t2 108.365
R10058 a_36888_19786.n1 a_36888_19786.n0 2.64217
R10059 a_36888_19786.n3 a_36888_19786.n2 2.64217
R10060 a_36888_19786.n3 a_36888_19786.n1 0.817167
R10061 a_36888_19786.n4 a_36888_19786.n3 0.302583
R10062 a_36888_19550.n1 a_36888_19550.t1 239.831
R10063 a_36888_19550.t0 a_36888_19550.n1 226.853
R10064 a_36888_19550.n0 a_36888_19550.t2 223.633
R10065 a_36888_19550.n0 a_36888_19550.t3 221.851
R10066 a_36888_19550.n1 a_36888_19550.n0 5.73071
R10067 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t3 232.214
R10068 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n0 191.1
R10069 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t4 159.915
R10070 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n1 152
R10071 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t1 140.53
R10072 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n3 46.4787
R10073 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n2 36.7299
R10074 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t0 26.5955
R10075 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t2 26.5955
R10076 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 16.5652
R10077 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n4 9.03579
R10078 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 2.27147
R10079 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 1.72748
R10080 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.t2 237.611
R10081 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.n1 237.554
R10082 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.t1 10.6569
R10083 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.t3 10.6569
R10084 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32.n0 3.36262
R10085 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31.n0 237.343
R10086 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31.t1 10.6247
R10087 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31.t2 10.5285
R10088 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t1 334.771
R10089 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t15 213.218
R10090 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t5 212.554
R10091 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t11 212.554
R10092 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t16 212.554
R10093 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t6 212.554
R10094 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t18 212.554
R10095 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t4 212.554
R10096 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t10 212.554
R10097 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t20 212.554
R10098 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t8 212.554
R10099 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t17 212.554
R10100 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t21 212.554
R10101 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t12 212.554
R10102 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t19 212.554
R10103 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t7 212.554
R10104 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t13 212.554
R10105 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t2 212.554
R10106 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t9 131.306
R10107 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t3 126.278
R10108 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t14 125.566
R10109 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t0 87.8231
R10110 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n16 71.2205
R10111 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n20 5.12863
R10112 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n18 4.68383
R10113 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n14 0.663962
R10114 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n13 0.663962
R10115 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n12 0.663962
R10116 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n11 0.663962
R10117 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n10 0.663962
R10118 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n9 0.663962
R10119 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n8 0.663962
R10120 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n0 0.663962
R10121 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n1 0.663962
R10122 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n2 0.663962
R10123 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n3 0.663962
R10124 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n4 0.663962
R10125 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n5 0.663962
R10126 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n6 0.663962
R10127 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n17 0.608192
R10128 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n7 0.542052
R10129 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.238481
R10130 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n19 0.177583
R10131 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n15 0.10936
R10132 a_24963_20174.n0 a_24963_20174.t1 250.252
R10133 a_24963_20174.t0 a_24963_20174.n1 245.975
R10134 a_24963_20174.n1 a_24963_20174.t2 240.382
R10135 a_24963_20174.n0 a_24963_20174.t3 240.165
R10136 a_24963_20174.n1 a_24963_20174.n0 4.27758
R10137 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.t2 240.311
R10138 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.n0 10.6068
R10139 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.t1 10.599
R10140 top_DAC_0/top_final_switch_0.VOUT[0].n2 top_DAC_0/top_final_switch_0.VOUT[0].n0 603.66
R10141 top_DAC_0/top_final_switch_0.VOUT[0].n2 top_DAC_0/top_final_switch_0.VOUT[0].n1 202.21
R10142 top_DAC_0/top_final_switch_0.VOUT[0].n3 top_DAC_0/top_final_switch_0.VOUT[0].t7 172.237
R10143 top_DAC_0/top_final_switch_0.VOUT[0].n4 top_DAC_0/top_final_switch_0.VOUT[0].t11 171.161
R10144 top_DAC_0/top_final_switch_0.VOUT[0].n3 top_DAC_0/top_final_switch_0.VOUT[0].t5 170.625
R10145 top_DAC_0/top_final_switch_0.VOUT[0].n4 top_DAC_0/top_final_switch_0.VOUT[0].t10 170.625
R10146 top_DAC_0/top_final_switch_0.VOUT[0].n7 top_DAC_0/top_final_switch_0.VOUT[0].t6 121.868
R10147 top_DAC_0/top_final_switch_0.VOUT[0].n6 top_DAC_0/top_final_switch_0.VOUT[0].t9 120.793
R10148 top_DAC_0/top_final_switch_0.VOUT[0].n7 top_DAC_0/top_final_switch_0.VOUT[0].t4 120.255
R10149 top_DAC_0/top_final_switch_0.VOUT[0].n6 top_DAC_0/top_final_switch_0.VOUT[0].t8 120.255
R10150 top_DAC_0/top_final_switch_0.VOUT[0].n0 top_DAC_0/top_final_switch_0.VOUT[0].t2 65.941
R10151 top_DAC_0/top_final_switch_0.VOUT[0].n0 top_DAC_0/top_final_switch_0.VOUT[0].t3 65.941
R10152 top_DAC_0/top_final_switch_0.VOUT[0].n1 top_DAC_0/top_final_switch_0.VOUT[0].t1 39.3576
R10153 top_DAC_0/top_final_switch_0.VOUT[0].n1 top_DAC_0/top_final_switch_0.VOUT[0].t0 39.3576
R10154 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_final_switch_0.VOUT[0].n9 18.838
R10155 top_DAC_0/top_final_switch_0.VOUT[0].n5 top_DAC_0/top_final_switch_0.VOUT[0].n3 8.69842
R10156 top_DAC_0/top_final_switch_0.VOUT[0].n8 top_DAC_0/top_final_switch_0.VOUT[0].n6 7.53592
R10157 top_DAC_0/top_final_switch_0.VOUT[0].n10 top_DAC_0/top_final_switch_0.VOUT[0] 6.22508
R10158 top_DAC_0/top_final_switch_0.VOUT[0].n5 top_DAC_0/top_final_switch_0.VOUT[0].n4 5.82758
R10159 top_DAC_0/top_final_switch_0.VOUT[0].n8 top_DAC_0/top_final_switch_0.VOUT[0].n7 5.29008
R10160 top_DAC_0/top_final_switch_0.VOUT[0].n9 top_DAC_0/top_final_switch_0.VOUT[0].n5 1.31717
R10161 top_DAC_0/top_final_switch_0.VOUT[0].n9 top_DAC_0/top_final_switch_0.VOUT[0].n8 0.4005
R10162 top_DAC_0/top_final_switch_0.VOUT[0].n10 top_DAC_0/top_final_switch_0.VOUT[0].n2 0.233364
R10163 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_final_switch_0.VOUT[0].n10 0.0275606
R10164 a_5050_12595.n3 a_5050_12595.t5 238.363
R10165 a_5050_12595.n3 a_5050_12595.t4 237.559
R10166 a_5050_12595.n6 a_5050_12595.n5 71.3963
R10167 a_5050_12595.n2 a_5050_12595.n1 71.3963
R10168 a_5050_12595.n2 a_5050_12595.n0 71.3963
R10169 a_5050_12595.n7 a_5050_12595.n6 71.3963
R10170 a_5050_12595.n5 a_5050_12595.t6 16.5305
R10171 a_5050_12595.n5 a_5050_12595.t2 16.5305
R10172 a_5050_12595.n1 a_5050_12595.t0 16.5305
R10173 a_5050_12595.n1 a_5050_12595.t8 16.5305
R10174 a_5050_12595.n0 a_5050_12595.t9 16.5305
R10175 a_5050_12595.n0 a_5050_12595.t1 16.5305
R10176 a_5050_12595.t3 a_5050_12595.n7 16.5305
R10177 a_5050_12595.n7 a_5050_12595.t7 16.5305
R10178 a_5050_12595.n4 a_5050_12595.n3 5.18724
R10179 a_5050_12595.n6 a_5050_12595.n4 0.3505
R10180 a_5050_12595.n4 a_5050_12595.n2 0.3505
R10181 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t1 227.856
R10182 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n2 152.333
R10183 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t2 140.382
R10184 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t3 114.031
R10185 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t0 83.3993
R10186 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t4 81.5883
R10187 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n3 14.4422
R10188 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n1 7.56882
R10189 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n0 5.08175
R10190 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R10191 a_43724_15312.t0 a_43724_15312.t1 55.3905
R10192 a_43698_14716.t0 a_43698_14716.n0 228.04
R10193 a_43698_14716.n0 a_43698_14716.t2 145.648
R10194 a_43698_14716.n0 a_43698_14716.t1 83.2159
R10195 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11.t2 248.95
R10196 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11.t1 10.5761
R10197 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11.t0 10.5739
R10198 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11.n0 2.84608
R10199 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.t1 249.594
R10200 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.t2 10.5307
R10201 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.t0 10.5295
R10202 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.n0 2.17402
R10203 top_DAC_0/top_final_switch_0.VOUT[4].n2 top_DAC_0/top_final_switch_0.VOUT[4].n0 603.644
R10204 top_DAC_0/top_final_switch_0.VOUT[4].n2 top_DAC_0/top_final_switch_0.VOUT[4].n1 202.21
R10205 top_DAC_0/top_final_switch_0.VOUT[4].n3 top_DAC_0/top_final_switch_0.VOUT[4].t9 172.237
R10206 top_DAC_0/top_final_switch_0.VOUT[4].n4 top_DAC_0/top_final_switch_0.VOUT[4].t11 171.161
R10207 top_DAC_0/top_final_switch_0.VOUT[4].n3 top_DAC_0/top_final_switch_0.VOUT[4].t7 170.625
R10208 top_DAC_0/top_final_switch_0.VOUT[4].n4 top_DAC_0/top_final_switch_0.VOUT[4].t5 170.625
R10209 top_DAC_0/top_final_switch_0.VOUT[4].n7 top_DAC_0/top_final_switch_0.VOUT[4].t8 121.868
R10210 top_DAC_0/top_final_switch_0.VOUT[4].n6 top_DAC_0/top_final_switch_0.VOUT[4].t10 120.793
R10211 top_DAC_0/top_final_switch_0.VOUT[4].n7 top_DAC_0/top_final_switch_0.VOUT[4].t6 120.255
R10212 top_DAC_0/top_final_switch_0.VOUT[4].n6 top_DAC_0/top_final_switch_0.VOUT[4].t4 120.255
R10213 top_DAC_0/top_final_switch_0.VOUT[4].n0 top_DAC_0/top_final_switch_0.VOUT[4].t2 65.941
R10214 top_DAC_0/top_final_switch_0.VOUT[4].n0 top_DAC_0/top_final_switch_0.VOUT[4].t3 65.941
R10215 top_DAC_0/top_final_switch_0.VOUT[4].n1 top_DAC_0/top_final_switch_0.VOUT[4].t1 39.3576
R10216 top_DAC_0/top_final_switch_0.VOUT[4].n1 top_DAC_0/top_final_switch_0.VOUT[4].t0 39.3576
R10217 top_DAC_0/top_final_switch_0.VOUT[4].n5 top_DAC_0/top_final_switch_0.VOUT[4].n3 8.69842
R10218 top_DAC_0/top_final_switch_0.VOUT[4].n8 top_DAC_0/top_final_switch_0.VOUT[4].n6 7.53592
R10219 top_DAC_0/top_final_switch_0.VOUT[4].n11 top_DAC_0/top_final_switch_0.VOUT[4].n10 6.56586
R10220 top_DAC_0/top_final_switch_0.VOUT[4].n5 top_DAC_0/top_final_switch_0.VOUT[4].n4 5.82758
R10221 top_DAC_0/top_final_switch_0.VOUT[4].n8 top_DAC_0/top_final_switch_0.VOUT[4].n7 5.29008
R10222 top_DAC_0/top_final_switch_0.VOUT[4].n10 top_DAC_0/top_final_switch_0.VOUT[4].n9 4.5005
R10223 top_DAC_0/top_final_switch_0.VOUT[4].n9 top_DAC_0/top_final_switch_0.VOUT[4].n8 1.13383
R10224 top_DAC_0/top_final_switch_0.VOUT[4].n9 top_DAC_0/top_final_switch_0.VOUT[4].n5 0.583833
R10225 top_DAC_0/top_final_switch_0.VOUT[4].n11 top_DAC_0/top_final_switch_0.VOUT[4].n2 0.23296
R10226 top_DAC_0/top_final_switch_0.VOUT[4].n10 top_DAC_0/top_final_switch_0.VOUT[4] 0.063
R10227 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_final_switch_0.VOUT[4].n11 0.0275606
R10228 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45.n0 238.496
R10229 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45.t1 10.7258
R10230 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45.t2 10.6617
R10231 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t7 141.129
R10232 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t4 141.129
R10233 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t5 139.808
R10234 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t6 139.808
R10235 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t1 134.732
R10236 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t2 134.732
R10237 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t0 134.732
R10238 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n5 134.732
R10239 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n4 9.87092
R10240 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n0 9.44517
R10241 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n1 5.85274
R10242 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n2 3.923
R10243 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n3 1.25383
R10244 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t1 334.822
R10245 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t17 213.218
R10246 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t5 213.218
R10247 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t15 213.218
R10248 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t6 212.864
R10249 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t12 212.554
R10250 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t10 212.554
R10251 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t7 212.554
R10252 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t13 212.554
R10253 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t4 212.554
R10254 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t23 212.554
R10255 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t20 212.554
R10256 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t24 212.554
R10257 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t14 212.554
R10258 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t21 212.554
R10259 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t11 212.554
R10260 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t16 208.054
R10261 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t2 208.054
R10262 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t8 208.054
R10263 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n21 152
R10264 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t9 126.27
R10265 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t3 125.558
R10266 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t22 125.558
R10267 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t18 114.031
R10268 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t0 87.8063
R10269 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t19 81.5883
R10270 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n4 47.4151
R10271 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n20 21.8672
R10272 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 13.9702
R10273 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 12.6356
R10274 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n22 11.4706
R10275 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n2 5.73592
R10276 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n3 5.66196
R10277 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 4.85387
R10278 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n16 4.5005
R10279 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n18 4.5005
R10280 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 4.48881
R10281 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n17 2.588
R10282 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n23 1.02238
R10283 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.7755
R10284 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n1 0.713
R10285 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n15 0.663962
R10286 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n14 0.663962
R10287 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n13 0.663962
R10288 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n12 0.663962
R10289 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n11 0.663962
R10290 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n5 0.663962
R10291 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n6 0.663962
R10292 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n7 0.663962
R10293 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n8 0.663962
R10294 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n9 0.663962
R10295 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n10 0.663962
R10296 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n19 0.311626
R10297 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n0 0.197295
R10298 a_29780_7686.n2 a_29780_7686.t4 245.879
R10299 a_29780_7686.n0 a_29780_7686.t2 241.619
R10300 a_29780_7686.n0 a_29780_7686.t1 240.234
R10301 a_29780_7686.n1 a_29780_7686.t3 238.593
R10302 a_29780_7686.t0 a_29780_7686.n2 238.593
R10303 a_29780_7686.n2 a_29780_7686.n1 6.788
R10304 a_29780_7686.n1 a_29780_7686.n0 4.94008
R10305 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.t0 249.738
R10306 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.t1 13.4579
R10307 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.t2 10.7848
R10308 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.n0 4.72836
R10309 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31.t1 240.469
R10310 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31.t2 10.6701
R10311 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31.n0 10.5739
R10312 a_31870_7686.n2 a_31870_7686.t3 247.161
R10313 a_31870_7686.n0 a_31870_7686.t2 244.589
R10314 a_31870_7686.n0 a_31870_7686.t1 240.337
R10315 a_31870_7686.n1 a_31870_7686.t4 239.875
R10316 a_31870_7686.t0 a_31870_7686.n2 239.875
R10317 a_31870_7686.n2 a_31870_7686.n1 6.788
R10318 a_31870_7686.n1 a_31870_7686.n0 1.86925
R10319 top_DAC_0/top_rseg_n_dcell_0.SH[3].n2 top_DAC_0/top_rseg_n_dcell_0.SH[3].n1 863.124
R10320 top_DAC_0/top_rseg_n_dcell_0.SH[3].n1 top_DAC_0/top_rseg_n_dcell_0.SH[3].n0 585
R10321 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.SH[3].t0 495.469
R10322 top_DAC_0/top_rseg_n_dcell_0.SH[3].n4 top_DAC_0/top_rseg_n_dcell_0.SH[3].t3 213.375
R10323 top_DAC_0/top_rseg_n_dcell_0.SH[3].n7 top_DAC_0/top_rseg_n_dcell_0.SH[3].t5 212.393
R10324 top_DAC_0/top_rseg_n_dcell_0.SH[3].n6 top_DAC_0/top_rseg_n_dcell_0.SH[3].t2 212.393
R10325 top_DAC_0/top_rseg_n_dcell_0.SH[3].n5 top_DAC_0/top_rseg_n_dcell_0.SH[3].t4 212.393
R10326 top_DAC_0/top_rseg_n_dcell_0.SH[3].n4 top_DAC_0/top_rseg_n_dcell_0.SH[3].t6 212.393
R10327 top_DAC_0/top_rseg_n_dcell_0.SH[3].n3 top_DAC_0/top_rseg_n_dcell_0.SH[3].t1 141.189
R10328 top_DAC_0/top_rseg_n_dcell_0.SH[3].n1 top_DAC_0/top_rseg_n_dcell_0.SH[3].t0 140.738
R10329 top_DAC_0/top_rseg_n_dcell_0.SH[3].n8 top_DAC_0/top_rseg_n_dcell_0.SH[3] 14.5776
R10330 top_DAC_0/top_rseg_n_dcell_0.SH[3].n2 top_DAC_0/top_rseg_n_dcell_0.SH[3] 11.6369
R10331 top_DAC_0/top_rseg_n_dcell_0.SH[3].n0 top_DAC_0/top_rseg_n_dcell_0.SH[3] 10.1408
R10332 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.SH[3].n8 8.14595
R10333 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.SH[3].n3 7.94225
R10334 top_DAC_0/top_rseg_n_dcell_0.SH[3].n8 top_DAC_0/top_rseg_n_dcell_0.SH[3] 6.20656
R10335 top_DAC_0/top_rseg_n_dcell_0.SH[3].n3 top_DAC_0/top_rseg_n_dcell_0.SH[3] 6.14988
R10336 top_DAC_0/top_rseg_n_dcell_0.SH[3].n0 top_DAC_0/top_rseg_n_dcell_0.SH[3] 2.16154
R10337 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.SH[3].n7 1.39101
R10338 top_DAC_0/top_rseg_n_dcell_0.SH[3].n5 top_DAC_0/top_rseg_n_dcell_0.SH[3].n4 0.982408
R10339 top_DAC_0/top_rseg_n_dcell_0.SH[3].n6 top_DAC_0/top_rseg_n_dcell_0.SH[3].n5 0.982408
R10340 top_DAC_0/top_rseg_n_dcell_0.SH[3].n7 top_DAC_0/top_rseg_n_dcell_0.SH[3].n6 0.982408
R10341 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.SH[3].n2 0.665435
R10342 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.VL3.t4 666.389
R10343 top_DAC_0/top_rseg_n_dcell_0.VL3.n2 top_DAC_0/top_rseg_n_dcell_0.VL3.t2 661.157
R10344 top_DAC_0/top_rseg_n_dcell_0.VL3.n1 top_DAC_0/top_rseg_n_dcell_0.VL3.t0 660.744
R10345 top_DAC_0/top_rseg_n_dcell_0.VL3.n5 top_DAC_0/top_rseg_n_dcell_0.VL3.t1 660.24
R10346 top_DAC_0/top_rseg_n_dcell_0.VL3.n4 top_DAC_0/top_rseg_n_dcell_0.VL3.t6 660.24
R10347 top_DAC_0/top_rseg_n_dcell_0.VL3.n3 top_DAC_0/top_rseg_n_dcell_0.VL3.t5 660.24
R10348 top_DAC_0/top_rseg_n_dcell_0.VL3.n2 top_DAC_0/top_rseg_n_dcell_0.VL3.t3 660.24
R10349 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.VL3.n1 25.6261
R10350 top_DAC_0/top_rseg_n_dcell_0.VL3.n1 top_DAC_0/top_rseg_n_dcell_0.VL3.n0 4.5005
R10351 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.VL3.n5 1.53057
R10352 top_DAC_0/top_rseg_n_dcell_0.VL3.n3 top_DAC_0/top_rseg_n_dcell_0.VL3.n2 1.33338
R10353 top_DAC_0/top_rseg_n_dcell_0.VL3.n4 top_DAC_0/top_rseg_n_dcell_0.VL3.n3 0.63637
R10354 top_DAC_0/top_rseg_n_dcell_0.VL3.n5 top_DAC_0/top_rseg_n_dcell_0.VL3.n4 0.63637
R10355 top_DAC_0/top_rseg_n_dcell_0.VL3.n0 top_DAC_0/top_rseg_n_dcell_0.VL3 0.063
R10356 top_DAC_0/top_rseg_n_dcell_0.VL3.n0 top_DAC_0/top_rseg_n_dcell_0.VL3 0.013
R10357 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39.t2 248.075
R10358 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39.t1 10.575
R10359 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39.t0 10.5739
R10360 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39.n0 4.2135
R10361 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38.t1 246.885
R10362 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38.t0 10.5306
R10363 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38.t2 10.5285
R10364 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38.n0 3.53633
R10365 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n1 267.599
R10366 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t5 229.369
R10367 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n0 202.094
R10368 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t6 157.07
R10369 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n3 152
R10370 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t3 132.982
R10371 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n5 61.3652
R10372 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t4 32.5055
R10373 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t1 32.5055
R10374 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t2 26.5955
R10375 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t0 26.5955
R10376 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n4 19.8407
R10377 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 5.92643
R10378 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n6 4.04261
R10379 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n2 1.12991
R10380 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t3 146.321
R10381 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t2 144.415
R10382 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t0 143.702
R10383 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n1 143.431
R10384 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n0 0.7525
R10385 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n2 271.668
R10386 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t1 258.846
R10387 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t4 228.649
R10388 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n5 224.775
R10389 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t3 156.35
R10390 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n0 152
R10391 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n1 35.7621
R10392 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t2 26.5955
R10393 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t0 26.5955
R10394 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 6.13383
R10395 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n4 3.76521
R10396 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n3 3.03935
R10397 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 2.30266
R10398 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.921363
R10399 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.368845
R10400 a_44255_4614.t0 a_44255_4614.t1 60.9236
R10401 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t7 752.615
R10402 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n5 258.361
R10403 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t5 230.576
R10404 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n4 202.095
R10405 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t6 158.275
R10406 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n0 152
R10407 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t1 126.469
R10408 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n6 62.4946
R10409 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t2 32.5055
R10410 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t4 32.5055
R10411 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t0 26.5955
R10412 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t3 26.5955
R10413 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[2] 13.6567
R10414 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n1 12.0102
R10415 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n2 9.82192
R10416 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.A 6.66717
R10417 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n3 6.51278
R10418 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n7 4.04261
R10419 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[2] 0.853179
R10420 top_DAC_0/top_rseg_n_dcell_0.VL2.n0 top_DAC_0/top_rseg_n_dcell_0.VL2.t6 240.29
R10421 top_DAC_0/top_rseg_n_dcell_0.VL2.n1 top_DAC_0/top_rseg_n_dcell_0.VL2.t8 239.082
R10422 top_DAC_0/top_rseg_n_dcell_0.VL2.n0 top_DAC_0/top_rseg_n_dcell_0.VL2.t1 239.082
R10423 top_DAC_0/top_rseg_n_dcell_0.VL2.n4 top_DAC_0/top_rseg_n_dcell_0.VL2.t5 236.407
R10424 top_DAC_0/top_rseg_n_dcell_0.VL2.n3 top_DAC_0/top_rseg_n_dcell_0.VL2.t4 234.582
R10425 top_DAC_0/top_rseg_n_dcell_0.VL2.n6 top_DAC_0/top_rseg_n_dcell_0.VL2.t2 233.657
R10426 top_DAC_0/top_rseg_n_dcell_0.VL2.n5 top_DAC_0/top_rseg_n_dcell_0.VL2.t3 233.657
R10427 top_DAC_0/top_rseg_n_dcell_0.VL2.n4 top_DAC_0/top_rseg_n_dcell_0.VL2.t7 233.657
R10428 top_DAC_0/top_rseg_n_dcell_0.VL2.n7 top_DAC_0/top_rseg_n_dcell_0.VL2.t0 233.657
R10429 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.VL2.n3 30.513
R10430 top_DAC_0/top_rseg_n_dcell_0.VL2.n3 top_DAC_0/top_rseg_n_dcell_0.VL2.n2 4.5005
R10431 top_DAC_0/top_rseg_n_dcell_0.VL2.n1 top_DAC_0/top_rseg_n_dcell_0.VL2.n0 1.20883
R10432 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.VL2.n7 1.00675
R10433 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.VL2.n1 0.94425
R10434 top_DAC_0/top_rseg_n_dcell_0.VL2.n5 top_DAC_0/top_rseg_n_dcell_0.VL2.n4 0.63637
R10435 top_DAC_0/top_rseg_n_dcell_0.VL2.n6 top_DAC_0/top_rseg_n_dcell_0.VL2.n5 0.63637
R10436 top_DAC_0/top_rseg_n_dcell_0.VL2.n7 top_DAC_0/top_rseg_n_dcell_0.VL2.n6 0.63637
R10437 top_DAC_0/top_rseg_n_dcell_0.VL2.n2 top_DAC_0/top_rseg_n_dcell_0.VL2 0.265083
R10438 top_DAC_0/top_rseg_n_dcell_0.VL2.n2 top_DAC_0/top_rseg_n_dcell_0.VL2 0.063
R10439 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3.t2 245.726
R10440 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3.t0 10.5816
R10441 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3.t1 10.5739
R10442 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3.n0 1.48638
R10443 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4.t1 247.869
R10444 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4.t2 10.5339
R10445 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4.t0 10.5295
R10446 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4.n0 2.21785
R10447 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t21 244.881
R10448 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t23 222.089
R10449 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t1 134.738
R10450 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t16 134.738
R10451 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t0 134.738
R10452 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t15 134.738
R10453 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t19 134.734
R10454 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t11 134.734
R10455 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t17 134.734
R10456 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t18 134.734
R10457 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t9 134.734
R10458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t10 134.734
R10459 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t2 134.734
R10460 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t3 134.734
R10461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t14 134.734
R10462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t7 134.734
R10463 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t12 134.734
R10464 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t6 134.734
R10465 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t8 134.734
R10466 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t4 134.734
R10467 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t5 134.734
R10468 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t13 134.734
R10469 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t20 15.2609
R10470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t24 15.2609
R10471 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n0 11.485
R10472 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n23 11.0892
R10473 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n19 9.71425
R10474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n1 7.63383
R10475 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n10 7.63383
R10476 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n18 7.15217
R10477 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n9 6.46995
R10478 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n2 4.5005
R10479 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n4 4.5005
R10480 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n6 4.5005
R10481 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n8 4.5005
R10482 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n11 4.5005
R10483 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n13 4.5005
R10484 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n17 4.5005
R10485 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n15 4.5005
R10486 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t25 4.23377
R10487 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t22 4.23377
R10488 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n3 3.13383
R10489 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n5 3.13383
R10490 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n7 3.13383
R10491 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n12 3.13383
R10492 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n14 3.13383
R10493 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n16 3.13383
R10494 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n20 3.05467
R10495 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n21 0.965083
R10496 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n22 0.646333
R10497 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n24 0.063
R10498 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n0 194.3
R10499 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n67 194.3
R10500 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t52 135.499
R10501 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t47 135.499
R10502 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t7 134.715
R10503 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t4 134.715
R10504 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t27 111.398
R10505 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t56 111.398
R10506 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t59 111.398
R10507 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t5 111.398
R10508 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t16 111.398
R10509 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n61 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t33 111.398
R10510 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t36 111.398
R10511 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t35 110.615
R10512 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t54 110.615
R10513 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t12 110.615
R10514 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t41 110.615
R10515 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t65 110.615
R10516 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t14 110.615
R10517 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t23 110.615
R10518 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t45 110.615
R10519 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t22 110.615
R10520 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t20 110.615
R10521 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t61 110.615
R10522 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t8 110.615
R10523 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t28 110.615
R10524 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t42 110.615
R10525 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t49 110.615
R10526 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t6 110.615
R10527 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t25 110.615
R10528 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t55 110.615
R10529 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t15 110.615
R10530 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t26 110.615
R10531 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t40 110.615
R10532 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t64 110.615
R10533 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t39 110.615
R10534 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t38 110.615
R10535 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t10 110.615
R10536 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t21 110.615
R10537 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t44 110.615
R10538 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t24 110.615
R10539 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n47 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t46 110.615
R10540 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t13 110.615
R10541 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t32 110.615
R10542 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t48 110.615
R10543 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t63 110.615
R10544 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t17 110.615
R10545 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t60 110.615
R10546 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t58 110.615
R10547 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t30 110.615
R10548 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t43 110.615
R10549 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t67 110.615
R10550 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n61 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t31 110.615
R10551 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t9 110.615
R10552 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t50 110.615
R10553 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t34 110.615
R10554 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t11 110.615
R10555 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t53 110.615
R10556 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n58 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t51 110.615
R10557 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t29 110.615
R10558 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n56 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t66 110.615
R10559 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n55 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t57 110.615
R10560 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t19 110.615
R10561 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t18 110.615
R10562 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t62 110.615
R10563 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n51 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t37 110.615
R10564 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t2 27.5505
R10565 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t0 27.5505
R10566 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t1 27.5505
R10567 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t3 27.5505
R10568 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n30 13.3067
R10569 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n29 6.23592
R10570 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n28 5.8755
R10571 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n2 5.04842
R10572 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n1 5.04633
R10573 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n68 5.04633
R10574 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n73 4.98592
R10575 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n18 3.84917
R10576 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n71 3.62129
R10577 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n65 3.4105
R10578 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n49 3.4105
R10579 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n35 3.4105
R10580 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n70 3.4105
R10581 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n71 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n66 1.97948
R10582 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.860917
R10583 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n4 0.783833
R10584 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n5 0.783833
R10585 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n6 0.783833
R10586 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n7 0.783833
R10587 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n8 0.783833
R10588 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n9 0.783833
R10589 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n10 0.783833
R10590 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n11 0.783833
R10591 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n12 0.783833
R10592 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n16 0.783833
R10593 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n15 0.783833
R10594 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n14 0.783833
R10595 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n19 0.783833
R10596 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n20 0.783833
R10597 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n21 0.783833
R10598 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n22 0.783833
R10599 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n23 0.783833
R10600 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n24 0.783833
R10601 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n25 0.783833
R10602 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n26 0.783833
R10603 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n33 0.783833
R10604 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n32 0.783833
R10605 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n31 0.783833
R10606 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n37 0.783833
R10607 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n38 0.783833
R10608 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n39 0.783833
R10609 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n40 0.783833
R10610 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n41 0.783833
R10611 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n42 0.783833
R10612 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n43 0.783833
R10613 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n44 0.783833
R10614 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n48 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n47 0.783833
R10615 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n47 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n46 0.783833
R10616 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n52 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n51 0.783833
R10617 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n53 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n52 0.783833
R10618 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n53 0.783833
R10619 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n55 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n54 0.783833
R10620 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n56 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n55 0.783833
R10621 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n56 0.783833
R10622 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n58 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n57 0.783833
R10623 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n58 0.783833
R10624 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n60 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n59 0.783833
R10625 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n64 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n63 0.783833
R10626 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n63 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n62 0.783833
R10627 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n61 0.783833
R10628 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n50 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n36 0.642121
R10629 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n72 0.548417
R10630 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n2 0.548417
R10631 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n72 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n3 0.546333
R10632 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n70 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n69 0.546333
R10633 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n73 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n2 0.492167
R10634 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n3 0.492167
R10635 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n66 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n50 0.439167
R10636 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n13 0.413
R10637 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n27 0.413
R10638 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n45 0.413
R10639 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n60 0.413
R10640 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n17 0.371333
R10641 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n34 0.371333
R10642 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n48 0.371333
R10643 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n65 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n64 0.371333
R10644 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n1 0.063
R10645 top_DAC_0/top_rseg_n_dcell_0.SH[2].n2 top_DAC_0/top_rseg_n_dcell_0.SH[2].n1 863.124
R10646 top_DAC_0/top_rseg_n_dcell_0.SH[2].n1 top_DAC_0/top_rseg_n_dcell_0.SH[2].n0 585
R10647 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.SH[2].t1 495.469
R10648 top_DAC_0/top_rseg_n_dcell_0.SH[2].t0 top_DAC_0/top_rseg_n_dcell_0.SH[2] 291.983
R10649 top_DAC_0/top_rseg_n_dcell_0.SH[2].n8 top_DAC_0/top_rseg_n_dcell_0.SH[2].t0 285
R10650 top_DAC_0/top_rseg_n_dcell_0.SH[2].n3 top_DAC_0/top_rseg_n_dcell_0.SH[2].t4 209.036
R10651 top_DAC_0/top_rseg_n_dcell_0.SH[2].n6 top_DAC_0/top_rseg_n_dcell_0.SH[2].t6 208.054
R10652 top_DAC_0/top_rseg_n_dcell_0.SH[2].n5 top_DAC_0/top_rseg_n_dcell_0.SH[2].t3 208.054
R10653 top_DAC_0/top_rseg_n_dcell_0.SH[2].n4 top_DAC_0/top_rseg_n_dcell_0.SH[2].t5 208.054
R10654 top_DAC_0/top_rseg_n_dcell_0.SH[2].n3 top_DAC_0/top_rseg_n_dcell_0.SH[2].t2 208.054
R10655 top_DAC_0/top_rseg_n_dcell_0.SH[2].n1 top_DAC_0/top_rseg_n_dcell_0.SH[2].t1 140.738
R10656 top_DAC_0/top_rseg_n_dcell_0.SH[2].n7 top_DAC_0/top_rseg_n_dcell_0.SH[2] 14.5776
R10657 top_DAC_0/top_rseg_n_dcell_0.SH[2].n8 top_DAC_0/top_rseg_n_dcell_0.SH[2] 12.4126
R10658 top_DAC_0/top_rseg_n_dcell_0.SH[2].n2 top_DAC_0/top_rseg_n_dcell_0.SH[2] 11.6369
R10659 top_DAC_0/top_rseg_n_dcell_0.SH[2].n0 top_DAC_0/top_rseg_n_dcell_0.SH[2] 10.1408
R10660 top_DAC_0/top_rseg_n_dcell_0.SH[2].n7 top_DAC_0/top_rseg_n_dcell_0.SH[2] 8.14595
R10661 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.SH[2].n7 6.20656
R10662 top_DAC_0/top_rseg_n_dcell_0.SH[2].n0 top_DAC_0/top_rseg_n_dcell_0.SH[2] 2.16154
R10663 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.SH[2].n8 1.93989
R10664 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.SH[2].n6 1.30619
R10665 top_DAC_0/top_rseg_n_dcell_0.SH[2].n4 top_DAC_0/top_rseg_n_dcell_0.SH[2].n3 0.982408
R10666 top_DAC_0/top_rseg_n_dcell_0.SH[2].n5 top_DAC_0/top_rseg_n_dcell_0.SH[2].n4 0.982408
R10667 top_DAC_0/top_rseg_n_dcell_0.SH[2].n6 top_DAC_0/top_rseg_n_dcell_0.SH[2].n5 0.982408
R10668 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.SH[2].n2 0.665435
R10669 top_DAC_0/top_final_switch_0.VOUT[3].n2 top_DAC_0/top_final_switch_0.VOUT[3].n0 603.66
R10670 top_DAC_0/top_final_switch_0.VOUT[3].n2 top_DAC_0/top_final_switch_0.VOUT[3].n1 202.21
R10671 top_DAC_0/top_final_switch_0.VOUT[3].n3 top_DAC_0/top_final_switch_0.VOUT[3].t9 172.237
R10672 top_DAC_0/top_final_switch_0.VOUT[3].n4 top_DAC_0/top_final_switch_0.VOUT[3].t8 171.161
R10673 top_DAC_0/top_final_switch_0.VOUT[3].n3 top_DAC_0/top_final_switch_0.VOUT[3].t5 170.625
R10674 top_DAC_0/top_final_switch_0.VOUT[3].n4 top_DAC_0/top_final_switch_0.VOUT[3].t11 170.625
R10675 top_DAC_0/top_final_switch_0.VOUT[3].n7 top_DAC_0/top_final_switch_0.VOUT[3].t7 121.868
R10676 top_DAC_0/top_final_switch_0.VOUT[3].n6 top_DAC_0/top_final_switch_0.VOUT[3].t6 120.793
R10677 top_DAC_0/top_final_switch_0.VOUT[3].n7 top_DAC_0/top_final_switch_0.VOUT[3].t4 120.255
R10678 top_DAC_0/top_final_switch_0.VOUT[3].n6 top_DAC_0/top_final_switch_0.VOUT[3].t10 120.255
R10679 top_DAC_0/top_final_switch_0.VOUT[3].n0 top_DAC_0/top_final_switch_0.VOUT[3].t3 65.941
R10680 top_DAC_0/top_final_switch_0.VOUT[3].n0 top_DAC_0/top_final_switch_0.VOUT[3].t2 65.941
R10681 top_DAC_0/top_final_switch_0.VOUT[3].n1 top_DAC_0/top_final_switch_0.VOUT[3].t0 39.3576
R10682 top_DAC_0/top_final_switch_0.VOUT[3].n1 top_DAC_0/top_final_switch_0.VOUT[3].t1 39.3576
R10683 top_DAC_0/top_final_switch_0.VOUT[3].n5 top_DAC_0/top_final_switch_0.VOUT[3].n3 8.69842
R10684 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_final_switch_0.VOUT[3].n9 8.038
R10685 top_DAC_0/top_final_switch_0.VOUT[3].n8 top_DAC_0/top_final_switch_0.VOUT[3].n6 7.53592
R10686 top_DAC_0/top_final_switch_0.VOUT[3].n10 top_DAC_0/top_final_switch_0.VOUT[3] 6.273
R10687 top_DAC_0/top_final_switch_0.VOUT[3].n5 top_DAC_0/top_final_switch_0.VOUT[3].n4 5.82758
R10688 top_DAC_0/top_final_switch_0.VOUT[3].n8 top_DAC_0/top_final_switch_0.VOUT[3].n7 5.29008
R10689 top_DAC_0/top_final_switch_0.VOUT[3].n9 top_DAC_0/top_final_switch_0.VOUT[3].n8 0.9505
R10690 top_DAC_0/top_final_switch_0.VOUT[3].n9 top_DAC_0/top_final_switch_0.VOUT[3].n5 0.767167
R10691 top_DAC_0/top_final_switch_0.VOUT[3].n10 top_DAC_0/top_final_switch_0.VOUT[3].n2 0.233364
R10692 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_final_switch_0.VOUT[3].n10 0.0275606
R10693 a_14615_14034.n0 a_14615_14034.t1 439.543
R10694 a_14615_14034.n0 a_14615_14034.t2 39.3576
R10695 a_14615_14034.t0 a_14615_14034.n0 39.3576
R10696 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n1 863.124
R10697 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n0 585
R10698 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t0 495.469
R10699 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t2 217.555
R10700 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t7 217.042
R10701 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t10 216.893
R10702 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t4 216.893
R10703 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t11 216.63
R10704 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t5 213.218
R10705 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t6 213.218
R10706 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t3 212.554
R10707 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t8 212.393
R10708 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t9 208.054
R10709 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t1 141.189
R10710 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t0 140.738
R10711 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n9 33.8463
R10712 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n13 19.6734
R10713 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 14.3755
R10714 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 12.1234
R10715 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 11.6369
R10716 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n12 11.5776
R10717 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n8 11.5588
R10718 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 10.1408
R10719 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n14 8.53383
R10720 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n3 7.94225
R10721 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 6.14988
R10722 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 5.81868
R10723 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n7 4.5005
R10724 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n11 4.5005
R10725 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n4 3.57326
R10726 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 2.16154
R10727 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n2 0.665435
R10728 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n5 0.663962
R10729 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n6 0.663962
R10730 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.380308
R10731 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n10 0.284154
R10732 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.180788
R10733 a_18724_8950.n0 a_18724_8950.t2 670.153
R10734 a_18724_8950.t0 a_18724_8950.n0 669.817
R10735 a_18724_8950.n0 a_18724_8950.t1 666.441
R10736 a_20932_10031.n0 a_20932_10031.t1 667.659
R10737 a_20932_10031.n0 a_20932_10031.t2 665.933
R10738 a_20932_10031.t0 a_20932_10031.n0 665.299
R10739 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t7 739.449
R10740 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t6 230.155
R10741 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t8 229.369
R10742 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 203.922
R10743 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 157.927
R10744 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t4 157.856
R10745 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t5 157.07
R10746 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 152
R10747 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 101.49
R10748 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 28.9524
R10749 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t3 26.5955
R10750 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t0 26.5955
R10751 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t1 24.9236
R10752 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t2 24.9236
R10753 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 14.4113
R10754 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y 13.0565
R10755 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 12.5635
R10756 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[1] 12.4026
R10757 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y 10.7525
R10758 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.B 7.11161
R10759 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y 6.6565
R10760 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 5.04292
R10761 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 4.3525
R10762 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 2.5605
R10763 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.A 2.13383
R10764 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y 1.93989
R10765 a_45023_18840.t0 a_45023_18840.t1 49.8467
R10766 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 593.396
R10767 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 268.077
R10768 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 258.846
R10769 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 231.554
R10770 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 26.5955
R10771 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 26.5955
R10772 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 16.5652
R10773 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 9.03579
R10774 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 8.8386
R10775 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 6.02403
R10776 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 1.72748
R10777 a_24135_20174.n0 a_24135_20174.t1 249.153
R10778 a_24135_20174.n1 a_24135_20174.t2 247.62
R10779 a_24135_20174.t0 a_24135_20174.n1 241.482
R10780 a_24135_20174.n0 a_24135_20174.t3 239.065
R10781 a_24135_20174.n1 a_24135_20174.n0 1.53175
R10782 a_15098_19866.t0 a_15098_19866.n0 670.881
R10783 a_15098_19866.n0 a_15098_19866.t2 668.149
R10784 a_15098_19866.n0 a_15098_19866.t1 665.133
R10785 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.t2 240.143
R10786 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.t1 10.575
R10787 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.n0 10.5739
R10788 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.t2 239.279
R10789 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.n0 10.681
R10790 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.t1 10.5753
R10791 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t10 231.017
R10792 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t14 230.155
R10793 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t9 229.369
R10794 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t7 229.369
R10795 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t13 229.369
R10796 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t6 229.369
R10797 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t11 228.649
R10798 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n0 203.923
R10799 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t16 158.716
R10800 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n14 157.927
R10801 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t5 157.856
R10802 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t15 157.07
R10803 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t12 157.07
R10804 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t17 157.07
R10805 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t8 157.07
R10806 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t4 156.35
R10807 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n2 156.268
R10808 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n5 153.423
R10809 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n15 152
R10810 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n12 152
R10811 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n9 152
R10812 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n3 152
R10813 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n21 101.49
R10814 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 53.8309
R10815 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n19 43.993
R10816 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t2 26.5955
R10817 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t3 26.5955
R10818 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t0 24.9236
R10819 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t1 24.9236
R10820 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n10 18.4368
R10821 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n4 16.4183
R10822 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n6 14.4998
R10823 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n16 13.1513
R10824 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n20 13.0565
R10825 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n13 11.3143
R10826 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n1 10.7525
R10827 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n17 9.3005
R10828 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 7.11161
R10829 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 6.6565
R10830 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n18 6.60324
R10831 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 5.92643
R10832 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 5.92643
R10833 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 5.04292
R10834 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 4.5042
R10835 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 4.3525
R10836 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 2.5605
R10837 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 2.3045
R10838 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n22 1.93989
R10839 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 1.43334
R10840 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n8 1.13136
R10841 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n7 1.10597
R10842 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n11 0.699719
R10843 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.529797
R10844 a_43391_3326.t0 a_43391_3326.t1 60.9236
R10845 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n4 267.599
R10846 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t0 257
R10847 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t0 249
R10848 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t5 230.155
R10849 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n0 196.889
R10850 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t6 157.856
R10851 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n1 152
R10852 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n5 62.4946
R10853 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t1 32.5055
R10854 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t2 32.5055
R10855 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n2 30.2423
R10856 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t4 26.5955
R10857 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t3 26.5955
R10858 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n6 6.51278
R10859 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n3 5.2056
R10860 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n7 4.04261
R10861 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 2.3045
R10862 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t1 231.236
R10863 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t0 231.129
R10864 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t3 230.782
R10865 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t2 230.272
R10866 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n0 1.03165
R10867 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n1 0.550258
R10868 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t1 334.771
R10869 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t15 213.218
R10870 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t4 212.554
R10871 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t12 212.554
R10872 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t3 212.554
R10873 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t5 212.554
R10874 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t17 212.554
R10875 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t7 212.554
R10876 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t11 212.554
R10877 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t18 212.554
R10878 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t9 212.554
R10879 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t16 212.554
R10880 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t14 212.554
R10881 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t21 212.554
R10882 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t8 212.554
R10883 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t19 212.554
R10884 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t10 212.554
R10885 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t6 208.054
R10886 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t20 126.278
R10887 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t13 125.566
R10888 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t2 125.566
R10889 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t0 87.8568
R10890 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n16 62.8505
R10891 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n20 5.04008
R10892 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n19 4.68383
R10893 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n15 4.5005
R10894 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n17 0.876942
R10895 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n18 0.713
R10896 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n0 0.663962
R10897 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n1 0.663962
R10898 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n2 0.663962
R10899 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n3 0.663962
R10900 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n4 0.663962
R10901 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n14 0.663962
R10902 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n13 0.663962
R10903 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n12 0.663962
R10904 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n11 0.663962
R10905 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n10 0.663962
R10906 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n9 0.663962
R10907 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n8 0.663962
R10908 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n7 0.663962
R10909 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n6 0.663962
R10910 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n5 0.663962
R10911 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.209635
R10912 a_42724_21320.t0 a_42724_21320.t1 65.941
R10913 a_42982_21320.t0 a_42982_21320.t1 65.941
R10914 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t10 142.458
R10915 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t7 142.458
R10916 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t21 141.674
R10917 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t16 141.674
R10918 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t13 140.891
R10919 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t4 140.891
R10920 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t28 139.879
R10921 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t19 139.879
R10922 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t26 139.879
R10923 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t23 139.879
R10924 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t25 139.879
R10925 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t17 139.879
R10926 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t31 139.879
R10927 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t29 139.879
R10928 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t24 139.879
R10929 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t18 139.879
R10930 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t27 135.441
R10931 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t22 135.441
R10932 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t30 135.435
R10933 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t20 135.435
R10934 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t6 134.732
R10935 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t5 134.732
R10936 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t1 134.732
R10937 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t3 134.732
R10938 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t8 134.732
R10939 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t0 134.732
R10940 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t9 134.732
R10941 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n29 134.732
R10942 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t12 134.712
R10943 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t2 134.712
R10944 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t14 134.712
R10945 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t11 134.712
R10946 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n20 5.61925
R10947 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n5 4.9505
R10948 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n2 4.57291
R10949 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n23 4.57291
R10950 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n19 4.5005
R10951 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n21 4.5005
R10952 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n0 4.5005
R10953 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n28 4.5005
R10954 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n3 4.05258
R10955 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n26 4.02292
R10956 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n27 3.78175
R10957 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n10 3.67541
R10958 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n11 3.5885
R10959 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n6 3.5885
R10960 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n17 3.4105
R10961 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n25 3.4105
R10962 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n14 3.38383
R10963 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n22 3.13383
R10964 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n1 3.13383
R10965 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n16 3.113
R10966 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n24 2.21508
R10967 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n12 1.79633
R10968 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n7 1.79633
R10969 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n18 1.56717
R10970 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n9 1.54633
R10971 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n13 1.338
R10972 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n15 1.338
R10973 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n4 1.338
R10974 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n8 1.338
R10975 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t0 227.856
R10976 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n2 152.333
R10977 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t4 140.382
R10978 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t3 114.031
R10979 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t1 83.3993
R10980 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t2 81.5883
R10981 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n3 14.4422
R10982 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n1 7.56882
R10983 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n0 5.08175
R10984 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R10985 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n1 863.124
R10986 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n0 585
R10987 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t0 495.469
R10988 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t6 216.893
R10989 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t4 216.893
R10990 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t5 215.142
R10991 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t2 213.042
R10992 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t9 212.393
R10993 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t8 208.054
R10994 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n10 152
R10995 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t1 141.189
R10996 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t0 140.738
R10997 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t3 114.031
R10998 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t7 81.5883
R10999 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n7 32.6672
R11000 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n9 25.5255
R11001 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 16.7132
R11002 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 13.7979
R11003 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 13.1884
R11004 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 11.6369
R11005 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n8 11.0276
R11006 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n6 11.0088
R11007 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 10.1408
R11008 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 8.97342
R11009 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n3 7.94225
R11010 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 6.14988
R11011 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n5 5.16396
R11012 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 4.67598
R11013 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n4 4.23576
R11014 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 2.16154
R11015 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 2.16154
R11016 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n11 1.16414
R11017 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n2 0.665435
R11018 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n12 0.582318
R11019 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.166365
R11020 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t26 85.4005
R11021 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t21 84.4381
R11022 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t14 84.4381
R11023 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t17 84.4381
R11024 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t16 84.4381
R11025 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t12 84.4381
R11026 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t20 84.4381
R11027 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t1 84.4381
R11028 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t25 84.4381
R11029 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t3 84.4381
R11030 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n4 75.1793
R11031 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n3 75.1793
R11032 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n2 75.1793
R11033 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n0 75.1793
R11034 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n42 75.1793
R11035 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t8 65.5634
R11036 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t9 65.0567
R11037 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n26 59.2318
R11038 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n24 49.0864
R11039 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n25 49.0864
R11040 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n23 24.3828
R11041 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n32 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n31 19.7755
R11042 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n28 18.0943
R11043 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n34 10.5047
R11044 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n38 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n37 10.5047
R11045 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n41 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n40 10.5047
R11046 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n45 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n44 10.5047
R11047 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t6 10.3318
R11048 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t5 10.3318
R11049 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t22 10.3318
R11050 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t23 10.3318
R11051 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t10 10.3318
R11052 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t4 10.3318
R11053 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n33 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 10.0234
R11054 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n36 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 10.0234
R11055 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n39 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 10.0234
R11056 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 10.0234
R11057 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n1 10.0214
R11058 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t15 9.23217
R11059 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t18 9.23217
R11060 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t11 9.23217
R11061 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t13 9.23217
R11062 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t7 9.23217
R11063 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t19 9.23217
R11064 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t27 9.23217
R11065 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t24 9.23217
R11066 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t0 9.23217
R11067 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n42 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t2 9.23217
R11068 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 5.863
R11069 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n29 5.72967
R11070 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n31 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n30 5.20675
R11071 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n7 3.90596
R11072 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n22 3.4105
R11073 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n18 3.4105
R11074 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n14 3.4105
R11075 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n10 3.4105
R11076 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n33 0.962993
R11077 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n37 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n36 0.962993
R11078 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n40 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n39 0.962993
R11079 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n44 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n43 0.962974
R11080 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n27 0.955189
R11081 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t37 0.523604
R11082 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t36 0.523604
R11083 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t40 0.523604
R11084 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t38 0.523604
R11085 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t33 0.523604
R11086 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t31 0.523604
R11087 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t30 0.523604
R11088 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t28 0.523604
R11089 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t47 0.523604
R11090 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t46 0.523604
R11091 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n11 0.495958
R11092 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n15 0.495958
R11093 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n19 0.495958
R11094 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t43 0.28175
R11095 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t29 0.28175
R11096 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t45 0.28175
R11097 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t32 0.28175
R11098 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t39 0.28175
R11099 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t44 0.28175
R11100 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t35 0.28175
R11101 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t42 0.28175
R11102 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t34 0.28175
R11103 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t41 0.28175
R11104 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n32 0.188
R11105 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n35 0.188
R11106 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n38 0.188
R11107 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n41 0.188
R11108 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n45 0.188
R11109 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n5 0.121427
R11110 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n6 0.121427
R11111 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n8 0.121427
R11112 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n9 0.121427
R11113 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n12 0.121427
R11114 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n13 0.121427
R11115 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n16 0.121427
R11116 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n17 0.121427
R11117 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n20 0.121427
R11118 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n21 0.121427
R11119 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t6 118.626
R11120 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t8 118.626
R11121 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t7 118.005
R11122 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t9 118.005
R11123 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t4 70.0103
R11124 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t3 69.7645
R11125 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t1 69.6506
R11126 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t0 59.4447
R11127 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t2 50.8563
R11128 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t5 49.6789
R11129 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n0 16.5734
R11130 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n1 11.3963
R11131 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n6 9.83175
R11132 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n3 2.93383
R11133 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n2 2.42967
R11134 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n7 2.11508
R11135 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n4 0.629667
R11136 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n5 0.629667
R11137 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t7 739.265
R11138 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t12 230.155
R11139 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t6 229.369
R11140 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t4 212.081
R11141 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t10 212.081
R11142 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 203.923
R11143 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 186.001
R11144 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 157.927
R11145 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t9 157.856
R11146 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t11 157.07
R11147 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 152
R11148 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t8 139.78
R11149 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t5 139.78
R11150 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 101.49
R11151 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 61.346
R11152 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t1 26.5955
R11153 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t2 26.5955
R11154 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t3 24.9236
R11155 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t0 24.9236
R11156 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 19.6746
R11157 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 19.6318
R11158 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.B 14.4147
R11159 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 13.5685
R11160 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[1] 11.5193
R11161 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 10.7525
R11162 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 9.64425
R11163 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 9.30224
R11164 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y 6.6565
R11165 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y 5.04292
R11166 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y 3.8405
R11167 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.A 3.0725
R11168 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y 2.5605
R11169 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.A 2.13383
R11170 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 1.93989
R11171 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t3 228.496
R11172 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t2 228.496
R11173 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t1 227.538
R11174 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t0 227.538
R11175 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t4 221.974
R11176 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t5 221.974
R11177 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t7 221.851
R11178 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t6 221.851
R11179 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n4 9.92404
R11180 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n3 9.90278
R11181 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n0 6.28466
R11182 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n1 4.10425
R11183 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n2 0.404985
R11184 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n5 0.299591
R11185 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59.t1 248.95
R11186 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59.t2 10.6701
R11187 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59.t0 10.5739
R11188 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59.n0 2.77016
R11189 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60.t1 249.148
R11190 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60.t0 10.6257
R11191 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60.t2 10.5285
R11192 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60.n0 2.09277
R11193 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n1 863.124
R11194 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n0 585
R11195 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t0 495.469
R11196 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t8 217.555
R11197 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t10 216.893
R11198 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t3 216.893
R11199 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t2 216.893
R11200 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t9 216.893
R11201 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t4 216.893
R11202 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t7 216.893
R11203 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t11 216.893
R11204 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t5 216.893
R11205 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n13 152
R11206 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t1 141.189
R11207 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t0 140.738
R11208 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t12 114.031
R11209 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t6 81.5883
R11210 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n12 73.9371
R11211 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 16.7132
R11212 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 13.7979
R11213 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 13.1884
R11214 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 11.6369
R11215 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 10.1408
R11216 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n3 7.94225
R11217 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 6.14988
R11218 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 2.16154
R11219 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 2.16154
R11220 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n14 1.16414
R11221 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n2 0.665435
R11222 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n9 0.663962
R11223 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n8 0.663962
R11224 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n7 0.663962
R11225 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n6 0.663962
R11226 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n5 0.663962
R11227 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n4 0.663962
R11228 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n10 0.658467
R11229 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n15 0.582318
R11230 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.155033
R11231 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n11 0.0138929
R11232 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.n0 679.191
R11233 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.t1 10.7575
R11234 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.t2 10.7275
R11235 a_15224_18696.n0 a_15224_18696.t2 671.891
R11236 a_15224_18696.n0 a_15224_18696.t1 666.433
R11237 a_15224_18696.t0 a_15224_18696.n0 666.404
R11238 DIN1.n1 DIN1.t0 212.081
R11239 DIN1.n0 DIN1.t3 212.081
R11240 DIN1.n2 DIN1.n1 183.185
R11241 DIN1.n1 DIN1.t2 139.78
R11242 DIN1.n0 DIN1.t1 139.78
R11243 DIN1.n1 DIN1.n0 61.346
R11244 DIN1 DIN1.n2 14.2776
R11245 DIN1.n2 DIN1 5.8885
R11246 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t4 757.36
R11247 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t6 212.081
R11248 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t5 212.081
R11249 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 203.923
R11250 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 186.001
R11251 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t8 139.78
R11252 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t7 139.78
R11253 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 101.49
R11254 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 61.346
R11255 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t2 26.5955
R11256 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t3 26.5955
R11257 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t1 24.9236
R11258 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t0 24.9236
R11259 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 13.5685
R11260 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 10.7525
R11261 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 9.64425
R11262 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 9.30224
R11263 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y 6.6565
R11264 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y 5.04292
R11265 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y 3.8405
R11266 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.A 3.0725
R11267 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y 2.5605
R11268 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 1.93989
R11269 a_44234_11946.t0 a_44234_11946.t1 114.052
R11270 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t1 675.533
R11271 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t2 10.7601
R11272 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t0 10.7161
R11273 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.n0 2.73056
R11274 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t1 676.553
R11275 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t2 10.7798
R11276 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t0 10.6302
R11277 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.n0 3.43637
R11278 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n1 863.124
R11279 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n0 585
R11280 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t0 495.469
R11281 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t14 217.555
R11282 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t12 217.555
R11283 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t6 217.555
R11284 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t10 216.893
R11285 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t16 216.893
R11286 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t15 216.893
R11287 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t11 216.893
R11288 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t5 216.893
R11289 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t7 216.893
R11290 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t4 216.893
R11291 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t2 216.893
R11292 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t17 216.893
R11293 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t13 216.893
R11294 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t3 216.893
R11295 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t9 216.893
R11296 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t8 216.893
R11297 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t1 141.189
R11298 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t0 140.738
R11299 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n18 65.2685
R11300 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 14.7463
R11301 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 11.6369
R11302 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 10.1408
R11303 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n3 7.94225
R11304 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n19 7.75808
R11305 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 6.59444
R11306 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n17 6.48592
R11307 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 6.37342
R11308 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 6.14988
R11309 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 2.16154
R11310 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n2 0.665435
R11311 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n15 0.663962
R11312 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n14 0.663962
R11313 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n11 0.663962
R11314 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n12 0.663962
R11315 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n4 0.663962
R11316 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n5 0.663962
R11317 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n6 0.663962
R11318 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n7 0.663962
R11319 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n8 0.663962
R11320 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n9 0.663962
R11321 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n16 0.320692
R11322 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n13 0.320692
R11323 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n10 0.274859
R11324 a_15629_7686.n0 a_15629_7686.t2 671.846
R11325 a_15629_7686.n2 a_15629_7686.t4 667.794
R11326 a_15629_7686.t0 a_15629_7686.n2 667.572
R11327 a_15629_7686.n0 a_15629_7686.t1 665.36
R11328 a_15629_7686.n1 a_15629_7686.t3 665.36
R11329 a_15629_7686.n1 a_15629_7686.n0 6.63383
R11330 a_15629_7686.n2 a_15629_7686.n1 4.51925
R11331 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t2 675.929
R11332 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t1 10.7912
R11333 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t0 10.6717
R11334 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.n0 4.09783
R11335 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30.t1 249.358
R11336 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30.t2 10.5296
R11337 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30.t0 10.5295
R11338 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30.n0 0.905521
R11339 a_31594_7686.n2 a_31594_7686.t3 246.978
R11340 a_31594_7686.n0 a_31594_7686.t1 244.013
R11341 a_31594_7686.n0 a_31594_7686.t2 240.072
R11342 a_31594_7686.n1 a_31594_7686.t4 239.692
R11343 a_31594_7686.t0 a_31594_7686.n2 239.692
R11344 a_31594_7686.n2 a_31594_7686.n1 6.788
R11345 a_31594_7686.n1 a_31594_7686.n0 2.26092
R11346 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46.n0 238.37
R11347 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46.t2 10.7799
R11348 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46.t1 10.7013
R11349 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47.n0 237.56
R11350 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47.t1 10.5728
R11351 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47.t2 10.5285
R11352 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t5 230.155
R11353 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t13 230.155
R11354 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t7 229.369
R11355 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t12 212.081
R11356 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t11 212.081
R11357 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n16 203.922
R11358 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n3 186.001
R11359 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n8 157.927
R11360 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t6 157.856
R11361 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t4 157.856
R11362 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t10 157.07
R11363 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n5 153.338
R11364 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n9 152
R11365 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t9 139.78
R11366 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t8 139.78
R11367 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n0 101.49
R11368 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n2 61.346
R11369 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n11 31.3499
R11370 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n12 29.8627
R11371 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t0 26.5955
R11372 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t2 26.5955
R11373 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t3 24.9236
R11374 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t1 24.9236
R11375 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n6 17.8391
R11376 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 13.5685
R11377 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 11.0938
R11378 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 10.7525
R11379 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n10 9.9845
R11380 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n13 9.64425
R11381 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n4 9.30224
R11382 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 6.6565
R11383 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n15 5.04292
R11384 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n14 3.8405
R11385 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 3.0725
R11386 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 3.05722
R11387 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n1 2.5605
R11388 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 2.3045
R11389 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n7 2.24073
R11390 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 1.93989
R11391 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.600109
R11392 a_44255_3438.t0 a_44255_3438.t1 49.8467
R11393 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t0 272.038
R11394 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t0 258.846
R11395 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t3 241.536
R11396 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n0 224.776
R11397 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t4 169.237
R11398 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n2 153.032
R11399 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n3 32.3107
R11400 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t1 26.5955
R11401 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t2 26.5955
R11402 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 24.8072
R11403 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 3.76521
R11404 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n5 2.30266
R11405 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n4 1.65805
R11406 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n1 1.38179
R11407 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.921363
R11408 a_44479_3254.t0 a_44479_3254.t1 49.8467
R11409 a_44234_10322.t0 a_44234_10322.t1 114.052
R11410 a_43698_9766.t0 a_43698_9766.n0 228.04
R11411 a_43698_9766.n0 a_43698_9766.t2 145.648
R11412 a_43698_9766.n0 a_43698_9766.t1 83.2159
R11413 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n1 863.124
R11414 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n0 585
R11415 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t0 495.469
R11416 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t4 217.555
R11417 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t6 216.893
R11418 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t5 216.893
R11419 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t2 216.893
R11420 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t3 212.393
R11421 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t1 141.189
R11422 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t0 140.738
R11423 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n8 90.6776
R11424 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 14.3755
R11425 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 11.6369
R11426 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 10.1408
R11427 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n9 8.53383
R11428 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n3 7.94225
R11429 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 6.14988
R11430 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 5.81868
R11431 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n7 4.5005
R11432 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 2.16154
R11433 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n2 0.665435
R11434 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n4 0.663962
R11435 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n5 0.663962
R11436 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n6 0.663962
R11437 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.325019
R11438 a_17148_18696.t0 a_17148_18696.n0 670.792
R11439 a_17148_18696.n0 a_17148_18696.t2 666.963
R11440 a_17148_18696.n0 a_17148_18696.t1 665.304
R11441 a_14514_18696.t0 a_14514_18696.n0 671.227
R11442 a_14514_18696.n0 a_14514_18696.t1 665.75
R11443 a_14514_18696.n0 a_14514_18696.t2 665.298
R11444 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14.n0 678.111
R11445 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14.t2 10.7803
R11446 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14.t1 10.7023
R11447 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15.t1 666.722
R11448 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15.n0 10.6331
R11449 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15.t2 10.5285
R11450 DIN5.n1 DIN5.t3 212.081
R11451 DIN5.n0 DIN5.t2 212.081
R11452 DIN5.n2 DIN5.n1 183.185
R11453 DIN5.n1 DIN5.t1 139.78
R11454 DIN5.n0 DIN5.t0 139.78
R11455 DIN5.n1 DIN5.n0 61.346
R11456 DIN5 DIN5.n2 14.2776
R11457 DIN5.n2 DIN5 5.8885
R11458 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.n0 679.261
R11459 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.t2 10.7728
R11460 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.t1 10.7357
R11461 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.n0 677.365
R11462 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.t1 10.79
R11463 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.t2 10.6292
R11464 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t15 140.945
R11465 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t11 140.945
R11466 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t12 140.945
R11467 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t13 140.945
R11468 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t14 139.635
R11469 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t9 139.635
R11470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t10 139.625
R11471 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t8 139.625
R11472 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t1 134.712
R11473 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t3 134.712
R11474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t6 134.712
R11475 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t4 134.712
R11476 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t2 134.712
R11477 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t0 134.712
R11478 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t5 134.712
R11479 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n13 134.712
R11480 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n0 11.8254
R11481 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n9 10.2587
R11482 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n8 9.9879
R11483 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n12 8.42123
R11484 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n5 6.5255
R11485 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n2 4.95883
R11486 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n1 4.688
R11487 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n3 4.42741
R11488 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n11 4.14826
R11489 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n6 3.4105
R11490 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n10 3.4105
R11491 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n4 3.12133
R11492 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n7 1.1285
R11493 a_38672_20477.n0 a_38672_20477.t2 233.361
R11494 a_38672_20477.t1 a_38672_20477.n0 229.339
R11495 a_38672_20477.n0 a_38672_20477.t0 227.399
R11496 a_21375_20174.n0 a_21375_20174.t2 251.903
R11497 a_21375_20174.t0 a_21375_20174.n1 248.659
R11498 a_21375_20174.n0 a_21375_20174.t3 241.815
R11499 a_21375_20174.n1 a_21375_20174.t1 238.732
R11500 a_21375_20174.n1 a_21375_20174.n0 3.24425
R11501 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.t3 237.774
R11502 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.t2 237.685
R11503 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.t1 10.6569
R11504 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.n1 10.6569
R11505 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16.n0 3.39554
R11506 DIN8.n1 DIN8.t3 212.081
R11507 DIN8.n0 DIN8.t2 212.081
R11508 DIN8.n2 DIN8.n1 183.185
R11509 DIN8.n1 DIN8.t1 139.78
R11510 DIN8.n0 DIN8.t0 139.78
R11511 DIN8.n1 DIN8.n0 61.346
R11512 DIN8 DIN8.n2 14.2776
R11513 DIN8.n2 DIN8 5.8885
R11514 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t2 676.497
R11515 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t1 10.7163
R11516 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t0 10.676
R11517 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.n0 2.06176
R11518 a_16615_7686.n1 a_16615_7686.t2 672.396
R11519 a_16615_7686.n0 a_16615_7686.t4 669.848
R11520 a_16615_7686.n0 a_16615_7686.t1 666.222
R11521 a_16615_7686.n1 a_16615_7686.t3 665.909
R11522 a_16615_7686.t0 a_16615_7686.n2 665.909
R11523 a_16615_7686.n2 a_16615_7686.n1 6.63383
R11524 a_16615_7686.n2 a_16615_7686.n0 3.01508
R11525 a_43724_15866.t0 a_43724_15866.t1 55.3905
R11526 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t1 230.518
R11527 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t3 229.369
R11528 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t4 229.369
R11529 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t0 157.62
R11530 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t5 157.07
R11531 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t2 157.07
R11532 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n0 152.712
R11533 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n2 152.475
R11534 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 24.2121
R11535 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n5 23.559
R11536 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n7 11.6875
R11537 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n1 10.2234
R11538 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n3 9.77342
R11539 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 7.23528
R11540 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 5.45235
R11541 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 5.21532
R11542 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 5.04292
R11543 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n6 4.73093
R11544 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n4 4.6005
R11545 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.31925
R11546 a_45023_21136.t0 a_45023_21136.t1 49.8467
R11547 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n1 863.124
R11548 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n0 585
R11549 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t0 495.469
R11550 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t11 219.499
R11551 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t12 217.555
R11552 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t15 217.555
R11553 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t17 216.893
R11554 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t13 216.893
R11555 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t19 216.893
R11556 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t18 216.893
R11557 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t5 216.893
R11558 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t9 216.893
R11559 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t6 213.218
R11560 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t4 213.218
R11561 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t22 212.554
R11562 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t7 212.554
R11563 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t3 212.554
R11564 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t20 212.554
R11565 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t16 212.554
R11566 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t8 212.393
R11567 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t14 212.393
R11568 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t2 208.054
R11569 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n24 152
R11570 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t1 141.189
R11571 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t0 140.738
R11572 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t21 114.031
R11573 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t10 81.5883
R11574 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n23 29.1651
R11575 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n15 18.9547
R11576 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 16.7132
R11577 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n5 14.8692
R11578 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n22 14.013
R11579 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n14 13.9942
R11580 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 13.7979
R11581 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 13.1884
R11582 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 11.6369
R11583 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 10.1408
R11584 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 10.0338
R11585 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n6 8.81508
R11586 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n3 7.94225
R11587 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 6.14988
R11588 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n4 4.5005
R11589 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n13 4.5005
R11590 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n21 4.5005
R11591 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 2.16154
R11592 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 2.16154
R11593 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n25 1.16414
R11594 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n2 0.665435
R11595 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n7 0.663962
R11596 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n8 0.663962
R11597 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n12 0.663962
R11598 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n11 0.663962
R11599 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n10 0.663962
R11600 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n9 0.663962
R11601 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n16 0.663962
R11602 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n18 0.663962
R11603 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n19 0.663962
R11604 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n20 0.663962
R11605 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n26 0.582318
R11606 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.541365
R11607 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.310596
R11608 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.293769
R11609 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n17 0.123096
R11610 a_27620_6250.n2 a_27620_6250.t2 247.553
R11611 a_27620_6250.n0 a_27620_6250.t1 245.569
R11612 a_27620_6250.n1 a_27620_6250.t3 244.964
R11613 a_27620_6250.n0 a_27620_6250.t4 238.899
R11614 a_27620_6250.t0 a_27620_6250.n2 238.899
R11615 a_27620_6250.n1 a_27620_6250.n0 5.463
R11616 a_27620_6250.n2 a_27620_6250.n1 1.55883
R11617 a_33634_8950.n0 a_33634_8950.t2 244.725
R11618 a_33634_8950.n0 a_33634_8950.t1 242.994
R11619 a_33634_8950.t0 a_33634_8950.n0 239.673
R11620 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27.t0 248.95
R11621 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27.t2 10.6701
R11622 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27.t1 10.5739
R11623 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27.n0 2.76539
R11624 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t0 230.71
R11625 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t6 230.576
R11626 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t9 230.155
R11627 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t5 230.155
R11628 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n7 205.28
R11629 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t4 158.275
R11630 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t7 157.856
R11631 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t8 157.856
R11632 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n8 153.067
R11633 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n2 152
R11634 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n0 152
R11635 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t2 135.947
R11636 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n11 67.4857
R11637 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n10 44.0818
R11638 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n6 33.5064
R11639 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t3 26.5955
R11640 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t1 26.5955
R11641 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n5 23.9017
R11642 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n9 19.3316
R11643 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 16.4149
R11644 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n1 12.2559
R11645 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n3 11.0199
R11646 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 5.6005
R11647 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n4 5.0505
R11648 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 2.10199
R11649 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 2.10199
R11650 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.05675
R11651 a_24687_20174.n0 a_24687_20174.t2 249.886
R11652 a_24687_20174.t0 a_24687_20174.n1 247.333
R11653 a_24687_20174.n1 a_24687_20174.t1 240.75
R11654 a_24687_20174.n0 a_24687_20174.t3 239.798
R11655 a_24687_20174.n1 a_24687_20174.n0 2.55258
R11656 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t0 675.929
R11657 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t2 10.8219
R11658 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t1 10.6741
R11659 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.n0 4.11026
R11660 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t0 676.321
R11661 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t2 13.4699
R11662 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t1 10.7776
R11663 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.n0 4.72836
R11664 a_43391_3794.t0 a_43391_3794.t1 49.8467
R11665 a_43391_3878.t0 a_43391_3878.t1 60.9236
R11666 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n1 863.124
R11667 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n0 585
R11668 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t0 495.469
R11669 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t3 223.035
R11670 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t4 216.893
R11671 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t5 215.142
R11672 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t7 208.054
R11673 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n8 152
R11674 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t1 141.189
R11675 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t0 140.738
R11676 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t2 114.031
R11677 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t6 81.5883
R11678 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n5 32.088
R11679 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n7 29.0609
R11680 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUTB 16.7132
R11681 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.A 13.7979
R11682 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 13.1884
R11683 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 11.6369
R11684 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n6 10.6609
R11685 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 10.1408
R11686 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n3 7.94225
R11687 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n5 top_DAC_0/top_final_switch_0.bb[0] 7.39217
R11688 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 6.14988
R11689 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.bb[0] 4.5606
R11690 top_DAC_0/top_final_switch_0.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n4 4.25242
R11691 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 2.16154
R11692 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 2.16154
R11693 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n9 1.16414
R11694 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n2 0.665435
R11695 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n10 0.582318
R11696 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUTB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.bb[0] 0.185917
R11697 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t1 672.309
R11698 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t2 10.7751
R11699 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t0 10.6965
R11700 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.n0 1.35813
R11701 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t0 672.795
R11702 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t1 10.7151
R11703 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t2 10.6674
R11704 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.n0 2.05222
R11705 a_8506_12595.n4 a_8506_12595.t4 221.916
R11706 a_8506_12595.n3 a_8506_12595.t2 221.913
R11707 a_8506_12595.n3 a_8506_12595.t5 221.91
R11708 a_8506_12595.n4 a_8506_12595.t3 221.909
R11709 a_8506_12595.n8 a_8506_12595.n7 71.3963
R11710 a_8506_12595.n2 a_8506_12595.n1 71.3963
R11711 a_8506_12595.n2 a_8506_12595.n0 71.3963
R11712 a_8506_12595.n9 a_8506_12595.n8 71.3963
R11713 a_8506_12595.n7 a_8506_12595.t9 16.5305
R11714 a_8506_12595.n7 a_8506_12595.t7 16.5305
R11715 a_8506_12595.n1 a_8506_12595.t11 16.5305
R11716 a_8506_12595.n1 a_8506_12595.t1 16.5305
R11717 a_8506_12595.n0 a_8506_12595.t6 16.5305
R11718 a_8506_12595.n0 a_8506_12595.t8 16.5305
R11719 a_8506_12595.t0 a_8506_12595.n9 16.5305
R11720 a_8506_12595.n9 a_8506_12595.t10 16.5305
R11721 a_8506_12595.n5 a_8506_12595.n4 9.24407
R11722 a_8506_12595.n5 a_8506_12595.n3 7.48275
R11723 a_8506_12595.n6 a_8506_12595.n5 4.33483
R11724 a_8506_12595.n6 a_8506_12595.n2 0.3505
R11725 a_8506_12595.n8 a_8506_12595.n6 0.3505
R11726 a_34304_8950.n0 a_34304_8950.t2 245.95
R11727 a_34304_8950.n0 a_34304_8950.t1 243.918
R11728 a_34304_8950.t0 a_34304_8950.n0 239.124
R11729 a_28606_6250.n2 a_28606_6250.t2 248.102
R11730 a_28606_6250.n0 a_28606_6250.t1 246.119
R11731 a_28606_6250.n1 a_28606_6250.t3 245.203
R11732 a_28606_6250.n0 a_28606_6250.t4 239.45
R11733 a_28606_6250.t0 a_28606_6250.n2 239.45
R11734 a_28606_6250.n2 a_28606_6250.n1 6.32758
R11735 a_28606_6250.n1 a_28606_6250.n0 0.69425
R11736 a_5111_10963.n1 a_5111_10963.t0 133.338
R11737 a_5111_10963.n2 a_5111_10963.t2 133.338
R11738 a_5111_10963.n1 a_5111_10963.n0 48.5755
R11739 a_5111_10963.n3 a_5111_10963.n2 48.5755
R11740 a_5111_10963.n0 a_5111_10963.t1 10.3318
R11741 a_5111_10963.n0 a_5111_10963.t4 10.3318
R11742 a_5111_10963.n3 a_5111_10963.t5 10.3318
R11743 a_5111_10963.t3 a_5111_10963.n3 10.3318
R11744 a_5111_10963.n2 a_5111_10963.n1 10.0148
R11745 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t4 147.899
R11746 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t5 146.752
R11747 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n2 79.7972
R11748 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n1 79.7972
R11749 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n3 79.7972
R11750 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n0 79.6389
R11751 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t7 9.23217
R11752 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t0 9.23217
R11753 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t8 9.23217
R11754 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t1 9.23217
R11755 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t2 9.23217
R11756 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t9 9.23217
R11757 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t3 9.23217
R11758 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t6 9.23217
R11759 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n5 4.68805
R11760 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n6 0.429667
R11761 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n4 0.429667
R11762 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n7 0.158833
R11763 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t26 94.4233
R11764 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t25 84.4574
R11765 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t16 84.4574
R11766 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t14 84.4574
R11767 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t20 84.4574
R11768 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t10 84.4574
R11769 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t18 84.4381
R11770 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t13 84.4381
R11771 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t21 84.4381
R11772 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t11 84.4381
R11773 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n4 75.1793
R11774 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n3 75.1793
R11775 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n2 75.1793
R11776 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n1 75.1793
R11777 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n0 75.1793
R11778 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t5 65.725
R11779 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t4 65.2617
R11780 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n26 50.072
R11781 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n25 49.0864
R11782 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n28 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n27 49.0864
R11783 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n23 24.7318
R11784 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n29 17.6109
R11785 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n7 10.5047
R11786 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n11 10.5047
R11787 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n15 10.5047
R11788 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n19 10.5047
R11789 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t2 10.3318
R11790 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n25 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t6 10.3318
R11791 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t3 10.3318
R11792 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n26 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t7 10.3318
R11793 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t0 10.3318
R11794 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n27 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t1 10.3318
R11795 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n28 9.98768
R11796 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n8 9.98569
R11797 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n12 9.98569
R11798 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n16 9.98569
R11799 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n20 9.98569
R11800 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t27 9.23217
R11801 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t24 9.23217
R11802 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t15 9.23217
R11803 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t17 9.23217
R11804 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t12 9.23217
R11805 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t23 9.23217
R11806 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t19 9.23217
R11807 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t22 9.23217
R11808 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t9 9.23217
R11809 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t8 9.23217
R11810 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n30 5.913
R11811 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n24 5.67967
R11812 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n21 0.773962
R11813 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n5 0.757842
R11814 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n9 0.757842
R11815 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n13 0.757842
R11816 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n17 0.757842
R11817 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n6 0.306265
R11818 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n10 0.306265
R11819 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n14 0.306265
R11820 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n18 0.306265
R11821 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n23 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n22 0.30484
R11822 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n22 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.0174229
R11823 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.016045
R11824 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.016045
R11825 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.016045
R11826 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.016045
R11827 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t10 134.734
R11828 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t7 134.734
R11829 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t11 134.734
R11830 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t9 134.734
R11831 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t6 134.734
R11832 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t5 134.734
R11833 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t4 134.734
R11834 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t8 134.734
R11835 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n12 79.7972
R11836 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n2 79.7972
R11837 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n1 79.7972
R11838 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n0 79.6389
R11839 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t14 9.23217
R11840 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t1 9.23217
R11841 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t2 9.23217
R11842 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t13 9.23217
R11843 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t15 9.23217
R11844 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t0 9.23217
R11845 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t3 9.23217
R11846 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t12 9.23217
R11847 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n4 9.2005
R11848 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n7 9.2005
R11849 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n6 6.63891
R11850 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n10 5.06405
R11851 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n5 4.5005
R11852 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n8 4.5005
R11853 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n9 4.43133
R11854 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n11 0.429667
R11855 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n3 0.429667
R11856 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n13 0.158833
R11857 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t1 227.707
R11858 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t5 227.707
R11859 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t7 227.707
R11860 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t2 227.707
R11861 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t6 226.386
R11862 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t3 226.386
R11863 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t4 226.386
R11864 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t0 226.386
R11865 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t11 221.911
R11866 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t14 221.911
R11867 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t8 221.911
R11868 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t13 221.911
R11869 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t15 221.911
R11870 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t12 221.911
R11871 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t9 221.911
R11872 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t10 221.911
R11873 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n8 9.59425
R11874 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n10 8.80675
R11875 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n11 8.02758
R11876 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n7 7.24008
R11877 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n4 4.43383
R11878 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n2 4.17674
R11879 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n9 3.92608
R11880 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n0 3.64633
R11881 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n12 3.4105
R11882 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n5 3.4105
R11883 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n1 2.86717
R11884 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n3 2.07967
R11885 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n6 0.718318
R11886 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n13 0.424924
R11887 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12.t1 239.088
R11888 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12.n0 10.5771
R11889 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12.t2 10.5739
R11890 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13.t2 238.671
R11891 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13.t1 10.5309
R11892 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13.n0 10.5295
R11893 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33.t2 236.65
R11894 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33.t1 10.6732
R11895 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33.n0 10.5739
R11896 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34.t1 246.804
R11897 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34.t0 10.6257
R11898 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34.t2 10.5285
R11899 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34.n0 0.86158
R11900 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t3 221.851
R11901 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t1 221.851
R11902 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t4 140.061
R11903 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t5 139.566
R11904 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t15 120.969
R11905 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t11 120.969
R11906 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t6 120.969
R11907 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t9 120.969
R11908 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t12 120.969
R11909 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t14 120.969
R11910 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t17 120.969
R11911 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t8 120.969
R11912 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t7 120.969
R11913 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t13 120.969
R11914 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t10 120.969
R11915 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t16 120.969
R11916 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t2 108.365
R11917 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t0 108.365
R11918 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n0 15.3463
R11919 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n15 13.5257
R11920 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n20 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n19 8.1267
R11921 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n17 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n16 5.84703
R11922 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n1 4.95104
R11923 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n19 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n18 4.79425
R11924 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n20 1.21717
R11925 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n3 0.713
R11926 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n4 0.713
R11927 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n5 0.713
R11928 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n13 0.713
R11929 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n12 0.713
R11930 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n11 0.713
R11931 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n9 0.713
R11932 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n8 0.713
R11933 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n7 0.713
R11934 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n10 0.690083
R11935 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.598417
R11936 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n0 0.557293
R11937 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n17 0.546515
R11938 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.523417
R11939 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n15 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n14 0.167167
R11940 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n6 0.140083
R11941 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.140083
R11942 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.140083
R11943 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n21 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.08175
R11944 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n21 0.063
R11945 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.0525833
R11946 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n16 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n2 0.0143889
R11947 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n10 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t3 221.913
R11948 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t0 221.913
R11949 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n10 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t4 221.911
R11950 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t2 221.911
R11951 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n12 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t6 221.851
R11952 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n8 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t5 221.851
R11953 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t1 221.851
R11954 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n13 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t7 221.851
R11955 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t12 214.787
R11956 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t13 214.787
R11957 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t14 214.005
R11958 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t15 214.005
R11959 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t10 212.323
R11960 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t8 212.042
R11961 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t11 48.2714
R11962 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n17 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t9 48.2714
R11963 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n2 17.7367
R11964 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n5 9.98379
R11965 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n11 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n10 9.98379
R11966 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n16 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n15 9.65976
R11967 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n15 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n9 8.23783
R11968 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n0 7.77967
R11969 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n1 7.65675
R11970 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n15 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n14 5.65425
R11971 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n14 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n13 4.73193
R11972 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n9 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n8 4.73193
R11973 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n6 4.73193
R11974 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n12 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n11 4.73193
R11975 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n16 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n4 2.42885
R11976 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n17 1.47876
R11977 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n17 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n16 1.40802
R11978 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n3 1.09089
R11979 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n9 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n6 0.246333
R11980 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n14 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n11 0.246333
R11981 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n8 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n7 0.123417
R11982 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n13 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n12 0.123417
R11983 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 0.0734167
R11984 a_23859_20174.n0 a_23859_20174.t1 248.969
R11985 a_23859_20174.n1 a_23859_20174.t2 246.287
R11986 a_23859_20174.t0 a_23859_20174.n1 241.666
R11987 a_23859_20174.n0 a_23859_20174.t3 238.881
R11988 a_23859_20174.n1 a_23859_20174.n0 2.68175
R11989 top_DAC_0/top_final_switch_0.VOUT[2].n2 top_DAC_0/top_final_switch_0.VOUT[2].n0 603.66
R11990 top_DAC_0/top_final_switch_0.VOUT[2].n2 top_DAC_0/top_final_switch_0.VOUT[2].n1 202.21
R11991 top_DAC_0/top_final_switch_0.VOUT[2].n3 top_DAC_0/top_final_switch_0.VOUT[2].t8 172.237
R11992 top_DAC_0/top_final_switch_0.VOUT[2].n4 top_DAC_0/top_final_switch_0.VOUT[2].t6 171.161
R11993 top_DAC_0/top_final_switch_0.VOUT[2].n3 top_DAC_0/top_final_switch_0.VOUT[2].t9 170.625
R11994 top_DAC_0/top_final_switch_0.VOUT[2].n4 top_DAC_0/top_final_switch_0.VOUT[2].t11 170.625
R11995 top_DAC_0/top_final_switch_0.VOUT[2].n7 top_DAC_0/top_final_switch_0.VOUT[2].t5 121.868
R11996 top_DAC_0/top_final_switch_0.VOUT[2].n6 top_DAC_0/top_final_switch_0.VOUT[2].t4 120.793
R11997 top_DAC_0/top_final_switch_0.VOUT[2].n7 top_DAC_0/top_final_switch_0.VOUT[2].t7 120.255
R11998 top_DAC_0/top_final_switch_0.VOUT[2].n6 top_DAC_0/top_final_switch_0.VOUT[2].t10 120.255
R11999 top_DAC_0/top_final_switch_0.VOUT[2].n0 top_DAC_0/top_final_switch_0.VOUT[2].t3 65.941
R12000 top_DAC_0/top_final_switch_0.VOUT[2].n0 top_DAC_0/top_final_switch_0.VOUT[2].t2 65.941
R12001 top_DAC_0/top_final_switch_0.VOUT[2].n1 top_DAC_0/top_final_switch_0.VOUT[2].t0 39.3576
R12002 top_DAC_0/top_final_switch_0.VOUT[2].n1 top_DAC_0/top_final_switch_0.VOUT[2].t1 39.3576
R12003 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_final_switch_0.VOUT[2].n9 11.638
R12004 top_DAC_0/top_final_switch_0.VOUT[2].n5 top_DAC_0/top_final_switch_0.VOUT[2].n3 8.69842
R12005 top_DAC_0/top_final_switch_0.VOUT[2].n8 top_DAC_0/top_final_switch_0.VOUT[2].n6 7.53592
R12006 top_DAC_0/top_final_switch_0.VOUT[2].n10 top_DAC_0/top_final_switch_0.VOUT[2] 5.92848
R12007 top_DAC_0/top_final_switch_0.VOUT[2].n5 top_DAC_0/top_final_switch_0.VOUT[2].n4 5.82758
R12008 top_DAC_0/top_final_switch_0.VOUT[2].n8 top_DAC_0/top_final_switch_0.VOUT[2].n7 5.29008
R12009 top_DAC_0/top_final_switch_0.VOUT[2].n9 top_DAC_0/top_final_switch_0.VOUT[2].n5 0.9505
R12010 top_DAC_0/top_final_switch_0.VOUT[2].n9 top_DAC_0/top_final_switch_0.VOUT[2].n8 0.767167
R12011 top_DAC_0/top_final_switch_0.VOUT[2].n10 top_DAC_0/top_final_switch_0.VOUT[2].n2 0.233364
R12012 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_final_switch_0.VOUT[2].n10 0.0275606
R12013 a_35132_8950.n0 a_35132_8950.t2 246.316
R12014 a_35132_8950.n0 a_35132_8950.t1 244.469
R12015 a_35132_8950.t0 a_35132_8950.n0 238.573
R12016 a_29434_6250.n2 a_29434_6250.t2 248.653
R12017 a_29434_6250.n0 a_29434_6250.t1 246.668
R12018 a_29434_6250.n1 a_29434_6250.t3 243.488
R12019 a_29434_6250.n0 a_29434_6250.t4 240
R12020 a_29434_6250.t0 a_29434_6250.n2 240
R12021 a_29434_6250.n2 a_29434_6250.n1 5.15258
R12022 a_29434_6250.n1 a_29434_6250.n0 1.86925
R12023 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t15 135.254
R12024 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t12 135.254
R12025 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n8 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t17 135.254
R12026 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t13 135.254
R12027 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t14 134.715
R12028 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t8 134.715
R12029 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t7 134.715
R12030 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t6 134.715
R12031 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n8 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t16 134.715
R12032 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n9 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t11 134.715
R12033 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t10 134.715
R12034 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t9 134.715
R12035 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n14 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t5 69.7645
R12036 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n11 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t1 60.7715
R12037 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n13 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t2 59.8932
R12038 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t4 59.8849
R12039 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n11 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t0 59.464
R12040 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t3 49.6789
R12041 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n0 15.0818
R12042 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n14 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n13 12.9172
R12043 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n12 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n11 9.36508
R12044 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n12 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n10 7.19425
R12045 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n14 3.55675
R12046 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n13 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n12 2.72758
R12047 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n10 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n5 1.9005
R12048 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n1 0.538
R12049 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n3 0.538
R12050 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n6 0.538
R12051 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n9 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n8 0.538
R12052 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n2 0.26925
R12053 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n4 0.26925
R12054 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n10 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n7 0.26925
R12055 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n10 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n9 0.26925
R12056 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 272.038
R12057 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t0 258.846
R12058 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t3 230.363
R12059 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n0 224.776
R12060 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t4 158.064
R12061 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n1 152.292
R12062 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t1 26.5955
R12063 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t2 26.5955
R12064 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 24.0946
R12065 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n2 20.0033
R12066 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 6.4005
R12067 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 3.76521
R12068 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n4 3.03935
R12069 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 2.30266
R12070 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n3 1.50638
R12071 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n5 0.921363
R12072 a_42982_22004.t0 a_42982_22004.t1 65.941
R12073 a_43240_22004.t0 a_43240_22004.t1 65.941
R12074 a_44255_3714.t0 a_44255_3714.t1 49.8467
R12075 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t0 272.038
R12076 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t0 258.846
R12077 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t3 241.536
R12078 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n0 224.776
R12079 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t4 169.237
R12080 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n1 152
R12081 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n2 31.596
R12082 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t1 26.5955
R12083 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t2 26.5955
R12084 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n3 22.9652
R12085 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 3.87418
R12086 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 3.76521
R12087 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n4 3.03935
R12088 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 2.63579
R12089 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n5 2.30266
R12090 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.921363
R12091 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t8 761.269
R12092 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t6 212.081
R12093 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t5 212.081
R12094 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 203.922
R12095 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 186.001
R12096 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t4 139.78
R12097 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t7 139.78
R12098 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 101.49
R12099 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 61.346
R12100 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t0 26.5955
R12101 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t1 26.5955
R12102 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t2 24.9236
R12103 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t3 24.9236
R12104 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y 13.5685
R12105 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y 10.7525
R12106 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 9.64425
R12107 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 9.30224
R12108 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y 6.6565
R12109 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 5.04292
R12110 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 3.8405
R12111 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.A 3.0725
R12112 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 2.5605
R12113 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y 1.93989
R12114 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t4 769.742
R12115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 203.923
R12116 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 101.49
R12117 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t3 26.5955
R12118 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t2 26.5955
R12119 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t0 24.9236
R12120 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t1 24.9236
R12121 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 13.0565
R12122 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 10.7525
R12123 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y 6.6565
R12124 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y 5.04292
R12125 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y 4.3525
R12126 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y 2.5605
R12127 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 1.93989
R12128 a_34856_8950.n0 a_34856_8950.t2 246.133
R12129 a_34856_8950.n0 a_34856_8950.t1 244.286
R12130 a_34856_8950.t0 a_34856_8950.n0 238.756
R12131 a_35453_10031.n0 a_35453_10031.t2 242.075
R12132 a_35453_10031.t0 a_35453_10031.n0 241.441
R12133 a_35453_10031.n0 a_35453_10031.t1 239.083
R12134 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.n0 680.072
R12135 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.t1 10.7276
R12136 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.t2 10.6922
R12137 a_15374_19866.n0 a_15374_19866.t1 671.848
R12138 a_15374_19866.n0 a_15374_19866.t2 666.814
R12139 a_15374_19866.t0 a_15374_19866.n0 665.327
R12140 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t1 334.788
R12141 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t8 213.218
R12142 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t22 213.218
R12143 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t19 213.218
R12144 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t6 212.887
R12145 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t13 212.554
R12146 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t12 212.554
R12147 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t9 212.554
R12148 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t7 212.554
R12149 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t4 212.554
R12150 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t23 212.554
R12151 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t5 212.554
R12152 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t2 212.554
R12153 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t24 212.554
R12154 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t21 212.554
R12155 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t20 212.554
R12156 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t14 208.054
R12157 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t11 208.054
R12158 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t10 208.054
R12159 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n21 152
R12160 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t3 126.27
R12161 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t15 125.558
R12162 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t18 121.127
R12163 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t16 114.031
R12164 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t0 87.8063
R12165 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t17 81.5883
R12166 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n4 39.4293
R12167 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n20 28.2979
R12168 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 15.1345
R12169 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 13.0029
R12170 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n22 11.4706
R12171 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n2 5.73592
R12172 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n3 5.388
R12173 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 4.83223
R12174 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n16 4.5005
R12175 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n18 4.5005
R12176 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 4.48881
R12177 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n17 2.59281
R12178 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n23 1.02758
R12179 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.7755
R12180 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n15 0.663962
R12181 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n14 0.663962
R12182 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n13 0.663962
R12183 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n12 0.663962
R12184 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n11 0.663962
R12185 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n5 0.663962
R12186 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n6 0.663962
R12187 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n7 0.663962
R12188 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n8 0.663962
R12189 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n9 0.663962
R12190 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n10 0.663962
R12191 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n0 0.322615
R12192 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n19 0.291365
R12193 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n1 0.177583
R12194 a_30608_7686.n2 a_30608_7686.t3 246.429
R12195 a_30608_7686.n0 a_30608_7686.t1 241.959
R12196 a_30608_7686.n0 a_30608_7686.t2 239.822
R12197 a_30608_7686.n1 a_30608_7686.t4 239.143
R12198 a_30608_7686.t0 a_30608_7686.n2 239.143
R12199 a_30608_7686.n2 a_30608_7686.n1 6.788
R12200 a_30608_7686.n1 a_30608_7686.n0 3.76508
R12201 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43.t2 248.95
R12202 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43.t1 10.575
R12203 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43.t0 10.5739
R12204 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43.n0 2.81389
R12205 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t2 676.833
R12206 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t1 10.7929
R12207 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.n0 10.5295
R12208 a_44062_18449.t0 a_44062_18449.t1 129.28
R12209 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 593.396
R12210 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 231.554
R12211 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 140.53
R12212 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 26.5955
R12213 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 26.5955
R12214 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 16.5652
R12215 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 9.03579
R12216 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 6.02403
R12217 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 1.72748
R12218 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 593.158
R12219 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 231.554
R12220 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 140.53
R12221 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 26.5955
R12222 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 26.5955
R12223 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 16.5652
R12224 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 9.03579
R12225 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 6.02403
R12226 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 1.72748
R12227 a_44062_18093.t0 a_44062_18093.t1 129.28
R12228 a_16596_18696.t0 a_16596_18696.n0 671.159
R12229 a_16596_18696.n0 a_16596_18696.t2 666.597
R12230 a_16596_18696.n0 a_16596_18696.t1 665.672
R12231 a_15066_18696.n0 a_15066_18696.t1 669.294
R12232 a_15066_18696.t0 a_15066_18696.n1 666.299
R12233 a_15066_18696.n1 a_15066_18696.t2 665.667
R12234 a_15066_18696.n0 a_15066_18696.t3 665.664
R12235 a_15066_18696.n1 a_15066_18696.n0 2.7505
R12236 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t5 230.155
R12237 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t2 229.369
R12238 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t1 221.538
R12239 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n0 157.927
R12240 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t3 157.856
R12241 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t4 157.07
R12242 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t0 152.889
R12243 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n1 152
R12244 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n3 24.6696
R12245 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n2 19.6746
R12246 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 17.3671
R12247 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n4 14.023
R12248 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 13.8127
R12249 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n5 2.22659
R12250 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 2.13383
R12251 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 1.55202
R12252 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.602583
R12253 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 593.165
R12254 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 268.077
R12255 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 258.846
R12256 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 237.577
R12257 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 26.5955
R12258 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 26.5955
R12259 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 16.5652
R12260 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 9.03579
R12261 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 8.8386
R12262 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 1.72748
R12263 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n1 863.124
R12264 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n0 585
R12265 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t0 495.469
R12266 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t2 220.327
R12267 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t8 217.555
R12268 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t13 217.555
R12269 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t17 216.893
R12270 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t14 216.893
R12271 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t4 216.893
R12272 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t7 216.893
R12273 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t11 216.893
R12274 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t3 216.893
R12275 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t6 213.218
R12276 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t18 212.77
R12277 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t15 212.554
R12278 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t19 212.554
R12279 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t16 212.554
R12280 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t5 212.554
R12281 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t9 212.554
R12282 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t20 212.393
R12283 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t10 212.393
R12284 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t12 208.054
R12285 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t1 141.189
R12286 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t0 140.738
R12287 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n15 39.9172
R12288 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n23 18.2588
R12289 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n14 14.6859
R12290 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 14.3755
R12291 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n22 14.1963
R12292 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n11 14.1776
R12293 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 11.6369
R12294 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 10.1408
R12295 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n24 8.53383
R12296 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n3 7.94225
R12297 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 7.20675
R12298 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 6.14988
R12299 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 5.81868
R12300 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n13 4.5005
R12301 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n10 4.5005
R12302 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n21 4.5005
R12303 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 2.16154
R12304 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n12 1.47133
R12305 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n2 0.665435
R12306 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n4 0.663962
R12307 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n5 0.663962
R12308 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n6 0.663962
R12309 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n7 0.663962
R12310 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n8 0.663962
R12311 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n9 0.663962
R12312 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n16 0.663962
R12313 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n17 0.663962
R12314 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n18 0.663962
R12315 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n19 0.663962
R12316 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n20 0.663962
R12317 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.447615
R12318 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.322615
R12319 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.226462
R12320 a_14615_14283.t0 a_14615_14283.n0 439.543
R12321 a_14615_14283.n0 a_14615_14283.t2 39.3576
R12322 a_14615_14283.n0 a_14615_14283.t1 39.3576
R12323 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t2 673.212
R12324 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t0 10.7613
R12325 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t1 10.7113
R12326 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.n0 2.72292
R12327 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t2 673.572
R12328 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t1 10.7178
R12329 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t0 10.6903
R12330 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.n0 3.41701
R12331 a_20823_20174.t0 a_20823_20174.n2 251.168
R12332 a_20823_20174.n0 a_20823_20174.t3 250.329
R12333 a_20823_20174.n2 a_20823_20174.t4 241.082
R12334 a_20823_20174.n1 a_20823_20174.t2 239.465
R12335 a_20823_20174.n0 a_20823_20174.t1 239.465
R12336 a_20823_20174.n1 a_20823_20174.n0 0.633833
R12337 a_20823_20174.n2 a_20823_20174.n1 0.20675
R12338 a_14055_6250.n2 a_14055_6250.t4 672.278
R12339 a_14055_6250.n0 a_14055_6250.t3 671.904
R12340 a_14055_6250.n1 a_14055_6250.t2 671.547
R12341 a_14055_6250.n0 a_14055_6250.t1 665.484
R12342 a_14055_6250.t0 a_14055_6250.n2 665.484
R12343 a_14055_6250.n2 a_14055_6250.n1 4.99842
R12344 a_14055_6250.n1 a_14055_6250.n0 1.563
R12345 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t2 663.232
R12346 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t1 10.6701
R12347 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.n0 10.5739
R12348 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1.t1 236.657
R12349 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1.n0 10.6906
R12350 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1.t2 10.5739
R12351 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2.t2 248.405
R12352 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2.t1 10.5394
R12353 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2.t0 10.5295
R12354 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2.n0 0.791214
R12355 a_42982_18130.t0 a_42982_18130.t1 65.941
R12356 a_43240_18130.t0 a_43240_18130.t1 65.941
R12357 a_42982_19896.t0 a_42982_19896.t1 65.941
R12358 a_43240_19896.t0 a_43240_19896.t1 65.941
R12359 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t1 134.734
R12360 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t2 134.734
R12361 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t0 134.734
R12362 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t3 134.734
R12363 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n1 79.7972
R12364 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n3 79.7972
R12365 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n2 79.7972
R12366 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n0 79.6389
R12367 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n5 11.8125
R12368 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t11 9.23217
R12369 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t6 9.23217
R12370 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t5 9.23217
R12371 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t8 9.23217
R12372 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t7 9.23217
R12373 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t10 9.23217
R12374 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t9 9.23217
R12375 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t4 9.23217
R12376 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n6 8.03342
R12377 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n7 5.19579
R12378 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n8 0.429667
R12379 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n4 0.429667
R12380 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n9 0.158833
R12381 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t1 672.309
R12382 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t0 10.8249
R12383 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t2 10.5739
R12384 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.n0 1.38332
R12385 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t1 673.491
R12386 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t2 10.7472
R12387 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t0 10.6536
R12388 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.n0 0.679794
R12389 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t2 227.827
R12390 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t1 227.827
R12391 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t5 227.827
R12392 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t4 227.827
R12393 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t6 226.506
R12394 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t3 226.506
R12395 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t7 226.506
R12396 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t0 226.506
R12397 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t14 221.911
R12398 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t8 221.911
R12399 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t12 221.911
R12400 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t13 221.911
R12401 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t11 221.911
R12402 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t15 221.911
R12403 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t9 221.911
R12404 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t10 221.911
R12405 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n10 8.30397
R12406 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n8 6.99147
R12407 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n7 6.73731
R12408 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n11 5.4248
R12409 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n2 4.30208
R12410 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n9 4.05141
R12411 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n12 3.4105
R12412 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n5 3.4105
R12413 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n0 3.12967
R12414 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n4 1.81717
R12415 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n3 1.563
R12416 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n6 0.655651
R12417 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n13 0.362258
R12418 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n1 0.2505
R12419 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t14 142.597
R12420 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t15 141.03
R12421 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t3 139.588
R12422 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t1 139.588
R12423 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t13 134.712
R12424 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n12 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t4 134.712
R12425 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t8 134.712
R12426 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n14 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t6 134.712
R12427 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t10 134.712
R12428 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n16 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t5 134.712
R12429 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t2 134.712
R12430 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t12 134.712
R12431 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t0 134.712
R12432 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t9 134.712
R12433 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t11 134.712
R12434 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n9 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t7 134.712
R12435 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n1 79.7972
R12436 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n3 79.7972
R12437 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n2 79.7972
R12438 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n0 79.6389
R12439 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t20 9.23217
R12440 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t17 9.23217
R12441 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t18 9.23217
R12442 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t23 9.23217
R12443 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t16 9.23217
R12444 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t21 9.23217
R12445 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t22 9.23217
R12446 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t19 9.23217
R12447 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n6 7.83383
R12448 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n15 7.83383
R12449 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n19 5.12671
R12450 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n12 4.61407
R12451 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n14 4.61407
R12452 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n17 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n16 4.61407
R12453 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n5 4.61407
R12454 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n8 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n7 4.61407
R12455 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n9 4.61407
R12456 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n11 3.97054
R12457 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n18 3.45425
R12458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n10 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n8 3.13383
R12459 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n15 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n13 3.13383
R12460 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n18 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n17 3.01092
R12461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n10 1.44425
R12462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n21 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n20 0.429667
R12463 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n20 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n4 0.429667
R12464 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n21 0.158833
R12465 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.n0 677.378
R12466 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.t2 10.7234
R12467 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.t1 10.6683
R12468 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.t1 249.345
R12469 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.t0 10.575
R12470 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.t2 10.5739
R12471 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.n0 4.20587
R12472 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58.t1 249.886
R12473 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58.t0 10.6257
R12474 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58.t2 10.5285
R12475 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58.n0 3.48476
R12476 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.n0 239.32
R12477 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.t1 10.716
R12478 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.t2 10.6698
R12479 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14.t1 238.232
R12480 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14.t2 10.5771
R12481 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14.n0 10.5739
R12482 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15.t1 237.542
R12483 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15.n0 10.5334
R12484 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15.t2 10.5312
R12485 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4.t1 677.225
R12486 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4.t2 10.7534
R12487 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4.n0 10.7113
R12488 a_14672_18696.n1 a_14672_18696.t2 671.525
R12489 a_14672_18696.n0 a_14672_18696.t1 668.735
R12490 a_14672_18696.t0 a_14672_18696.n1 666.038
R12491 a_14672_18696.n0 a_14672_18696.t3 665.865
R12492 a_14672_18696.n1 a_14672_18696.n0 0.365083
R12493 a_35757_10031.t0 a_35757_10031.n0 241.258
R12494 a_35757_10031.n0 a_35757_10031.t2 240.909
R12495 a_35757_10031.n0 a_35757_10031.t1 238.899
R12496 a_43724_12342.t0 a_43724_12342.t1 55.3905
R12497 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 272.038
R12498 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t1 258.846
R12499 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t3 230.363
R12500 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n5 224.775
R12501 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t4 158.064
R12502 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n0 153.28
R12503 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t2 26.5955
R12504 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t0 26.5955
R12505 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n1 19.4367
R12506 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 5.1205
R12507 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n4 3.76521
R12508 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n3 3.03935
R12509 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n2 1.56597
R12510 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.921363
R12511 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n2 0.737191
R12512 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t4 151.438
R12513 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t5 149.923
R12514 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n6 79.7972
R12515 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n2 79.7972
R12516 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n1 79.7972
R12517 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n0 79.6389
R12518 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t6 9.23217
R12519 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t2 9.23217
R12520 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t0 9.23217
R12521 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t8 9.23217
R12522 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t9 9.23217
R12523 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t1 9.23217
R12524 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t3 9.23217
R12525 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t7 9.23217
R12526 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n4 4.75071
R12527 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n7 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n5 0.429667
R12528 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n5 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n3 0.429667
R12529 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n7 0.158833
R12530 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t4 748.038
R12531 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 237.577
R12532 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t3 230.576
R12533 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t5 158.275
R12534 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 152.8
R12535 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t1 139.514
R12536 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t2 26.5955
R12537 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t0 26.5955
R12538 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y 16.1887
R12539 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 10.0771
R12540 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 9.63258
R12541 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 9.41227
R12542 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y 6.98232
R12543 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_0.A 5.86717
R12544 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[3] 5.74157
R12545 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y 2.23542
R12546 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[3] 0.830857
R12547 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 0.508436
R12548 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 0.291409
R12549 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7.t2 248.075
R12550 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7.t1 10.5773
R12551 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7.t0 10.5739
R12552 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7.n0 4.31612
R12553 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.t1 249.738
R12554 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.t2 13.5844
R12555 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.t0 10.8964
R12556 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.n0 4.7255
R12557 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t0 227.856
R12558 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n2 152.333
R12559 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t3 140.382
R12560 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t4 114.031
R12561 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t1 83.3993
R12562 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t2 81.5883
R12563 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n3 14.4422
R12564 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n1 7.56882
R12565 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n0 5.08175
R12566 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R12567 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t0 673.212
R12568 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t2 10.7577
R12569 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t1 10.7161
R12570 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.n0 2.72817
R12571 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49.n0 236.649
R12572 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49.t2 10.6713
R12573 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49.t1 10.5739
R12574 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50.t0 246.716
R12575 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50.t2 10.5296
R12576 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50.t1 10.5285
R12577 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50.n0 0.886534
R12578 a_43240_18814.t0 a_43240_18814.t1 65.941
R12579 a_21651_20174.n0 a_21651_20174.t2 251.719
R12580 a_21651_20174.t0 a_21651_20174.n1 248.475
R12581 a_21651_20174.n0 a_21651_20174.t3 241.631
R12582 a_21651_20174.n1 a_21651_20174.t1 238.916
R12583 a_21651_20174.n1 a_21651_20174.n0 3.24425
R12584 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t4 743.342
R12585 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n7 586.745
R12586 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n6 289.24
R12587 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t5 230.576
R12588 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t3 158.275
R12589 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n2 152
R12590 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n0 94.1864
R12591 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n5 82.6525
R12592 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t1 26.5955
R12593 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t2 24.9236
R12594 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t0 24.9236
R12595 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n4 21.3341
R12596 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n6 17.9639
R12597 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n3 9.3005
R12598 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_1.A 6.66717
R12599 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[1] 3.48572
R12600 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[1] 0.790679
R12601 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[1] 0.063
R12602 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n1 0.063
R12603 a_42847_4906.t0 a_42847_4906.t1 41.3705
R12604 a_30332_7686.n2 a_30332_7686.t2 246.244
R12605 a_30332_7686.n0 a_30332_7686.t1 241.385
R12606 a_30332_7686.n0 a_30332_7686.t3 240.358
R12607 a_30332_7686.n1 a_30332_7686.t4 238.959
R12608 a_30332_7686.t0 a_30332_7686.n2 238.959
R12609 a_30332_7686.n2 a_30332_7686.n1 6.788
R12610 a_30332_7686.n1 a_30332_7686.n0 4.15675
R12611 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.t2 250.332
R12612 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.t0 10.5317
R12613 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.t1 10.5285
R12614 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.n0 3.51046
R12615 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t4 739.633
R12616 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t9 229.369
R12617 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t12 229.369
R12618 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t7 212.081
R12619 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t6 212.081
R12620 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 203.922
R12621 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 186.001
R12622 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t5 157.07
R12623 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t8 157.07
R12624 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 152.712
R12625 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 152.475
R12626 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t11 139.78
R12627 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t10 139.78
R12628 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 101.49
R12629 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 61.346
R12630 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t0 26.5955
R12631 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t1 26.5955
R12632 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t2 24.9236
R12633 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t3 24.9236
R12634 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 15.8609
R12635 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[0] 13.7651
R12636 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y 13.5685
R12637 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y 10.7525
R12638 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 10.2234
R12639 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 9.77342
R12640 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 9.64425
R12641 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 9.30224
R12642 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y 6.6565
R12643 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.B 5.45235
R12644 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.B 5.21532
R12645 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 5.04292
R12646 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 4.91925
R12647 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 3.8405
R12648 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.A 3.0725
R12649 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 2.5605
R12650 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y 1.93989
R12651 a_44234_14916.t0 a_44234_14916.t1 114.052
R12652 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t2 274.793
R12653 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t4 232.214
R12654 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n0 205.28
R12655 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t1 169.452
R12656 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t5 159.915
R12657 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n2 152.207
R12658 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n1 54.4975
R12659 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t3 26.5955
R12660 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t0 26.5955
R12661 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n3 20.6093
R12662 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n4 12.9887
R12663 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 4.54244
R12664 a_44234_15906.t0 a_44234_15906.t1 114.052
R12665 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n1 863.124
R12666 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n0 585
R12667 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t0 495.469
R12668 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t5 217.555
R12669 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t4 217.555
R12670 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t3 217.555
R12671 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t17 216.893
R12672 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t15 216.893
R12673 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t7 216.893
R12674 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t10 216.893
R12675 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t9 216.893
R12676 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t11 216.893
R12677 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t16 216.893
R12678 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t14 216.893
R12679 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t6 216.893
R12680 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t2 216.893
R12681 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t12 216.893
R12682 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t13 212.393
R12683 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t8 212.393
R12684 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t1 141.189
R12685 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t0 140.738
R12686 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n18 109.279
R12687 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n19 13.9817
R12688 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 11.6369
R12689 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 10.1408
R12690 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n3 7.94225
R12691 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n20 7.56414
R12692 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 6.78838
R12693 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 6.14988
R12694 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n15 4.5005
R12695 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n17 4.5005
R12696 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 2.16154
R12697 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n16 1.88512
R12698 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.7755
R12699 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.6755
R12700 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n2 0.665435
R12701 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n14 0.663962
R12702 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n13 0.663962
R12703 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n12 0.663962
R12704 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n11 0.663962
R12705 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n10 0.663962
R12706 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n4 0.663962
R12707 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n5 0.663962
R12708 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n6 0.663962
R12709 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n7 0.663962
R12710 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n8 0.663962
R12711 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n9 0.663962
R12712 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53.t0 246.63
R12713 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53.t1 10.6701
R12714 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53.t2 10.5739
R12715 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53.n0 2.77493
R12716 a_28882_6250.n2 a_28882_6250.t2 248.286
R12717 a_28882_6250.n0 a_28882_6250.t1 246.303
R12718 a_28882_6250.n1 a_28882_6250.t3 244.629
R12719 a_28882_6250.n0 a_28882_6250.t4 239.633
R12720 a_28882_6250.t0 a_28882_6250.n2 239.633
R12721 a_28882_6250.n2 a_28882_6250.n1 5.93592
R12722 a_28882_6250.n1 a_28882_6250.n0 1.08592
R12723 a_44062_21653.t0 a_44062_21653.t1 129.28
R12724 a_39936_22083.t0 a_39936_22083.n0 356.854
R12725 a_39936_22083.n0 a_39936_22083.t2 15.3866
R12726 a_39936_22083.n0 a_39936_22083.t1 15.3866
R12727 a_8051_10107.n9 a_8051_10107.t9 221.913
R12728 a_8051_10107.n8 a_8051_10107.t8 221.913
R12729 a_8051_10107.n3 a_8051_10107.t6 221.913
R12730 a_8051_10107.n9 a_8051_10107.t7 221.911
R12731 a_8051_10107.n8 a_8051_10107.t11 221.911
R12732 a_8051_10107.n3 a_8051_10107.t10 221.911
R12733 a_8051_10107.n5 a_8051_10107.t4 221.851
R12734 a_8051_10107.n6 a_8051_10107.t5 221.851
R12735 a_8051_10107.n14 a_8051_10107.n13 71.3963
R12736 a_8051_10107.n2 a_8051_10107.n1 71.3963
R12737 a_8051_10107.n2 a_8051_10107.n0 71.3963
R12738 a_8051_10107.n15 a_8051_10107.n14 71.3963
R12739 a_8051_10107.n13 a_8051_10107.t14 16.5305
R12740 a_8051_10107.n13 a_8051_10107.t1 16.5305
R12741 a_8051_10107.n1 a_8051_10107.t2 16.5305
R12742 a_8051_10107.n1 a_8051_10107.t13 16.5305
R12743 a_8051_10107.n0 a_8051_10107.t15 16.5305
R12744 a_8051_10107.n0 a_8051_10107.t0 16.5305
R12745 a_8051_10107.t3 a_8051_10107.n15 16.5305
R12746 a_8051_10107.n15 a_8051_10107.t12 16.5305
R12747 a_8051_10107.n4 a_8051_10107.n3 6.97216
R12748 a_8051_10107.n10 a_8051_10107.n9 5.78883
R12749 a_8051_10107.n7 a_8051_10107.n6 4.97106
R12750 a_8051_10107.n5 a_8051_10107.n4 4.97106
R12751 a_8051_10107.n11 a_8051_10107.n7 4.69233
R12752 a_8051_10107.n12 a_8051_10107.n11 4.3975
R12753 a_8051_10107.n10 a_8051_10107.n8 3.69924
R12754 a_8051_10107.n11 a_8051_10107.n10 3.4105
R12755 a_8051_10107.n14 a_8051_10107.n12 0.3505
R12756 a_8051_10107.n12 a_8051_10107.n2 0.3505
R12757 a_8051_10107.n7 a_8051_10107.n4 0.246333
R12758 a_8051_10107.n6 a_8051_10107.n5 0.123417
R12759 a_44234_14282.t0 a_44234_14282.t1 114.052
R12760 a_43698_13726.t0 a_43698_13726.n0 228.04
R12761 a_43698_13726.n0 a_43698_13726.t2 145.648
R12762 a_43698_13726.n0 a_43698_13726.t1 83.2159
R12763 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55.t0 248.075
R12764 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55.t2 10.6701
R12765 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55.t1 10.5739
R12766 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55.n0 4.16691
R12767 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45.t1 249.321
R12768 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45.t2 10.6671
R12769 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45.t0 10.5769
R12770 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45.n0 1.55078
R12771 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44.t1 249.209
R12772 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44.t2 10.5296
R12773 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44.t0 10.5295
R12774 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44.n0 2.13671
R12775 top_DAC_0/top_rseg_n_dcell_0.VS4.n5 top_DAC_0/top_rseg_n_dcell_0.VS4.t0 665.933
R12776 top_DAC_0/top_rseg_n_dcell_0.VS4.n0 top_DAC_0/top_rseg_n_dcell_0.VS4.t6 660.876
R12777 top_DAC_0/top_rseg_n_dcell_0.VS4.n4 top_DAC_0/top_rseg_n_dcell_0.VS4.t1 660.799
R12778 top_DAC_0/top_rseg_n_dcell_0.VS4.n3 top_DAC_0/top_rseg_n_dcell_0.VS4.t3 660.24
R12779 top_DAC_0/top_rseg_n_dcell_0.VS4.n2 top_DAC_0/top_rseg_n_dcell_0.VS4.t5 660.24
R12780 top_DAC_0/top_rseg_n_dcell_0.VS4.n1 top_DAC_0/top_rseg_n_dcell_0.VS4.t2 660.24
R12781 top_DAC_0/top_rseg_n_dcell_0.VS4.n0 top_DAC_0/top_rseg_n_dcell_0.VS4.t4 660.24
R12782 top_DAC_0/top_rseg_n_dcell_0.VS4.n4 top_DAC_0/top_rseg_n_dcell_0.VS4 20.2526
R12783 top_DAC_0/top_rseg_n_dcell_0.VS4.n5 top_DAC_0/top_rseg_n_dcell_0.VS4.n4 4.5005
R12784 top_DAC_0/top_rseg_n_dcell_0.VS4.n1 top_DAC_0/top_rseg_n_dcell_0.VS4.n0 0.63637
R12785 top_DAC_0/top_rseg_n_dcell_0.VS4.n2 top_DAC_0/top_rseg_n_dcell_0.VS4.n1 0.63637
R12786 top_DAC_0/top_rseg_n_dcell_0.VS4.n3 top_DAC_0/top_rseg_n_dcell_0.VS4.n2 0.63637
R12787 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.VS4.n3 0.465083
R12788 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.VS4.n5 0.063
R12789 a_19468_10031.n0 a_19468_10031.t2 666.692
R12790 a_19468_10031.t0 a_19468_10031.n0 666.317
R12791 a_19468_10031.n0 a_19468_10031.t1 665.484
R12792 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.VH3.t3 666.581
R12793 top_DAC_0/top_rseg_n_dcell_0.VH3.n1 top_DAC_0/top_rseg_n_dcell_0.VH3.t4 660.933
R12794 top_DAC_0/top_rseg_n_dcell_0.VH3.n2 top_DAC_0/top_rseg_n_dcell_0.VH3.t1 660.876
R12795 top_DAC_0/top_rseg_n_dcell_0.VH3.n2 top_DAC_0/top_rseg_n_dcell_0.VH3.t2 660.24
R12796 top_DAC_0/top_rseg_n_dcell_0.VH3.n3 top_DAC_0/top_rseg_n_dcell_0.VH3.t0 660.24
R12797 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.VH3.n1 26.7547
R12798 top_DAC_0/top_rseg_n_dcell_0.VH3.n1 top_DAC_0/top_rseg_n_dcell_0.VH3.n0 4.5005
R12799 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.VH3.n3 1.5255
R12800 top_DAC_0/top_rseg_n_dcell_0.VH3.n3 top_DAC_0/top_rseg_n_dcell_0.VH3.n2 0.63637
R12801 top_DAC_0/top_rseg_n_dcell_0.VH3.n0 top_DAC_0/top_rseg_n_dcell_0.VH3 0.063
R12802 top_DAC_0/top_rseg_n_dcell_0.VH3.n0 top_DAC_0/top_rseg_n_dcell_0.VH3 0.0588333
R12803 a_15863_13287.t0 a_15863_13287.n0 1266.9
R12804 a_15863_13287.n0 a_15863_13287.t1 65.941
R12805 a_15863_13287.n0 a_15863_13287.t2 65.941
R12806 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t10 142.488
R12807 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t12 142.488
R12808 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t6 142.488
R12809 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t11 141.704
R12810 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t7 141.704
R12811 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t8 141.704
R12812 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t13 141.704
R12813 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t9 141.704
R12814 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t2 139.454
R12815 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t0 139.454
R12816 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t5 135.329
R12817 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t1 135.231
R12818 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t3 135.231
R12819 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t4 134.444
R12820 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n0 6.41092
R12821 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n11 4.563
R12822 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n8 2.2505
R12823 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n4 2.2505
R12824 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n5 0.829667
R12825 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n9 0.829667
R12826 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n6 0.783833
R12827 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n7 0.783833
R12828 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n1 0.783833
R12829 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n2 0.783833
R12830 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n3 0.783833
R12831 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n10 0.224458
R12832 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t0 158.145
R12833 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t2 142.477
R12834 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t3 140.496
R12835 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t1 140.082
R12836 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n0 7.35744
R12837 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n1 0.0463333
R12838 top_DAC_0/top_rseg_n_dcell_0.SH[4].n2 top_DAC_0/top_rseg_n_dcell_0.SH[4].n1 863.124
R12839 top_DAC_0/top_rseg_n_dcell_0.SH[4].n1 top_DAC_0/top_rseg_n_dcell_0.SH[4].n0 585
R12840 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.SH[4].t0 495.469
R12841 top_DAC_0/top_rseg_n_dcell_0.SH[4].n4 top_DAC_0/top_rseg_n_dcell_0.SH[4].t5 213.375
R12842 top_DAC_0/top_rseg_n_dcell_0.SH[4].n7 top_DAC_0/top_rseg_n_dcell_0.SH[4].t2 212.393
R12843 top_DAC_0/top_rseg_n_dcell_0.SH[4].n6 top_DAC_0/top_rseg_n_dcell_0.SH[4].t4 212.393
R12844 top_DAC_0/top_rseg_n_dcell_0.SH[4].n5 top_DAC_0/top_rseg_n_dcell_0.SH[4].t6 212.393
R12845 top_DAC_0/top_rseg_n_dcell_0.SH[4].n4 top_DAC_0/top_rseg_n_dcell_0.SH[4].t3 212.393
R12846 top_DAC_0/top_rseg_n_dcell_0.SH[4].n3 top_DAC_0/top_rseg_n_dcell_0.SH[4].t1 141.189
R12847 top_DAC_0/top_rseg_n_dcell_0.SH[4].n1 top_DAC_0/top_rseg_n_dcell_0.SH[4].t0 140.738
R12848 top_DAC_0/top_rseg_n_dcell_0.SH[4].n8 top_DAC_0/top_rseg_n_dcell_0.SH[4] 14.5776
R12849 top_DAC_0/top_rseg_n_dcell_0.SH[4].n2 top_DAC_0/top_rseg_n_dcell_0.SH[4] 11.6369
R12850 top_DAC_0/top_rseg_n_dcell_0.SH[4].n0 top_DAC_0/top_rseg_n_dcell_0.SH[4] 10.1408
R12851 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.SH[4].n8 8.14595
R12852 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.SH[4].n3 7.94225
R12853 top_DAC_0/top_rseg_n_dcell_0.SH[4].n8 top_DAC_0/top_rseg_n_dcell_0.SH[4] 6.20656
R12854 top_DAC_0/top_rseg_n_dcell_0.SH[4].n3 top_DAC_0/top_rseg_n_dcell_0.SH[4] 6.14988
R12855 top_DAC_0/top_rseg_n_dcell_0.SH[4].n0 top_DAC_0/top_rseg_n_dcell_0.SH[4] 2.16154
R12856 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.SH[4].n7 1.39101
R12857 top_DAC_0/top_rseg_n_dcell_0.SH[4].n5 top_DAC_0/top_rseg_n_dcell_0.SH[4].n4 0.982408
R12858 top_DAC_0/top_rseg_n_dcell_0.SH[4].n6 top_DAC_0/top_rseg_n_dcell_0.SH[4].n5 0.982408
R12859 top_DAC_0/top_rseg_n_dcell_0.SH[4].n7 top_DAC_0/top_rseg_n_dcell_0.SH[4].n6 0.982408
R12860 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.SH[4].n2 0.665435
R12861 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1.t1 663.775
R12862 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1.n0 10.6257
R12863 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1.t2 10.5285
R12864 a_16872_18696.n0 a_16872_18696.t1 670.976
R12865 a_16872_18696.n0 a_16872_18696.t2 666.78
R12866 a_16872_18696.t0 a_16872_18696.n0 665.487
R12867 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n1 863.124
R12868 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n0 585
R12869 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t0 495.469
R12870 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t10 217.555
R12871 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t2 216.893
R12872 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t7 216.893
R12873 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t4 216.893
R12874 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t6 216.893
R12875 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t9 216.893
R12876 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t5 216.893
R12877 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t8 216.893
R12878 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t3 216.893
R12879 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t1 141.189
R12880 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t0 140.738
R12881 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n12 79.1581
R12882 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 14.3755
R12883 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 11.6369
R12884 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 10.1408
R12885 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n13 8.53383
R12886 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n3 7.94225
R12887 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 6.14988
R12888 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 5.81868
R12889 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 2.16154
R12890 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n2 0.665435
R12891 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n10 0.663962
R12892 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n9 0.663962
R12893 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n8 0.663962
R12894 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n7 0.663962
R12895 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n6 0.663962
R12896 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n5 0.663962
R12897 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n4 0.663962
R12898 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n11 0.284841
R12899 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 0.0250536
R12900 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.t1 249.345
R12901 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.t2 10.6701
R12902 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.t0 10.5739
R12903 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.n0 4.15498
R12904 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26.t1 250.066
R12905 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26.t2 10.5296
R12906 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26.t0 10.5295
R12907 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26.n0 3.52631
R12908 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37.t2 246.63
R12909 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37.t1 10.575
R12910 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37.t0 10.5739
R12911 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37.n0 2.81913
R12912 DIN9.n1 DIN9.t2 212.081
R12913 DIN9.n0 DIN9.t0 212.081
R12914 DIN9.n2 DIN9.n1 183.185
R12915 DIN9.n1 DIN9.t1 139.78
R12916 DIN9.n0 DIN9.t3 139.78
R12917 DIN9.n1 DIN9.n0 61.346
R12918 DIN9 DIN9.n2 14.2776
R12919 DIN9.n2 DIN9 5.8885
R12920 top_DAC_0/top_rseg_n_dcell_0.SH[1].n2 top_DAC_0/top_rseg_n_dcell_0.SH[1].n1 863.124
R12921 top_DAC_0/top_rseg_n_dcell_0.SH[1].n1 top_DAC_0/top_rseg_n_dcell_0.SH[1].n0 585
R12922 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.SH[1].t0 495.469
R12923 top_DAC_0/top_rseg_n_dcell_0.SH[1].n4 top_DAC_0/top_rseg_n_dcell_0.SH[1].t2 209.036
R12924 top_DAC_0/top_rseg_n_dcell_0.SH[1].n7 top_DAC_0/top_rseg_n_dcell_0.SH[1].t4 208.054
R12925 top_DAC_0/top_rseg_n_dcell_0.SH[1].n6 top_DAC_0/top_rseg_n_dcell_0.SH[1].t6 208.054
R12926 top_DAC_0/top_rseg_n_dcell_0.SH[1].n5 top_DAC_0/top_rseg_n_dcell_0.SH[1].t3 208.054
R12927 top_DAC_0/top_rseg_n_dcell_0.SH[1].n4 top_DAC_0/top_rseg_n_dcell_0.SH[1].t5 208.054
R12928 top_DAC_0/top_rseg_n_dcell_0.SH[1].n3 top_DAC_0/top_rseg_n_dcell_0.SH[1].t1 141.189
R12929 top_DAC_0/top_rseg_n_dcell_0.SH[1].n1 top_DAC_0/top_rseg_n_dcell_0.SH[1].t0 140.738
R12930 top_DAC_0/top_rseg_n_dcell_0.SH[1].n8 top_DAC_0/top_rseg_n_dcell_0.SH[1] 14.5776
R12931 top_DAC_0/top_rseg_n_dcell_0.SH[1].n2 top_DAC_0/top_rseg_n_dcell_0.SH[1] 11.6369
R12932 top_DAC_0/top_rseg_n_dcell_0.SH[1].n0 top_DAC_0/top_rseg_n_dcell_0.SH[1] 10.1408
R12933 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.SH[1].n8 8.14595
R12934 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.SH[1].n3 7.94225
R12935 top_DAC_0/top_rseg_n_dcell_0.SH[1].n8 top_DAC_0/top_rseg_n_dcell_0.SH[1] 6.20656
R12936 top_DAC_0/top_rseg_n_dcell_0.SH[1].n3 top_DAC_0/top_rseg_n_dcell_0.SH[1] 6.14988
R12937 top_DAC_0/top_rseg_n_dcell_0.SH[1].n0 top_DAC_0/top_rseg_n_dcell_0.SH[1] 2.16154
R12938 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.SH[1].n7 1.30619
R12939 top_DAC_0/top_rseg_n_dcell_0.SH[1].n5 top_DAC_0/top_rseg_n_dcell_0.SH[1].n4 0.982408
R12940 top_DAC_0/top_rseg_n_dcell_0.SH[1].n6 top_DAC_0/top_rseg_n_dcell_0.SH[1].n5 0.982408
R12941 top_DAC_0/top_rseg_n_dcell_0.SH[1].n7 top_DAC_0/top_rseg_n_dcell_0.SH[1].n6 0.982408
R12942 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.SH[1].n2 0.665435
R12943 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.VS1.t1 239.155
R12944 top_DAC_0/top_rseg_n_dcell_0.VS1.n0 top_DAC_0/top_rseg_n_dcell_0.VS1.t6 234.293
R12945 top_DAC_0/top_rseg_n_dcell_0.VS1.n4 top_DAC_0/top_rseg_n_dcell_0.VS1.t0 234.216
R12946 top_DAC_0/top_rseg_n_dcell_0.VS1.n3 top_DAC_0/top_rseg_n_dcell_0.VS1.t4 233.657
R12947 top_DAC_0/top_rseg_n_dcell_0.VS1.n2 top_DAC_0/top_rseg_n_dcell_0.VS1.t3 233.657
R12948 top_DAC_0/top_rseg_n_dcell_0.VS1.n1 top_DAC_0/top_rseg_n_dcell_0.VS1.t5 233.657
R12949 top_DAC_0/top_rseg_n_dcell_0.VS1.n0 top_DAC_0/top_rseg_n_dcell_0.VS1.t2 233.657
R12950 top_DAC_0/top_rseg_n_dcell_0.VS1.n4 top_DAC_0/top_rseg_n_dcell_0.VS1 56.6505
R12951 top_DAC_0/top_rseg_n_dcell_0.VS1.n5 top_DAC_0/top_rseg_n_dcell_0.VS1.n4 4.5005
R12952 top_DAC_0/top_rseg_n_dcell_0.VS1.n1 top_DAC_0/top_rseg_n_dcell_0.VS1.n0 0.63637
R12953 top_DAC_0/top_rseg_n_dcell_0.VS1.n2 top_DAC_0/top_rseg_n_dcell_0.VS1.n1 0.63637
R12954 top_DAC_0/top_rseg_n_dcell_0.VS1.n3 top_DAC_0/top_rseg_n_dcell_0.VS1.n2 0.63637
R12955 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.VS1.n3 0.44425
R12956 top_DAC_0/top_rseg_n_dcell_0.VS1.n5 top_DAC_0/top_rseg_n_dcell_0.VS1 0.196333
R12957 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.VS1.n5 0.063
R12958 a_39306_20477.t0 a_39306_20477.n0 239.25
R12959 a_39306_20477.n0 a_39306_20477.t2 222.119
R12960 a_39306_20477.n0 a_39306_20477.t1 222.119
R12961 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n1 863.124
R12962 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n0 585
R12963 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t0 495.469
R12964 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t2 217.555
R12965 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t3 216.893
R12966 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t4 212.393
R12967 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t1 141.189
R12968 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t0 140.738
R12969 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n6 77.7359
R12970 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 14.3755
R12971 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 11.6369
R12972 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 10.1408
R12973 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n7 8.53383
R12974 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n3 7.94225
R12975 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 6.14988
R12976 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 5.81868
R12977 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n5 4.5005
R12978 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 2.16154
R12979 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n2 0.665435
R12980 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n4 0.663962
R12981 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.317808
R12982 a_16891_7686.n0 a_16891_7686.t1 672.581
R12983 a_16891_7686.n2 a_16891_7686.t3 670.423
R12984 a_16891_7686.t0 a_16891_7686.n2 666.391
R12985 a_16891_7686.n0 a_16891_7686.t4 666.092
R12986 a_16891_7686.n1 a_16891_7686.t2 666.092
R12987 a_16891_7686.n1 a_16891_7686.n0 6.63383
R12988 a_16891_7686.n2 a_16891_7686.n1 2.62342
R12989 a_43698_12736.t0 a_43698_12736.n0 228.04
R12990 a_43698_12736.n0 a_43698_12736.t2 145.648
R12991 a_43698_12736.n0 a_43698_12736.t1 83.2159
R12992 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t1 227.856
R12993 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n2 152.333
R12994 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t4 140.382
R12995 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t2 114.031
R12996 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t0 83.3993
R12997 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t3 81.5883
R12998 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n3 14.4422
R12999 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n1 7.56882
R13000 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n0 5.08175
R13001 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R13002 a_43724_12896.t0 a_43724_12896.t1 55.3905
R13003 a_17732_18696.n0 a_17732_18696.t2 667.216
R13004 a_17732_18696.n0 a_17732_18696.t1 666.692
R13005 a_17732_18696.t0 a_17732_18696.n0 665.433
R13006 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.t1 668.619
R13007 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.t0 238.077
R13008 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.t2 12.4069
R13009 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.t3 10.6569
R13010 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V48 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.n0 1.29821
R13011 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V48 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0.n1 0.397447
R13012 a_15353_7686.n1 a_15353_7686.t2 671.663
R13013 a_15353_7686.n0 a_15353_7686.t1 668.203
R13014 a_15353_7686.n0 a_15353_7686.t3 667.22
R13015 a_15353_7686.n1 a_15353_7686.t4 665.176
R13016 a_15353_7686.t0 a_15353_7686.n2 665.176
R13017 a_15353_7686.n2 a_15353_7686.n1 6.63383
R13018 a_15353_7686.n2 a_15353_7686.n0 4.91092
R13019 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t2 676.321
R13020 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t1 13.5968
R13021 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t0 10.7638
R13022 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.n0 4.72836
R13023 a_22203_20174.n0 a_22203_20174.t2 250.986
R13024 a_22203_20174.t0 a_22203_20174.n1 249.524
R13025 a_22203_20174.n0 a_22203_20174.t3 240.898
R13026 a_22203_20174.n1 a_22203_20174.t1 239.649
R13027 a_22203_20174.n1 a_22203_20174.n0 1.46092
R13028 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.t2 239.248
R13029 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.n0 10.7191
R13030 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.t1 10.6712
R13031 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2.t1 675.611
R13032 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2.t2 10.8307
R13033 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2.n0 10.5739
R13034 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3.t1 674.707
R13035 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3.n0 10.7559
R13036 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3.t2 10.6512
R13037 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n2 270.841
R13038 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t0 258.846
R13039 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t4 241.536
R13040 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n3 224.776
R13041 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t3 169.237
R13042 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n0 152
R13043 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n1 31.0273
R13044 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t1 26.5955
R13045 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t2 26.5955
R13046 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 3.92583
R13047 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 3.76521
R13048 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n4 3.03935
R13049 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n5 2.30266
R13050 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n2 1.19762
R13051 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.921363
R13052 a_27344_6250.n2 a_27344_6250.t2 247.369
R13053 a_27344_6250.n0 a_27344_6250.t1 245.386
R13054 a_27344_6250.n1 a_27344_6250.t3 244.766
R13055 a_27344_6250.n0 a_27344_6250.t4 238.716
R13056 a_27344_6250.t0 a_27344_6250.n2 238.716
R13057 a_27344_6250.n1 a_27344_6250.n0 5.07133
R13058 a_27344_6250.n2 a_27344_6250.n1 1.9505
R13059 a_33358_8950.n0 a_33358_8950.t2 244.542
R13060 a_33358_8950.n0 a_33358_8950.t1 242.81
R13061 a_33358_8950.t0 a_33358_8950.n0 239.857
R13062 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 593.154
R13063 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 268.077
R13064 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 258.846
R13065 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 231.554
R13066 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 26.5955
R13067 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 26.5955
R13068 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 16.5652
R13069 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 9.03579
R13070 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 8.8386
R13071 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 6.02403
R13072 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 1.72748
R13073 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.t2 238.876
R13074 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.t1 10.7601
R13075 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.n0 10.719
R13076 ROUT1.n1 ROUT1.t1 160.756
R13077 ROUT1.n1 ROUT1.t3 134.811
R13078 ROUT1.n3 ROUT1.t0 16.8154
R13079 ROUT1.n0 ROUT1.t4 16.8154
R13080 ROUT1.n2 ROUT1.n0 12.0038
R13081 ROUT1.n4 ROUT1.n3 6.5267
R13082 ROUT1.n3 ROUT1.t5 5.78822
R13083 ROUT1.n0 ROUT1.t2 5.78822
R13084 ROUT1.n4 ROUT1.n2 5.72758
R13085 ROUT1 ROUT1.n4 3.44682
R13086 ROUT1 ROUT1.n1 0.902583
R13087 ROUT1.n2 ROUT1 0.063
R13088 a_8473_23194.n1 a_8473_23194.n0 243.671
R13089 a_8473_23194.n0 a_8473_23194.t1 15.3866
R13090 a_8473_23194.n0 a_8473_23194.t3 15.3866
R13091 a_8473_23194.t0 a_8473_23194.n1 15.3866
R13092 a_8473_23194.n1 a_8473_23194.t2 15.3866
R13093 a_19552_8950.n0 a_19552_8950.t1 670.775
R13094 a_19552_8950.n0 a_19552_8950.t2 670.366
R13095 a_19552_8950.t0 a_19552_8950.n0 665.89
R13096 a_20076_10031.n0 a_20076_10031.t2 670.216
R13097 a_20076_10031.n0 a_20076_10031.t1 668.208
R13098 a_20076_10031.t0 a_20076_10031.n0 665.85
R13099 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t9 142.488
R13100 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t12 142.488
R13101 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t13 142.488
R13102 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t7 142.488
R13103 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t11 141.704
R13104 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t8 141.704
R13105 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t6 141.704
R13106 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t10 141.704
R13107 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t2 139.454
R13108 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t4 139.454
R13109 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t1 135.305
R13110 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t3 135.246
R13111 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t5 135.246
R13112 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t0 135.244
R13113 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n12 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n11 12.38
R13114 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n0 5.038
R13115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n10 4.5005
R13116 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n7 2.2505
R13117 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n3 2.2505
R13118 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n4 0.842167
R13119 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n8 0.842167
R13120 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n5 0.783833
R13121 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n6 0.783833
R13122 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n1 0.783833
R13123 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n2 0.783833
R13124 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n0 0.26925
R13125 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n9 0.26925
R13126 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n12 0.063
R13127 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t1 158.273
R13128 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t2 141.358
R13129 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t0 140.304
R13130 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t3 139.566
R13131 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n0 8.02027
R13132 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n1 0.063
R13133 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t8 217.037
R13134 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t9 217.037
R13135 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t6 211.755
R13136 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t7 211.755
R13137 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t0 60.8179
R13138 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t2 60.0612
R13139 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t5 59.4176
R13140 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t1 50.7632
R13141 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t4 50.7591
R13142 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t3 49.6518
R13143 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n2 13.3067
R13144 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n4 5.57275
R13145 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n0 5.26748
R13146 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n5 5.03383
R13147 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n7 4.92133
R13148 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n6 3.04842
R13149 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n1 0.565401
R13150 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n3 0.189786
R13151 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t1 227.856
R13152 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R13153 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t3 140.163
R13154 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t2 114.031
R13155 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t0 83.3993
R13156 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t4 81.5883
R13157 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R13158 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R13159 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R13160 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R13161 a_44234_6996.t0 a_44234_6996.t1 114.052
R13162 a_28172_6250.n2 a_28172_6250.t2 247.918
R13163 a_28172_6250.n0 a_28172_6250.t1 245.935
R13164 a_28172_6250.n1 a_28172_6250.t3 245.381
R13165 a_28172_6250.n0 a_28172_6250.t4 239.267
R13166 a_28172_6250.t0 a_28172_6250.n2 239.267
R13167 a_28172_6250.n1 a_28172_6250.n0 6.24633
R13168 a_28172_6250.n2 a_28172_6250.n1 0.7755
R13169 a_34186_8950.n0 a_34186_8950.t2 245.316
R13170 a_34186_8950.n0 a_34186_8950.t1 243.361
R13171 a_34186_8950.t0 a_34186_8950.n0 239.308
R13172 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t0 157.346
R13173 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t2 142.179
R13174 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t3 140.314
R13175 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t1 140.065
R13176 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n0 7.42011
R13177 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n2 0.063
R13178 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n1 0.0171667
R13179 a_23583_20174.n0 a_23583_20174.t1 249.335
R13180 a_23583_20174.n1 a_23583_20174.t2 247.23
R13181 a_23583_20174.t0 a_23583_20174.n1 241.299
R13182 a_23583_20174.n0 a_23583_20174.t3 239.248
R13183 a_23583_20174.n1 a_23583_20174.n0 2.10675
R13184 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.t1 239.53
R13185 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.t2 10.533
R13186 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.n0 10.5295
R13187 a_45343_4622.t0 a_45343_4622.t1 60.9236
R13188 a_43240_20238.t0 a_43240_20238.t1 65.941
R13189 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22.t0 247.119
R13190 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22.t2 10.5296
R13191 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22.t1 10.5285
R13192 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22.n0 3.54349
R13193 a_45023_20264.t0 a_45023_20264.t1 49.8467
R13194 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.t1 239.357
R13195 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.n0 10.7707
R13196 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.t2 10.7309
R13197 a_43724_9926.t0 a_43724_9926.t1 55.3905
R13198 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42.t2 249.947
R13199 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42.t0 10.5306
R13200 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42.t1 10.5285
R13201 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42.n0 3.5287
R13202 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32.t2 241.547
R13203 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32.t1 12.1521
R13204 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32.n0 12.0768
R13205 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t2 663.232
R13206 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.n0 10.6713
R13207 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t1 10.5739
R13208 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t2 673.259
R13209 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t1 10.7368
R13210 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t0 10.6531
R13211 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.n0 0.682657
R13212 a_23049_18133.t0 a_23049_18133.n3 242.181
R13213 a_23049_18133.n0 a_23049_18133.t5 240.082
R13214 a_23049_18133.n0 a_23049_18133.t1 239.415
R13215 a_23049_18133.n1 a_23049_18133.t3 239.248
R13216 a_23049_18133.n2 a_23049_18133.t2 239.248
R13217 a_23049_18133.n3 a_23049_18133.t4 239.248
R13218 a_23049_18133.n1 a_23049_18133.n0 3.40883
R13219 a_23049_18133.n3 a_23049_18133.n2 2.93383
R13220 a_23049_18133.n2 a_23049_18133.n1 2.93383
R13221 a_43724_16302.t0 a_43724_16302.t1 55.3905
R13222 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.t2 239.999
R13223 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.t1 10.5782
R13224 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.n0 10.5739
R13225 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.t2 240.44
R13226 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.n0 10.534
R13227 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.t1 10.5285
R13228 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t2 146.001
R13229 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t3 144.221
R13230 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n1 143.886
R13231 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t0 143.494
R13232 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n0 0.7525
R13233 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n1 863.124
R13234 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n0 585
R13235 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t0 495.469
R13236 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t5 217.555
R13237 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t6 217.042
R13238 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t3 216.63
R13239 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t4 212.911
R13240 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t2 212.393
R13241 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t7 208.054
R13242 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t1 141.189
R13243 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t0 140.738
R13244 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n7 30.2547
R13245 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n9 26.7318
R13246 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 14.3755
R13247 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 11.6369
R13248 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n8 11.2109
R13249 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n6 11.1922
R13250 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 10.1408
R13251 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 10.0547
R13252 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n10 8.53383
R13253 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n3 7.94225
R13254 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 6.14988
R13255 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 5.81868
R13256 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 4.80819
R13257 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n5 4.5005
R13258 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n4 3.57742
R13259 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 2.16154
R13260 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n2 0.665435
R13261 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.214442
R13262 a_45343_3530.t0 a_45343_3530.t1 49.8467
R13263 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t2 674.658
R13264 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t0 10.7653
R13265 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t1 10.7376
R13266 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.n0 4.0963
R13267 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t0 673.412
R13268 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t1 10.7203
R13269 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t2 10.6898
R13270 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.n0 3.42178
R13271 a_24411_20174.n0 a_24411_20174.t2 249.518
R13272 a_24411_20174.n1 a_24411_20174.t1 249.325
R13273 a_24411_20174.t0 a_24411_20174.n1 241.115
R13274 a_24411_20174.n0 a_24411_20174.t3 239.431
R13275 a_24411_20174.n1 a_24411_20174.n0 0.19425
R13276 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.t1 241.31
R13277 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.t2 10.5439
R13278 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.n0 10.5295
R13279 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n9 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t13 135.499
R13280 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n10 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t12 135.499
R13281 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t2 134.734
R13282 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t4 134.734
R13283 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t1 134.734
R13284 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n6 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t7 134.734
R13285 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t6 134.734
R13286 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n5 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t3 134.734
R13287 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t5 134.734
R13288 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n3 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t0 134.734
R13289 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n9 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t15 134.715
R13290 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n10 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t14 134.715
R13291 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t10 133.338
R13292 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n12 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t8 132.793
R13293 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t9 58.9067
R13294 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n0 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t11 58.9067
R13295 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n2 15.4672
R13296 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n5 15.4672
R13297 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n11 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 9.85842
R13298 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n12 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n11 8.58003
R13299 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n8 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n7 8.3355
R13300 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n8 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n4 7.15195
R13301 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n9 6.49842
R13302 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n10 6.33383
R13303 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n4 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n3 4.5005
R13304 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n7 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n6 4.5005
R13305 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n0 2.09724
R13306 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n11 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n8 1.70389
R13307 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n12 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n1 0.484196
R13308 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n12 0.0484167
R13309 a_43240_21320.t0 a_43240_21320.t1 65.941
R13310 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t0 272.038
R13311 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t0 258.846
R13312 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t3 230.363
R13313 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n0 201.161
R13314 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t4 158.064
R13315 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n1 155.328
R13316 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n2 29.1319
R13317 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t1 26.5955
R13318 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t2 26.5955
R13319 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n3 23.616
R13320 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 3.76521
R13321 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 3.0725
R13322 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n4 3.03935
R13323 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n5 2.30266
R13324 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.921363
R13325 a_23031_20174.t0 a_23031_20174.n1 250.069
R13326 a_23031_20174.n0 a_23031_20174.t2 249.745
R13327 a_23031_20174.n0 a_23031_20174.t1 240.565
R13328 a_23031_20174.n1 a_23031_20174.t3 239.982
R13329 a_23031_20174.n1 a_23031_20174.n0 0.323417
R13330 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.t2 240.188
R13331 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.n0 10.5827
R13332 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.t1 10.5739
R13333 a_34569_10031.n0 a_34569_10031.t1 240.108
R13334 a_34569_10031.t0 a_34569_10031.n0 239.733
R13335 a_34569_10031.n0 a_34569_10031.t2 238.899
R13336 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t1 227.856
R13337 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n2 152.333
R13338 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t4 140.382
R13339 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t2 114.031
R13340 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t0 83.3993
R13341 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t3 81.5883
R13342 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n3 14.4422
R13343 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n1 7.56882
R13344 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n0 5.08175
R13345 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R13346 a_45023_19712.t0 a_45023_19712.t1 49.8467
R13347 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t2 756.356
R13348 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t1 235.56
R13349 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t0 152.889
R13350 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[3] 14.6392
R13351 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 2.22659
R13352 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_0.Y 1.55202
R13353 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[3] 0.826393
R13354 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t5 753.758
R13355 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.Y 586.745
R13356 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 289.24
R13357 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t3 230.576
R13358 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t4 158.275
R13359 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 153.661
R13360 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 152
R13361 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t1 26.5955
R13362 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t2 24.9236
R13363 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t0 24.9236
R13364 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 23.1774
R13365 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[4] 18.1258
R13366 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.Y 17.9639
R13367 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 10.7516
R13368 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 10.238
R13369 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n6 6.66717
R13370 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[4] 0.7505
R13371 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.t1 680.375
R13372 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.t2 10.7835
R13373 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.n0 10.6741
R13374 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.t1 677.731
R13375 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.n0 10.7394
R13376 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.t2 10.6292
R13377 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t4 241.536
R13378 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n2 195.704
R13379 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t3 169.237
R13380 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n0 152
R13381 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t1 140.53
R13382 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n3 41.8732
R13383 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n1 28.2143
R13384 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t2 26.5955
R13385 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t0 26.5955
R13386 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 16.5652
R13387 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n4 9.03579
R13388 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 1.87783
R13389 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 1.72748
R13390 a_44234_9332.t0 a_44234_9332.t1 114.052
R13391 a_4415_23194.n2 a_4415_23194.t5 160.632
R13392 a_4415_23194.n5 a_4415_23194.t0 151.631
R13393 a_4415_23194.n2 a_4415_23194.t3 134.811
R13394 a_4415_23194.t1 a_4415_23194.n5 134.811
R13395 a_4415_23194.n0 a_4415_23194.t4 16.8154
R13396 a_4415_23194.n1 a_4415_23194.t6 16.8154
R13397 a_4415_23194.n3 a_4415_23194.n1 12.0038
R13398 a_4415_23194.n5 a_4415_23194.n4 6.72342
R13399 a_4415_23194.n4 a_4415_23194.n0 6.5892
R13400 a_4415_23194.n0 a_4415_23194.t7 5.78822
R13401 a_4415_23194.n1 a_4415_23194.t2 5.78822
R13402 a_4415_23194.n4 a_4415_23194.n3 5.66508
R13403 a_4415_23194.n3 a_4415_23194.n2 0.965083
R13404 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36.t2 246.268
R13405 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36.t0 10.5306
R13406 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36.t1 10.5285
R13407 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36.n0 2.15701
R13408 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t3 230.363
R13409 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n0 203.147
R13410 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t4 158.064
R13411 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n1 152
R13412 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t1 140.53
R13413 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n3 34.4304
R13414 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t2 26.5955
R13415 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t0 26.5955
R13416 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n2 24.0657
R13417 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 16.5652
R13418 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n4 9.03579
R13419 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 3.2005
R13420 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 1.72748
R13421 a_22469_18133.t0 a_22469_18133.n3 242.364
R13422 a_22469_18133.n0 a_22469_18133.t3 240.264
R13423 a_22469_18133.n0 a_22469_18133.t5 239.631
R13424 a_22469_18133.n1 a_22469_18133.t2 239.431
R13425 a_22469_18133.n2 a_22469_18133.t1 239.431
R13426 a_22469_18133.n3 a_22469_18133.t4 239.431
R13427 a_22469_18133.n1 a_22469_18133.n0 4.04217
R13428 a_22469_18133.n3 a_22469_18133.n2 2.93383
R13429 a_22469_18133.n2 a_22469_18133.n1 2.93383
R13430 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35.t2 245.728
R13431 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35.t1 10.5752
R13432 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35.t0 10.5739
R13433 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35.n0 1.55257
R13434 a_20547_20174.t0 a_20547_20174.n1 250.803
R13435 a_20547_20174.n0 a_20547_20174.t2 248.238
R13436 a_20547_20174.n1 a_20547_20174.t3 240.714
R13437 a_20547_20174.n0 a_20547_20174.t1 239.833
R13438 a_20547_20174.n1 a_20547_20174.n0 2.56508
R13439 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.n0 240.321
R13440 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.t1 10.7966
R13441 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.t2 10.6741
R13442 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.t2 240.931
R13443 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.t1 13.8869
R13444 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.n0 10.8444
R13445 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.t2 240.24
R13446 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.t1 10.7826
R13447 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.n0 10.6302
R13448 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 593.158
R13449 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 231.554
R13450 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 140.53
R13451 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 26.5955
R13452 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 26.5955
R13453 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 16.5652
R13454 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 9.03579
R13455 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 6.02403
R13456 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 1.72748
R13457 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.t2 240.773
R13458 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.t1 13.9942
R13459 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.n0 11.0596
R13460 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.t2 243.41
R13461 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.n0 10.5372
R13462 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.t1 10.5285
R13463 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t2 673.212
R13464 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t1 10.7631
R13465 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t0 10.7147
R13466 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.n0 2.72674
R13467 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t2 673.273
R13468 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t0 10.7808
R13469 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t1 10.6292
R13470 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.n0 3.43753
R13471 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 593.165
R13472 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 268.077
R13473 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 258.846
R13474 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 237.577
R13475 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 26.5955
R13476 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 26.5955
R13477 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 16.5652
R13478 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 9.03579
R13479 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 8.8386
R13480 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 1.72748
R13481 a_36033_10031.t0 a_36033_10031.n0 241.075
R13482 a_36033_10031.n0 a_36033_10031.t2 239.35
R13483 a_36033_10031.n0 a_36033_10031.t1 238.716
R13484 a_43167_4634.t0 a_43167_4634.t1 49.8467
R13485 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51.t0 245.726
R13486 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51.t1 10.575
R13487 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51.t2 10.5739
R13488 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51.n0 1.5626
R13489 a_14615_13785.t0 a_14615_13785.n0 439.543
R13490 a_14615_13785.n0 a_14615_13785.t1 39.3576
R13491 a_14615_13785.n0 a_14615_13785.t2 39.3576
R13492 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18.t2 238.254
R13493 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18.t1 10.5761
R13494 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18.n0 10.5739
R13495 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19.t2 248.799
R13496 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19.n0 10.6684
R13497 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19.t1 10.5285
R13498 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23.t0 248.075
R13499 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23.t2 10.6701
R13500 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23.t1 10.5739
R13501 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23.n0 4.17455
R13502 a_45023_19988.t0 a_45023_19988.t1 49.8467
R13503 a_20498_8950.n0 a_20498_8950.t1 671.928
R13504 a_20498_8950.n0 a_20498_8950.t2 671.475
R13505 a_20498_8950.t0 a_20498_8950.n0 665.158
R13506 a_15869_6250.n2 a_15869_6250.t3 673.378
R13507 a_15869_6250.n0 a_15869_6250.t2 673.005
R13508 a_15869_6250.n1 a_15869_6250.t1 669.523
R13509 a_15869_6250.n0 a_15869_6250.t4 666.583
R13510 a_15869_6250.t0 a_15869_6250.n2 666.583
R13511 a_15869_6250.n1 a_15869_6250.n0 4.60675
R13512 a_15869_6250.n2 a_15869_6250.n1 1.95467
R13513 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54.t0 246.798
R13514 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54.t2 10.6247
R13515 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54.t1 10.5285
R13516 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54.n0 3.49191
R13517 a_29158_6250.n2 a_29158_6250.t2 248.469
R13518 a_29158_6250.n0 a_29158_6250.t1 246.486
R13519 a_29158_6250.n1 a_29158_6250.t3 244.054
R13520 a_29158_6250.n0 a_29158_6250.t4 239.816
R13521 a_29158_6250.t0 a_29158_6250.n2 239.816
R13522 a_29158_6250.n2 a_29158_6250.n1 5.54425
R13523 a_29158_6250.n1 a_29158_6250.n0 1.47758
R13524 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.t0 249.738
R13525 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.t1 13.5018
R13526 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.t2 10.7924
R13527 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.n0 4.72836
R13528 a_43724_6956.t0 a_43724_6956.t1 55.3905
R13529 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t2 674.658
R13530 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t1 10.7625
R13531 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t0 10.7309
R13532 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.n0 4.09058
R13533 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5.t1 246.63
R13534 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5.t0 10.5795
R13535 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5.t2 10.5739
R13536 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5.n0 2.90483
R13537 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6.t2 248.484
R13538 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6.t0 10.5338
R13539 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6.t1 10.5285
R13540 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6.n0 3.63285
R13541 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t1 675.741
R13542 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t2 10.7126
R13543 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t0 10.6732
R13544 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.n0 2.0546
R13545 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 593.165
R13546 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 268.077
R13547 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 258.846
R13548 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 237.577
R13549 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 26.5955
R13550 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 26.5955
R13551 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 16.5652
R13552 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 9.03579
R13553 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 8.8386
R13554 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 1.72748
R13555 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t1 221.851
R13556 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t3 221.851
R13557 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t4 140.625
R13558 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t5 140.244
R13559 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t7 113.648
R13560 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t6 113.648
R13561 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t0 108.365
R13562 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t2 108.365
R13563 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n5 12.9957
R13564 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n4 1.60385
R13565 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n3 0.557293
R13566 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n1 0.557293
R13567 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n2 0.266714
R13568 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n0 0.063
R13569 DIN6.n1 DIN6.t1 212.081
R13570 DIN6.n0 DIN6.t0 212.081
R13571 DIN6.n2 DIN6.n1 183.185
R13572 DIN6.n1 DIN6.t3 139.78
R13573 DIN6.n0 DIN6.t2 139.78
R13574 DIN6.n1 DIN6.n0 61.346
R13575 DIN6 DIN6.n2 14.2776
R13576 DIN6.n2 DIN6 5.8885
R13577 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t2 672.956
R13578 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t0 10.717
R13579 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t1 10.6712
R13580 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.n0 2.0484
R13581 a_34873_10031.n0 a_34873_10031.t1 240.13
R13582 a_34873_10031.t0 a_34873_10031.n0 239.512
R13583 a_34873_10031.n0 a_34873_10031.t2 238.921
R13584 DIN4.n1 DIN4.t0 212.081
R13585 DIN4.n0 DIN4.t3 212.081
R13586 DIN4.n2 DIN4.n1 183.185
R13587 DIN4.n1 DIN4.t2 139.78
R13588 DIN4.n0 DIN4.t1 139.78
R13589 DIN4.n1 DIN4.n0 61.346
R13590 DIN4 DIN4.n2 14.2776
R13591 DIN4.n2 DIN4 5.8885
R13592 a_43698_15706.n0 a_43698_15706.t1 228.04
R13593 a_43698_15706.n0 a_43698_15706.t2 145.648
R13594 a_43698_15706.t0 a_43698_15706.n0 83.2159
R13595 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t2 667.052
R13596 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.n0 10.6701
R13597 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t1 10.5739
R13598 a_17443_7686.n1 a_17443_7686.t2 672.947
R13599 a_17443_7686.n0 a_17443_7686.t3 671.573
R13600 a_17443_7686.n0 a_17443_7686.t1 666.919
R13601 a_17443_7686.n1 a_17443_7686.t4 666.46
R13602 a_17443_7686.t0 a_17443_7686.n2 666.46
R13603 a_17443_7686.n2 a_17443_7686.n1 6.63383
R13604 a_17443_7686.n2 a_17443_7686.n0 1.84008
R13605 a_44062_20941.t0 a_44062_20941.t1 129.28
R13606 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t0 334.822
R13607 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t3 126.27
R13608 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t4 125.558
R13609 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t2 125.558
R13610 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n1 5.73592
R13611 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n2 5.66196
R13612 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n0 0.713
R13613 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t1 0.197295
R13614 DIN7.n1 DIN7.t0 212.081
R13615 DIN7.n0 DIN7.t3 212.081
R13616 DIN7.n2 DIN7.n1 183.185
R13617 DIN7.n1 DIN7.t2 139.78
R13618 DIN7.n0 DIN7.t1 139.78
R13619 DIN7.n1 DIN7.n0 61.346
R13620 DIN7 DIN7.n2 14.2776
R13621 DIN7.n2 DIN7 5.8885
R13622 a_35177_10031.n0 a_35177_10031.t2 243.633
R13623 a_35177_10031.t0 a_35177_10031.n0 241.625
R13624 a_35177_10031.n0 a_35177_10031.t1 239.267
R13625 a_45023_21412.t0 a_45023_21412.t1 49.8467
R13626 a_17167_7686.n1 a_17167_7686.t2 672.764
R13627 a_17167_7686.n0 a_17167_7686.t3 670.999
R13628 a_17167_7686.n0 a_17167_7686.t1 666.655
R13629 a_17167_7686.n1 a_17167_7686.t4 666.275
R13630 a_17167_7686.t0 a_17167_7686.n2 666.275
R13631 a_17167_7686.n2 a_17167_7686.n1 6.63383
R13632 a_17167_7686.n2 a_17167_7686.n0 2.23175
R13633 a_20222_8950.n0 a_20222_8950.t1 671.744
R13634 a_20222_8950.n0 a_20222_8950.t2 671.292
R13635 a_20222_8950.t0 a_20222_8950.n0 665.34
R13636 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t2 743.367
R13637 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t1 223.315
R13638 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t0 152.889
R13639 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[1] 15.4066
R13640 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n0 12.2462
R13641 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n1 2.22659
R13642 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_1.Y 1.55202
R13643 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[1] 0.84425
R13644 a_15863_13785.n0 a_15863_13785.t2 1266.96
R13645 a_15863_13785.t0 a_15863_13785.n0 65.941
R13646 a_15863_13785.n0 a_15863_13785.t1 65.941
R13647 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19.t1 245.726
R13648 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19.t0 10.6701
R13649 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19.t2 10.5739
R13650 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19.n0 1.51759
R13651 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18.t0 247.037
R13652 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18.t1 10.5307
R13653 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18.t2 10.5285
R13654 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18.n0 0.885467
R13655 a_42724_19156.t0 a_42724_19156.t1 65.941
R13656 a_42982_19156.t0 a_42982_19156.t1 65.941
R13657 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t2 675.77
R13658 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t0 10.7393
R13659 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t1 10.6502
R13660 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.n0 0.682179
R13661 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 593.396
R13662 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 268.077
R13663 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 258.846
R13664 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 231.554
R13665 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 26.5955
R13666 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 26.5955
R13667 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 16.5652
R13668 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 9.03579
R13669 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 8.8386
R13670 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 6.02403
R13671 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 1.72748
R13672 a_44234_12936.t0 a_44234_12936.t1 114.052
R13673 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.t1 239.483
R13674 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.t2 10.7256
R13675 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.n0 10.6908
R13676 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.n1 676.072
R13677 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t3 672.926
R13678 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t2 13.884
R13679 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t1 10.7934
R13680 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.n0 5.03253
R13681 a_44234_11312.t0 a_44234_11312.t1 114.052
R13682 a_43698_10756.t0 a_43698_10756.n0 228.04
R13683 a_43698_10756.n0 a_43698_10756.t2 145.648
R13684 a_43698_10756.n0 a_43698_10756.t1 83.2159
R13685 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.t2 249.738
R13686 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.t1 13.4746
R13687 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.t0 10.7886
R13688 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.n0 4.72836
R13689 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t4 766.463
R13690 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 203.923
R13691 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 101.49
R13692 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t3 26.5955
R13693 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t2 26.5955
R13694 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t1 24.9236
R13695 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t0 24.9236
R13696 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 13.0565
R13697 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 10.7525
R13698 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y 6.6565
R13699 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y 5.04292
R13700 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y 4.3525
R13701 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y 2.5605
R13702 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 1.93989
R13703 a_43724_16856.t0 a_43724_16856.t1 55.3905
R13704 a_43724_10362.t0 a_43724_10362.t1 55.3905
R13705 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t5 739.816
R13706 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t8 230.155
R13707 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t7 230.155
R13708 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 203.923
R13709 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t6 157.856
R13710 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t4 157.856
R13711 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 152
R13712 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 152
R13713 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 101.49
R13714 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t3 26.5955
R13715 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t2 26.5955
R13716 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 25.1816
R13717 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t1 24.9236
R13718 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t0 24.9236
R13719 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[0] 14.1609
R13720 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 13.0565
R13721 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 12.2559
R13722 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 11.0199
R13723 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 10.7525
R13724 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y 6.6565
R13725 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 5.10675
R13726 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y 5.04292
R13727 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y 4.3525
R13728 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y 2.5605
R13729 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.A 2.10199
R13730 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.A 2.10199
R13731 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 1.93989
R13732 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13.t2 676.942
R13733 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13.t1 10.7298
R13734 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13.n0 10.6646
R13735 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t2 668.13
R13736 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t1 12.1225
R13737 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.n0 12.0768
R13738 DIN0.n1 DIN0.t1 212.081
R13739 DIN0.n0 DIN0.t0 212.081
R13740 DIN0.n2 DIN0.n1 183.185
R13741 DIN0.n1 DIN0.t3 139.78
R13742 DIN0.n0 DIN0.t2 139.78
R13743 DIN0.n1 DIN0.n0 61.346
R13744 DIN0 DIN0.n2 14.2776
R13745 DIN0.n2 DIN0 5.8885
R13746 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t1 675.929
R13747 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t2 10.8167
R13748 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t0 10.6741
R13749 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.n0 4.10816
R13750 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t0 676.712
R13751 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t2 10.7718
R13752 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t1 10.6268
R13753 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.n0 3.43316
R13754 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t2 675.904
R13755 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t0 10.7799
R13756 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t1 10.6965
R13757 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.n0 1.35813
R13758 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n1 863.124
R13759 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n0 585
R13760 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t0 495.469
R13761 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t17 217.555
R13762 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t9 217.555
R13763 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t4 217.555
R13764 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t14 216.893
R13765 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t13 216.893
R13766 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t10 216.893
R13767 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t15 216.893
R13768 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t5 216.893
R13769 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t12 216.893
R13770 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t16 216.893
R13771 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t7 216.893
R13772 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t3 216.893
R13773 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t11 216.893
R13774 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t8 216.893
R13775 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t6 212.393
R13776 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t2 212.393
R13777 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t1 141.189
R13778 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t0 140.738
R13779 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n18 71.8985
R13780 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 14.7588
R13781 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 11.6369
R13782 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 10.1408
R13783 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n3 7.94225
R13784 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n19 7.75808
R13785 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 6.59444
R13786 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 6.14988
R13787 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n15 4.5005
R13788 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n17 4.5005
R13789 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 2.16154
R13790 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n16 1.89425
R13791 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n2 0.665435
R13792 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n14 0.663962
R13793 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n13 0.663962
R13794 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n12 0.663962
R13795 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n11 0.663962
R13796 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n10 0.663962
R13797 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n4 0.663962
R13798 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n5 0.663962
R13799 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n6 0.663962
R13800 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n7 0.663962
R13801 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n8 0.663962
R13802 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n9 0.663962
R13803 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.65675
R13804 a_15593_6250.n2 a_15593_6250.t3 673.193
R13805 a_15593_6250.n0 a_15593_6250.t2 672.821
R13806 a_15593_6250.n1 a_15593_6250.t1 670.087
R13807 a_15593_6250.n0 a_15593_6250.t4 666.399
R13808 a_15593_6250.t0 a_15593_6250.n2 666.399
R13809 a_15593_6250.n1 a_15593_6250.n0 4.99842
R13810 a_15593_6250.n2 a_15593_6250.n1 1.563
R13811 DIN3.n1 DIN3.t1 212.081
R13812 DIN3.n0 DIN3.t0 212.081
R13813 DIN3.n2 DIN3.n1 183.185
R13814 DIN3.n1 DIN3.t3 139.78
R13815 DIN3.n0 DIN3.t2 139.78
R13816 DIN3.n1 DIN3.n0 61.346
R13817 DIN3 DIN3.n2 14.3234
R13818 DIN3.n2 DIN3 5.8885
R13819 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t2 667.052
R13820 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.n0 10.6713
R13821 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t1 10.5739
R13822 a_44479_4170.t0 a_44479_4170.t1 49.8467
R13823 a_44479_4254.t0 a_44479_4254.t1 60.9236
R13824 a_44062_18805.t0 a_44062_18805.t1 129.28
R13825 a_44062_20229.t0 a_44062_20229.t1 129.28
R13826 a_43724_7392.t0 a_43724_7392.t1 55.3905
R13827 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 593.158
R13828 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 231.554
R13829 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 140.53
R13830 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 26.5955
R13831 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 26.5955
R13832 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 16.5652
R13833 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 9.03579
R13834 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 6.02403
R13835 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 1.72748
R13836 a_43167_3438.t0 a_43167_3438.t1 49.8467
R13837 a_27896_6250.n2 a_27896_6250.t2 247.736
R13838 a_27896_6250.n0 a_27896_6250.t1 245.752
R13839 a_27896_6250.n1 a_27896_6250.t3 245.172
R13840 a_27896_6250.n0 a_27896_6250.t4 239.083
R13841 a_27896_6250.t0 a_27896_6250.n2 239.083
R13842 a_27896_6250.n1 a_27896_6250.n0 5.85467
R13843 a_27896_6250.n2 a_27896_6250.n1 1.16717
R13844 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35.n0 238.345
R13845 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35.t1 10.7398
R13846 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35.t2 10.6488
R13847 a_43698_6796.n0 a_43698_6796.t1 228.04
R13848 a_43698_6796.n0 a_43698_6796.t2 145.648
R13849 a_43698_6796.t0 a_43698_6796.n0 83.2159
R13850 a_19670_8950.n0 a_19670_8950.t1 671.409
R13851 a_19670_8950.n0 a_19670_8950.t2 670.924
R13852 a_19670_8950.t0 a_19670_8950.n0 665.707
R13853 a_15041_6250.n2 a_15041_6250.t3 672.827
R13854 a_15041_6250.n0 a_15041_6250.t2 672.455
R13855 a_15041_6250.n1 a_15041_6250.t1 671.236
R13856 a_15041_6250.n0 a_15041_6250.t4 666.034
R13857 a_15041_6250.t0 a_15041_6250.n2 666.034
R13858 a_15041_6250.n1 a_15041_6250.n0 5.78175
R13859 a_15041_6250.n2 a_15041_6250.n1 0.779667
R13860 a_15317_6250.n2 a_15317_6250.t3 673.01
R13861 a_15317_6250.n0 a_15317_6250.t2 672.638
R13862 a_15317_6250.n1 a_15317_6250.t1 670.662
R13863 a_15317_6250.n0 a_15317_6250.t4 666.216
R13864 a_15317_6250.t0 a_15317_6250.n2 666.216
R13865 a_15317_6250.n1 a_15317_6250.n0 5.39008
R13866 a_15317_6250.n2 a_15317_6250.n1 1.17133
R13867 a_43724_13332.t0 a_43724_13332.t1 55.3905
R13868 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t0 231.016
R13869 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t1 230.996
R13870 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t3 230.959
R13871 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t2 230.272
R13872 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n0 0.968985
R13873 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n1 0.550258
R13874 a_22755_20174.n0 a_22755_20174.t3 250.435
R13875 a_22755_20174.t0 a_22755_20174.n2 249.549
R13876 a_22755_20174.n0 a_22755_20174.t4 240.347
R13877 a_22755_20174.n2 a_22755_20174.t1 240.2
R13878 a_22755_20174.n1 a_22755_20174.t2 240.2
R13879 a_22755_20174.n2 a_22755_20174.n1 0.633833
R13880 a_22755_20174.n1 a_22755_20174.n0 0.252583
R13881 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.n0 240.804
R13882 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.t2 13.9904
R13883 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.t1 10.8053
R13884 a_16181_7686.n1 a_16181_7686.t2 672.213
R13885 a_16181_7686.n0 a_16181_7686.t3 668.944
R13886 a_16181_7686.n0 a_16181_7686.t1 666.405
R13887 a_16181_7686.n1 a_16181_7686.t4 665.726
R13888 a_16181_7686.t0 a_16181_7686.n2 665.726
R13889 a_16181_7686.n2 a_16181_7686.n1 6.63383
R13890 a_16181_7686.n2 a_16181_7686.n0 3.73592
R13891 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t0 675.533
R13892 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t2 10.7625
R13893 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t1 10.7161
R13894 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.n0 2.72817
R13895 a_42724_19554.t0 a_42724_19554.t1 65.941
R13896 a_42982_19554.t0 a_42982_19554.t1 65.941
R13897 a_43391_3710.t0 a_43391_3710.t1 49.8467
R13898 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t2 675.533
R13899 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t1 10.7636
R13900 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t0 10.7261
R13901 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.n0 2.74248
R13902 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t2 677.236
R13903 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t0 10.7544
R13904 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t1 10.6216
R13905 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.n0 3.42573
R13906 a_42724_20978.t0 a_42724_20978.t1 65.941
R13907 a_42982_20978.t0 a_42982_20978.t1 65.941
R13908 a_31318_7686.n2 a_31318_7686.t2 246.794
R13909 a_31318_7686.n0 a_31318_7686.t1 243.439
R13910 a_31318_7686.n0 a_31318_7686.t3 239.809
R13911 a_31318_7686.n1 a_31318_7686.t4 239.51
R13912 a_31318_7686.t0 a_31318_7686.n2 239.51
R13913 a_31318_7686.n2 a_31318_7686.n1 6.788
R13914 a_31318_7686.n1 a_31318_7686.n0 2.65258
R13915 a_34580_8950.n0 a_34580_8950.t2 245.95
R13916 a_34580_8950.n0 a_34580_8950.t1 244.102
R13917 a_34580_8950.t0 a_34580_8950.n0 238.94
R13918 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.t1 240.298
R13919 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.t2 10.7108
R13920 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.n0 10.687
R13921 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t1 675.975
R13922 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t0 10.7163
R13923 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t2 10.6736
R13924 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.n0 2.05556
R13925 a_44234_15272.t0 a_44234_15272.t1 114.052
R13926 a_15863_13536.t0 a_15863_13536.n0 1266.83
R13927 a_15863_13536.n0 a_15863_13536.t2 65.941
R13928 a_15863_13536.n0 a_15863_13536.t1 65.941
R13929 a_20352_10031.n0 a_20352_10031.t2 668.659
R13930 a_20352_10031.n0 a_20352_10031.t1 668.024
R13931 a_20352_10031.t0 a_20352_10031.n0 665.667
R13932 a_16320_18696.t0 a_16320_18696.n0 671.341
R13933 a_16320_18696.n0 a_16320_18696.t2 666.413
R13934 a_16320_18696.n0 a_16320_18696.t1 665.855
R13935 a_45023_19116.t0 a_45023_19116.t1 49.8467
R13936 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 593.154
R13937 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 268.077
R13938 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 258.846
R13939 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 231.554
R13940 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 26.5955
R13941 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 26.5955
R13942 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 16.5652
R13943 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 9.03579
R13944 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 8.8386
R13945 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 6.02403
R13946 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 1.72748
R13947 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t2 667.057
R13948 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t1 10.6819
R13949 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.n0 10.5739
R13950 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t1 676.005
R13951 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t2 10.7345
R13952 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t0 10.6522
R13953 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.n0 0.683611
R13954 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62.t0 249.178
R13955 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62.t2 10.6247
R13956 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62.t1 10.5285
R13957 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62.n0 0.872789
R13958 a_15905_7686.n1 a_15905_7686.t2 672.03
R13959 a_15905_7686.n0 a_15905_7686.t3 668.37
R13960 a_15905_7686.n0 a_15905_7686.t1 666.942
R13961 a_15905_7686.n1 a_15905_7686.t4 665.543
R13962 a_15905_7686.t0 a_15905_7686.n2 665.543
R13963 a_15905_7686.n2 a_15905_7686.n1 6.63383
R13964 a_15905_7686.n2 a_15905_7686.n0 4.12758
R13965 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t1 676.48
R13966 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t0 10.7836
R13967 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t2 10.6316
R13968 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.n0 3.43753
R13969 a_19772_10031.n0 a_19772_10031.t2 666.712
R13970 a_19772_10031.t0 a_19772_10031.n0 666.096
R13971 a_19772_10031.n0 a_19772_10031.t1 665.505
R13972 a_45023_20540.t0 a_45023_20540.t1 49.8467
R13973 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t2 674.658
R13974 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t1 10.7657
R13975 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t0 10.7357
R13976 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.n0 4.09773
R13977 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17.n0 236.649
R13978 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17.t2 10.6701
R13979 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17.t1 10.5739
R13980 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t2 675.904
R13981 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t1 10.7856
R13982 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t0 10.6951
R13983 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.n0 1.35718
R13984 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t1 227.856
R13985 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n2 152.333
R13986 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t4 140.382
R13987 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t2 114.031
R13988 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t0 83.3993
R13989 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t3 81.5883
R13990 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n3 14.4422
R13991 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n1 7.56882
R13992 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n0 5.08175
R13993 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R13994 a_43724_13886.t0 a_43724_13886.t1 55.3905
R13995 a_45023_18288.t0 a_45023_18288.t1 49.8467
R13996 a_42847_3710.t0 a_42847_3710.t1 41.3705
R13997 a_33910_8950.n0 a_33910_8950.t2 244.909
R13998 a_33910_8950.n0 a_33910_8950.t1 243.178
R13999 a_33910_8950.t0 a_33910_8950.n0 239.489
R14000 a_13779_6250.n2 a_13779_6250.t3 672.093
R14001 a_13779_6250.n0 a_13779_6250.t2 671.721
R14002 a_13779_6250.n1 a_13779_6250.t1 671.35
R14003 a_13779_6250.n0 a_13779_6250.t4 665.299
R14004 a_13779_6250.t0 a_13779_6250.n2 665.299
R14005 a_13779_6250.n2 a_13779_6250.n1 4.60675
R14006 a_13779_6250.n1 a_13779_6250.n0 1.95467
R14007 a_19000_8950.n0 a_19000_8950.t1 670.336
R14008 a_19000_8950.n0 a_19000_8950.t2 670
R14009 a_19000_8950.t0 a_19000_8950.n0 666.258
R14010 a_24209_18133.n0 a_24209_18133.t3 241.857
R14011 a_24209_18133.t0 a_24209_18133.n2 241.815
R14012 a_24209_18133.n0 a_24209_18133.t2 238.881
R14013 a_24209_18133.n1 a_24209_18133.t1 238.881
R14014 a_24209_18133.n2 a_24209_18133.t4 238.881
R14015 a_24209_18133.n2 a_24209_18133.n1 2.93383
R14016 a_24209_18133.n1 a_24209_18133.n0 2.93383
R14017 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.t2 239.869
R14018 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.t1 10.8275
R14019 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.n0 10.677
R14020 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t2 675.814
R14021 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t1 10.7152
R14022 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t0 10.6722
R14023 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.n0 2.05317
R14024 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13.t1 249.321
R14025 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13.t0 10.575
R14026 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13.t2 10.5739
R14027 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13.n0 1.60689
R14028 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14.t2 249.623
R14029 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14.t0 10.5319
R14030 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14.t1 10.5285
R14031 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14.n0 0.915451
R14032 a_42724_18472.t0 a_42724_18472.t1 65.941
R14033 a_42982_18472.t0 a_42982_18472.t1 65.941
R14034 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t1 227.856
R14035 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R14036 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t3 140.163
R14037 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t2 114.031
R14038 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t0 83.3993
R14039 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t4 81.5883
R14040 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R14041 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R14042 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R14043 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R14044 a_44234_7986.t0 a_44234_7986.t1 114.052
R14045 a_14607_6250.n2 a_14607_6250.t3 672.644
R14046 a_14607_6250.n0 a_14607_6250.t2 672.27
R14047 a_14607_6250.n1 a_14607_6250.t1 671.963
R14048 a_14607_6250.n0 a_14607_6250.t4 665.85
R14049 a_14607_6250.t0 a_14607_6250.n2 665.85
R14050 a_14607_6250.n2 a_14607_6250.n1 5.78175
R14051 a_14607_6250.n1 a_14607_6250.n0 0.779667
R14052 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t2 672.309
R14053 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t0 10.7857
R14054 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t1 10.6946
R14055 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.n0 1.3567
R14056 a_44062_22009.t0 a_44062_22009.t1 129.28
R14057 a_45023_18564.t0 a_45023_18564.t1 49.8467
R14058 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t1 676.321
R14059 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t2 13.4994
R14060 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t0 10.7733
R14061 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.n0 4.72836
R14062 a_43724_17292.t0 a_43724_17292.t1 55.3905
R14063 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t2 753.312
R14064 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n0 268.349
R14065 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t0 268.077
R14066 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t1 230.518
R14067 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n1 27.3291
R14068 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[2] 12.4649
R14069 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.Y 11.6875
R14070 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n2 7.23528
R14071 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.Y 5.04292
R14072 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n0 3.68535
R14073 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[2] 0.90675
R14074 a_22479_20174.n0 a_22479_20174.t2 250.619
R14075 a_22479_20174.t0 a_22479_20174.n1 249.733
R14076 a_22479_20174.n0 a_22479_20174.t3 240.531
R14077 a_22479_20174.n1 a_22479_20174.t1 240.016
R14078 a_22479_20174.n1 a_22479_20174.n0 0.885917
R14079 a_43698_16696.t0 a_43698_16696.n0 228.04
R14080 a_43698_16696.n0 a_43698_16696.t2 145.648
R14081 a_43698_16696.n0 a_43698_16696.t1 83.2159
R14082 a_44255_3162.t0 a_44255_3162.t1 49.8467
R14083 a_18008_18696.n1 a_18008_18696.t3 667.399
R14084 a_18008_18696.n0 a_18008_18696.t2 666.116
R14085 a_18008_18696.t0 a_18008_18696.n1 665.615
R14086 a_18008_18696.n0 a_18008_18696.t1 665.484
R14087 a_18008_18696.n1 a_18008_18696.n0 1.39217
R14088 a_44234_7352.t0 a_44234_7352.t1 114.052
R14089 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52.t0 246.18
R14090 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52.t1 10.5296
R14091 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52.t2 10.5285
R14092 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52.n0 2.14387
R14093 a_37410_19098.n1 a_37410_19098.t0 229.328
R14094 a_37410_19098.t1 a_37410_19098.n1 226.986
R14095 a_37410_19098.n0 a_37410_19098.t3 127.692
R14096 a_37410_19098.n1 a_37410_19098.n0 12.484
R14097 a_37410_19098.n0 a_37410_19098.t2 10.584
R14098 a_43240_19156.t0 a_43240_19156.t1 65.941
R14099 a_21099_20174.n0 a_21099_20174.t2 251.536
R14100 a_21099_20174.t0 a_21099_20174.n1 250.017
R14101 a_21099_20174.n0 a_21099_20174.t3 241.447
R14102 a_21099_20174.n1 a_21099_20174.t1 239.1
R14103 a_21099_20174.n1 a_21099_20174.n0 1.51925
R14104 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30.t2 237.898
R14105 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30.n0 10.786
R14106 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30.t1 10.6951
R14107 a_43391_4174.t0 a_43391_4174.t1 49.8467
R14108 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t0 675.904
R14109 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t2 10.7766
R14110 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t1 10.6951
R14111 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.n0 1.35956
R14112 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t2 675.533
R14113 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t1 10.7605
R14114 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t0 10.7175
R14115 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.n0 2.73151
R14116 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48.t1 241.547
R14117 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48.t2 12.1321
R14118 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48.n0 12.0768
R14119 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t1 663.232
R14120 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t2 10.6713
R14121 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.n0 10.5739
R14122 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t1 668.13
R14123 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.n0 12.1402
R14124 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t2 12.0758
R14125 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t2 675.929
R14126 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t0 10.8299
R14127 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t1 10.6741
R14128 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.n0 4.11253
R14129 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29.t1 249.321
R14130 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29.t2 10.6701
R14131 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29.t0 10.5739
R14132 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29.n0 1.54779
R14133 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t2 752.994
R14134 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t1 230.518
R14135 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t0 162.351
R14136 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[4] 26.8833
R14137 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y 11.6875
R14138 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 7.23528
R14139 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y 3.10353
R14140 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 1.93989
R14141 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[4] 0.790679
R14142 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29.t2 238.269
R14143 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29.t1 10.7341
R14144 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29.n0 10.6526
R14145 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16.t1 241.547
R14146 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16.t2 12.2056
R14147 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16.n0 12.0768
R14148 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.t1 239.793
R14149 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.n0 10.7638
R14150 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.t2 10.7314
R14151 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15.t2 240.469
R14152 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15.t1 10.6713
R14153 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15.n0 10.5739
R14154 a_43724_7946.t0 a_43724_7946.t1 55.3905
R14155 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t2 668.13
R14156 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.n0 12.177
R14157 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t1 12.0758
R14158 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t2 676.321
R14159 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t0 13.4542
R14160 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t1 10.7771
R14161 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.n0 4.72836
R14162 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.t2 249.345
R14163 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.t0 10.575
R14164 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.t1 10.5739
R14165 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.n0 4.20348
R14166 a_45343_3894.t0 a_45343_3894.t1 49.8467
R14167 a_45343_3978.t0 a_45343_3978.t1 60.9236
R14168 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63.t1 240.469
R14169 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63.t2 10.6713
R14170 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63.n0 10.5739
R14171 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17.t2 242.349
R14172 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17.n0 10.6929
R14173 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17.t1 10.5285
R14174 a_42724_21662.t0 a_42724_21662.t1 65.941
R14175 a_42982_21662.t0 a_42982_21662.t1 65.941
R14176 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t2 673.212
R14177 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t0 10.7601
R14178 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t1 10.7161
R14179 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.n0 2.72817
R14180 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.t2 668.534
R14181 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.t1 668.481
R14182 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.n1 11.7566
R14183 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.t3 10.6569
R14184 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0.n0 5.86455
R14185 a_43240_19554.t0 a_43240_19554.t1 65.941
R14186 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t2 672.722
R14187 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t1 10.7152
R14188 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t0 10.6722
R14189 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.n0 2.05317
R14190 a_43240_20978.t0 a_43240_20978.t1 65.941
R14191 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t1 673.332
R14192 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t0 10.7393
R14193 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t2 10.6478
R14194 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.n0 0.682179
R14195 a_44234_13926.t0 a_44234_13926.t1 114.052
R14196 a_5111_8388.n2 a_5111_8388.t2 213.52
R14197 a_5111_8388.n1 a_5111_8388.t0 213.52
R14198 a_5111_8388.n1 a_5111_8388.n0 42.5016
R14199 a_5111_8388.n3 a_5111_8388.n2 42.5016
R14200 a_5111_8388.n2 a_5111_8388.n1 11.7539
R14201 a_5111_8388.n0 a_5111_8388.t4 5.77029
R14202 a_5111_8388.n0 a_5111_8388.t1 5.77029
R14203 a_5111_8388.t3 a_5111_8388.n3 5.77029
R14204 a_5111_8388.n3 a_5111_8388.t5 5.77029
R14205 a_44234_12302.t0 a_44234_12302.t1 114.052
R14206 a_43698_11746.t0 a_43698_11746.n0 228.04
R14207 a_43698_11746.n0 a_43698_11746.t2 145.648
R14208 a_43698_11746.n0 a_43698_11746.t1 83.2159
R14209 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.t1 237.625
R14210 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.t0 15.5077
R14211 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.t2 10.6569
R14212 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.n1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.n0 2.49239
R14213 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0.n1 0.252408
R14214 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.n0 240.44
R14215 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.t1 10.7488
R14216 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.t2 10.6292
R14217 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t1 157.49
R14218 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t2 142.079
R14219 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t0 140.304
R14220 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t3 139.327
R14221 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n0 7.54544
R14222 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n1 0.063
R14223 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t1 227.856
R14224 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n2 152.333
R14225 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t3 140.382
R14226 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t2 114.031
R14227 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t0 83.3993
R14228 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t4 81.5883
R14229 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n3 14.4422
R14230 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n1 7.56882
R14231 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n0 5.08175
R14232 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R14233 a_43724_10916.t0 a_43724_10916.t1 55.3905
R14234 a_42724_20580.t0 a_42724_20580.t1 65.941
R14235 a_42982_20580.t0 a_42982_20580.t1 65.941
R14236 a_44479_3530.t0 a_44479_3530.t1 49.8467
R14237 a_45023_21688.t0 a_45023_21688.t1 49.8467
R14238 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t2 663.232
R14239 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t1 10.6701
R14240 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.n0 10.5739
R14241 a_44479_3898.t0 a_44479_3898.t1 49.8467
R14242 a_43240_18472.t0 a_43240_18472.t1 65.941
R14243 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t2 274.793
R14244 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t4 231.017
R14245 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n3 205.28
R14246 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t5 158.716
R14247 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n0 153.347
R14248 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t1 130.49
R14249 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n4 67.4857
R14250 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n2 38.9629
R14251 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t3 26.5955
R14252 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t0 26.5955
R14253 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n1 22.1046
R14254 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 3.81804
R14255 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t2 675.843
R14256 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t1 10.7383
R14257 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t0 10.6488
R14258 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.n0 0.682179
R14259 a_45343_3254.t0 a_45343_3254.t1 49.8467
R14260 a_43724_8382.t0 a_43724_8382.t1 55.3905
R14261 a_44234_16896.t0 a_44234_16896.t1 114.052
R14262 a_44062_19161.t0 a_44062_19161.t1 129.28
R14263 a_43698_7786.n0 a_43698_7786.t1 228.04
R14264 a_43698_7786.n0 a_43698_7786.t2 145.648
R14265 a_43698_7786.t0 a_43698_7786.n0 83.2159
R14266 a_19276_8950.n0 a_19276_8950.t1 670.519
R14267 a_19276_8950.n0 a_19276_8950.t2 670.183
R14268 a_19276_8950.t0 a_19276_8950.n0 666.073
R14269 a_44062_20585.t0 a_44062_20585.t1 129.28
R14270 a_43724_14322.t0 a_43724_14322.t1 55.3905
R14271 a_44234_16262.t0 a_44234_16262.t1 114.052
R14272 ROUT2.n1 ROUT2.t1 134.847
R14273 ROUT2.n2 ROUT2.t3 134.246
R14274 ROUT2.n3 ROUT2 13.0108
R14275 ROUT2.n1 ROUT2.n0 8.36161
R14276 ROUT2.t5 ROUT2.t4 5.8809
R14277 ROUT2.t0 ROUT2.t5 5.0615
R14278 ROUT2.n0 ROUT2.t2 2.9407
R14279 ROUT2.n0 ROUT2.t0 2.9407
R14280 ROUT2.n2 ROUT2.n1 0.601043
R14281 ROUT2.n3 ROUT2.n2 0.271587
R14282 ROUT2 ROUT2.n3 0.023
R14283 a_43994_22522.n0 a_43994_22522.t3 135.572
R14284 a_43994_22522.t1 a_43994_22522.n1 135.572
R14285 a_43994_22522.n1 a_43994_22522.t0 134.246
R14286 a_43994_22522.n0 a_43994_22522.t2 134.246
R14287 a_43994_22522.n1 a_43994_22522.n0 1.1418
R14288 a_15342_18696.t0 a_15342_18696.n0 670.384
R14289 a_15342_18696.n0 a_15342_18696.t1 668.327
R14290 a_15342_18696.n0 a_15342_18696.t2 665.848
R14291 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.t2 675.904
R14292 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.t0 10.7652
R14293 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.t1 10.6927
R14294 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.n0 1.36672
R14295 a_44255_4530.t0 a_44255_4530.t1 49.8467
R14296 a_43724_11352.t0 a_43724_11352.t1 55.3905
R14297 a_43724_14876.t0 a_43724_14876.t1 55.3905
R14298 a_43391_3242.t0 a_43391_3242.t1 49.8467
R14299 a_44234_8976.t0 a_44234_8976.t1 114.052
R14300 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47.t2 240.469
R14301 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47.n0 10.6713
R14302 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47.t1 10.5739
R14303 a_42724_18814.t0 a_42724_18814.t1 65.941
R14304 a_42982_18814.t0 a_42982_18814.t1 65.941
R14305 a_43240_21662.t0 a_43240_21662.t1 65.941
R14306 a_44234_8342.t0 a_44234_8342.t1 114.052
R14307 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4.t1 239.142
R14308 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4.n0 10.5871
R14309 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4.t2 10.5739
R14310 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46.t2 249.239
R14311 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46.t1 10.6247
R14312 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46.t0 10.5295
R14313 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46.n0 0.872789
R14314 a_44234_10956.t0 a_44234_10956.t1 114.052
R14315 a_44255_4078.t0 a_44255_4078.t1 49.8467
R14316 a_44255_4162.t0 a_44255_4162.t1 60.9236
R14317 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61.t0 249.321
R14318 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61.t1 10.6701
R14319 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61.t2 10.5739
R14320 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61.n0 1.53658
R14321 a_44255_4446.t0 a_44255_4446.t1 49.8467
R14322 a_42724_20238.t0 a_42724_20238.t1 65.941
R14323 a_42982_20238.t0 a_42982_20238.t1 65.941
R14324 a_43391_3158.t0 a_43391_3158.t1 49.8467
R14325 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.t2 242.369
R14326 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.n0 10.5394
R14327 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.t1 10.5285
R14328 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20.t2 239.094
R14329 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20.n0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20.t1 10.6701
R14330 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20.t0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20.n0 10.5739
R14331 a_44062_19873.t0 a_44062_19873.t1 129.28
R14332 a_44234_13292.t0 a_44234_13292.t1 114.052
R14333 a_43724_11906.t0 a_43724_11906.t1 55.3905
R14334 a_42724_22004.t0 a_42724_22004.t1 65.941
R14335 a_44062_21297.t0 a_44062_21297.t1 129.28
R14336 a_42724_18130.t0 a_42724_18130.t1 65.941
R14337 a_42724_19896.t0 a_42724_19896.t1 65.941
C0 a_1896_16243# a_2678_16243# 0.02127f
C1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_39883_19479# 0.02736f
C2 a_44067_22496# ROUT2 0.08397f
C3 a_1896_20320# a_2678_20320# 0.02127f
C4 a_6445_14150# VDDH 0.49013f
C5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 0.15598f
C6 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_6445_15057# 0.04959f
C7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.04405f
C8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 VDDH 0.15179f
C9 a_2300_14353# VDDH 0.53441f
C10 a_1636_13708# a_1636_13352# 0.02286f
C11 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.06345f
C12 a_7625_12507# a_8173_12507# 0.0103f
C13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.64353f
C14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.13343f
C15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 1.47954f
C16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.02493f
C17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.02615f
C18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 1.3157f
C19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.02715f
C20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.21475f
C21 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.06917f
C22 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.05396f
C23 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.02122f
C24 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1636_14353# 0.03043f
C25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.14826f
C26 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 0.03135f
C27 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_final_switch_0.VOUT[4] 5.50358f
C28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.1245f
C29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.04779f
C30 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C31 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] DIN7 0.0349f
C32 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.05883f
C33 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.01796f
C34 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_5897_14150# 0.04959f
C35 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[2] 0.39626f
C36 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.06351f
C37 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 VDDH 0.10984f
C38 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.06278f
C39 DIN1 DIN2 0.33f
C40 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.18203f
C41 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.01389f
C42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 VDDH 0.14262f
C43 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 8.23983f
C44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 VDDH 0.47118f
C45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02077f
C46 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_2678_19053# 0.01343f
C47 a_11629_14150# VOUT 0.0409f
C48 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.19453f
C49 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 1.36438f
C50 a_39861_21457# VDDH 0.40618f
C51 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.01469f
C52 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.16626f
C53 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.VH3 0.05944f
C54 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_final_switch_0.VOUT[3] 0.05206f
C55 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 1.04282f
C56 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD 0.21766f
C57 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_final_switch_0.VOUT[4] 0.06373f
C58 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.055f
C59 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] VDD 3.68198f
C60 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_2678_12504# 0.04249f
C61 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.03552f
C62 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] VDDH 0.85743f
C63 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_final_switch_0.VOUT[1] 5.80043f
C64 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.40887f
C65 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.15968f
C66 a_11081_13005# a_11629_13005# 0.0103f
C67 a_39861_22496# VDDH 1.43189f
C68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN a_5642_8388# 0.01976f
C69 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.98493f
C70 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 1.15703f
C71 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.05159f
C72 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.12314f
C73 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD 0.23151f
C74 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 1.34913f
C75 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.09546f
C76 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_2678_20320# 0.05095f
C77 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.06812f
C78 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y VDD 0.49613f
C79 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.04851f
C80 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B VOUT 0.65147f
C81 top_DAC_0/top_final_switch_0.VOUT[1] VOUT 6.36642f
C82 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09271f
C83 VDD DIN5 0.67364f
C84 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD a_4717_15057# 0.01033f
C85 a_7625_14150# a_8173_14150# 0.0237f
C86 VDDH ROUT2 9.92565f
C87 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 0.04732f
C88 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 0.02163f
C89 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.10072f
C90 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 0.02198f
C91 a_4978_8388# a_5642_8388# 0.02543f
C92 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_7625_15057# 0.04959f
C93 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.08581f
C94 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 0.15788f
C95 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09013f
C96 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.0436f
C97 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.15473f
C98 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.01165f
C99 a_6445_12507# VOUT 0.03463f
C100 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.0436f
C101 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.0203f
C102 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.06158f
C103 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.03366f
C104 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 VDDH 0.16165f
C105 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C VDD 0.26024f
C106 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] VDDH 2.1111f
C107 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_39861_21457# 0.06598f
C108 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_final_switch_0.VOUT[1] 0.01647f
C109 top_DAC_0/top_final_switch_0.VOUT[3] a_11629_14150# 0.01208f
C110 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 1.57341f
C111 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 VOUT 0.13144f
C112 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.VL3 0.17935f
C113 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.77374f
C114 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 0.16476f
C115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.02121f
C116 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 3.28115f
C117 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.02001f
C118 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.43094f
C119 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 ROUT2 0.01358f
C120 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.05843f
C121 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09914f
C122 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.15972f
C123 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.0961f
C124 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 1.37492f
C125 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 VDDH 0.10118f
C126 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A VDD 0.32055f
C127 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 0.05551f
C128 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD 0.2275f
C129 a_2678_19053# VDDH 0.72825f
C130 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.04937f
C131 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.05186f
C132 top_DAC_0/top_rseg_n_dcell_0.SH[1] VDDH 1.78593f
C133 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.0119f
C134 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 1.24994f
C135 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_final_switch_0.VOUT[2] 0.01655f
C136 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 1.24591f
C137 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.05518f
C138 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.0239f
C139 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_11629_14150# 0.04994f
C140 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_final_switch_0.VOUT[3] 0.10582f
C141 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.05833f
C142 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.05877f
C143 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV ROUT2 0.25958f
C144 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1896_19053# 0.02486f
C145 a_8173_15057# VDDH 0.49886f
C146 top_DAC_0/top_final_switch_0.VOUT[0] a_6445_14150# 0.01199f
C147 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 0.09136f
C148 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.04834f
C149 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.049f
C150 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.07383f
C151 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.15469f
C152 a_2300_13708# a_2300_13352# 0.02286f
C153 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.17416f
C154 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.19079f
C155 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_final_switch_0.VOUT[2] 0.01823f
C156 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.0514f
C157 a_11629_12507# VOUT 0.03463f
C158 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.15992f
C159 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 1.1572f
C160 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] VDDH 0.88599f
C161 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.04929f
C162 a_44737_4828# VDD 0.02571f
C163 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 0.21283f
C164 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.06069f
C165 a_6445_14150# VOUT 0.0409f
C166 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.45991f
C167 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.VH2 0.05786f
C168 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.01132f
C169 VDD DIN6 0.70858f
C170 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04064f
C171 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.98671f
C172 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.05253f
C173 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 1.81035f
C174 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_2678_17510# 0.06357f
C175 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.0505f
C176 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04064f
C177 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.VH2 0.20766f
C178 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.5556f
C179 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.02079f
C180 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_final_switch_0.VOUT[1] 0.20373f
C181 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.20079f
C182 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.17825f
C183 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 0.01835f
C184 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.01887f
C185 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 0.04824f
C186 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 0.04313f
C187 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.06115f
C188 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.09544f
C189 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 0.48841f
C190 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.03009f
C191 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.11542f
C192 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1896_12504# 0.06294f
C193 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.VL3 0.06414f
C194 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.16951f
C195 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 VDDH 4.40766f
C196 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 0.57553f
C197 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.09312f
C198 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] VDDH 2.21503f
C199 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_20320# 0.06368f
C200 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A 0.90356f
C201 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.01068f
C202 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.12876f
C203 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 0.02615f
C204 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 0.02493f
C205 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 1.33973f
C206 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] VDDH 1.29039f
C207 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04362f
C208 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_4717_13005# 0.02092f
C209 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 VDDH 0.04651f
C210 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.34747f
C211 a_5897_15057# a_6445_15057# 0.0237f
C212 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_2678_11886# 0.04314f
C213 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 VDDH 1.16961f
C214 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 8.15945f
C215 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.03773f
C216 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 1.39623f
C217 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.05175f
C218 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VDDH 2.32693f
C219 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.04626f
C220 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.02139f
C221 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.0921f
C222 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.02163f
C223 a_44067_22496# VDDH 1.22217f
C224 DIN2 DIN3 0.33146f
C225 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.04736f
C226 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 1.34563f
C227 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.09544f
C228 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 VDDH 3.10831f
C229 a_1896_17510# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.06357f
C230 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.07752f
C231 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_2678_19053# 0.05235f
C232 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.02121f
C233 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.05719f
C234 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 3.18174f
C235 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 2.15109f
C236 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 VDDH 1.32603f
C237 a_9353_15057# VDDH 0.49783f
C238 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 1.97317f
C239 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.04843f
C240 a_36813_19760# a_36813_19462# 0.015f
C241 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 0.09964f
C242 a_1896_22970# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.06357f
C243 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 0.01142f
C244 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y VDD 0.33964f
C245 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 1.40678f
C246 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.12293f
C247 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.09992f
C248 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 2.90337f
C249 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.04875f
C250 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 0.28615f
C251 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 1.15763f
C252 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.21387f
C253 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 0.65201f
C254 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.17741f
C255 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 0.11135f
C256 a_11629_15057# top_DAC_0/top_final_switch_0.VOUT[4] 0.03029f
C257 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.09997f
C258 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_9901_13005# 0.0208f
C259 VDD DIN7 0.71581f
C260 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.07563f
C261 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.17417f
C262 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.02595f
C263 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD 0.21631f
C264 top_DAC_0/top_rseg_n_dcell_0.SH[3] VDDH 1.2895f
C265 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.05175f
C266 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 0.04684f
C267 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_6445_14150# 0.04994f
C268 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.03344f
C269 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 VDDH 0.14057f
C270 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 0.02106f
C271 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.09513f
C272 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 VDDH 0.15152f
C273 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.VL2 0.09426f
C274 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_2678_21703# 0.13435f
C275 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 3.48836f
C276 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.4572f
C277 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.06132f
C278 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.6765f
C279 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 1.16389f
C280 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.02213f
C281 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04066f
C282 top_DAC_0/top_rseg_n_dcell_0.VH2 VDDH 0.20437f
C283 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.05322f
C284 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.06276f
C285 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 1.79255f
C286 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.08855f
C287 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.24261f
C288 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 0.0658f
C289 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.VL2 0.06485f
C290 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 VDDH 7.284f
C291 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.44826f
C292 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B VDD 0.25715f
C293 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.09198f
C294 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.24881f
C295 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_9353_12507# 0.0208f
C296 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.0977f
C297 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.11523f
C298 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.05175f
C299 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.02611f
C300 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 1.34056f
C301 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.02537f
C302 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1896_17510# 0.06525f
C303 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 14.0478f
C304 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.01812f
C305 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 0.20729f
C306 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 0.0119f
C307 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 2.89925f
C308 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 0.06043f
C309 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_1896_21703# 0.06357f
C310 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 0.08427f
C311 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 2.07729f
C312 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.062f
C313 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 VDDH 0.14904f
C314 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.05882f
C315 top_DAC_0/top_final_switch_0.VOUT[4] a_11629_13005# 0.02842f
C316 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.01148f
C317 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.1111f
C318 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 0.0954f
C319 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 1.31906f
C320 a_1896_20320# VDDH 0.72706f
C321 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.04939f
C322 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.08478f
C323 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.1675f
C324 a_8173_15057# VOUT 0.01454f
C325 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD a_6445_15057# 0.01033f
C326 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] DIN7 0.01582f
C327 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.26736f
C328 a_5642_11461# a_5642_10963# 0.015f
C329 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.17828f
C330 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 1.45197f
C331 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.25426f
C332 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.10421f
C333 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.05223f
C334 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.08294f
C335 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.11848f
C336 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.04843f
C337 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.60845f
C338 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.05177f
C339 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 VDDH 2.20196f
C340 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.02015f
C341 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04363f
C342 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_final_switch_0.VOUT[4] 0.03109f
C343 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.09515f
C344 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.04736f
C345 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD a_8173_15057# 0.01033f
C346 top_DAC_0/top_final_switch_0.VOUT[4] a_12809_15057# 0.03952f
C347 VDD DIN8 0.72319f
C348 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.VS4 0.03139f
C349 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.18775f
C350 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.09076f
C351 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.02488f
C352 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 17.4806f
C353 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_5897_13005# 0.0208f
C354 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A VDDH 0.90751f
C355 VDD ROUT1 0.68441f
C356 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 VOUT 0.17766f
C357 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 0.87032f
C358 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_final_switch_0.VOUT[0] 0.20436f
C359 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH 17.253f
C360 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_45343_4828# 0.01719f
C361 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09344f
C362 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.06177f
C363 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 0.42912f
C364 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 14.96f
C365 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.87726f
C366 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.07232f
C367 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 1.7882f
C368 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 1.24741f
C369 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.84443f
C370 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 0.02575f
C371 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.14095f
C372 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 17.3231f
C373 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 VDDH 0.15933f
C374 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.VL2 0.11724f
C375 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD a_9901_15057# 0.01035f
C376 top_DAC_0/top_final_switch_0.VOUT[1] a_6445_13005# 0.02851f
C377 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 1.05222f
C378 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.VH3 1.53928f
C379 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD a_5897_15057# 0.01037f
C380 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.12764f
C381 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.26572f
C382 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 1.8611f
C383 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.06127f
C384 top_DAC_0/top_final_switch_0.VOUT[2] a_9901_15057# 0.01175f
C385 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.98866f
C386 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_12504# 0.05618f
C387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT 2.66242f
C388 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_38584_20389# 0.02882f
C389 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 1.19048f
C390 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[2] 0.59509f
C391 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.18445f
C392 a_9353_14150# VDDH 0.49013f
C393 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 0.02541f
C394 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 0.0266f
C395 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 1.34685f
C396 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.30079f
C397 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 VDDH 25.2932f
C398 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.08546f
C399 a_1896_21703# VDDH 0.73997f
C400 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.21776f
C401 a_37595_19760# a_37595_19462# 0.015f
C402 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05675f
C403 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.09505f
C404 a_1636_15118# a_2300_15118# 0.01589f
C405 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 0.29715f
C406 DIN3 DIN4 0.3362f
C407 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.04039f
C408 a_9353_13005# VOUT 0.02203f
C409 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.27678f
C410 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.06065f
C411 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.VS1 0.04711f
C412 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.49342f
C413 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.01687f
C414 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.11409f
C415 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.05759f
C416 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.61579f
C417 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.07707f
C418 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_1896_20320# 0.03145f
C419 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 4.13148f
C420 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 1.2875f
C421 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.09535f
C422 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.04858f
C423 a_9353_15057# VOUT 0.04641f
C424 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD a_7625_15057# 0.01033f
C425 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 0.02015f
C426 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_11081_13005# 0.0208f
C427 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.54094f
C428 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] DIN8 0.17935f
C429 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.07853f
C430 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04068f
C431 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.30168f
C432 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 VDDH 1.23475f
C433 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.11775f
C434 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.05178f
C435 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 1.30528f
C436 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 1.45085f
C437 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.09522f
C438 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_final_switch_0.VOUT[0] 0.01053f
C439 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 3.83937f
C440 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.15222f
C441 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 VDDH 0.04533f
C442 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.04851f
C443 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD a_9353_15057# 0.01034f
C444 VDD DIN9 0.75623f
C445 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.11848f
C446 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.09146f
C447 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 1.94253f
C448 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.11409f
C449 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] VDDH 0.18887f
C450 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.21309f
C451 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 1.27501f
C452 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04366f
C453 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_4978_9535# 0.11619f
C454 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_final_switch_0.VOUT[3] 0.20319f
C455 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.VH2 0.47348f
C456 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.30645f
C457 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.05434f
C458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_final_switch_0.VOUT[4] 0.5995f
C459 top_DAC_0/top_final_switch_0.VOUT[0] VDDH 1.7051f
C460 a_1896_22970# a_2678_22970# 0.02127f
C461 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 VOUT 0.13389f
C462 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.28212f
C463 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.13121f
C464 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.04792f
C465 top_DAC_0/top_final_switch_0.VOUT[4] a_12809_13005# 0.03376f
C466 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 0.39192f
C467 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 0.05585f
C468 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 1.789f
C469 a_4978_9535# VDDH 0.73032f
C470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD a_11081_15057# 0.01033f
C471 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.06231f
C472 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_final_switch_0.VOUT[1] 0.01878f
C473 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.VL2 0.05628f
C474 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 1.3467f
C475 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 0.10095f
C476 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.10297f
C477 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] VDDH 1.26896f
C478 VDDH VOUT 8.72574f
C479 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.06351f
C480 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 VDDH 0.08462f
C481 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD 0.2275f
C482 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.14576f
C483 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 0.09468f
C484 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.13341f
C485 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 1.73459f
C486 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.4235f
C487 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.06152f
C488 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 1.31964f
C489 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.04789f
C490 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 0.69962f
C491 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.05177f
C492 a_38584_20665# a_38584_20389# 0.02286f
C493 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] VDD 1.60464f
C494 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.05177f
C495 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 2.46853f
C496 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.05653f
C497 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 1.45233f
C498 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C499 top_DAC_0/top_final_switch_0.VOUT[4] a_12809_14150# 0.01964f
C500 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.06598f
C501 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.06661f
C502 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05322f
C503 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.09358f
C504 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.VL3 0.1844f
C505 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.02015f
C506 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_39883_19854# 0.02806f
C507 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VDDH 0.63882f
C508 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.10024f
C509 a_6445_15057# top_DAC_0/top_final_switch_0.VOUT[1] 0.03029f
C510 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD 0.23023f
C511 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 0.05743f
C512 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.04969f
C513 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_final_switch_0.VOUT[3] 0.01337f
C514 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax VDDH 4.75556f
C515 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.18677f
C516 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 1.44458f
C517 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04071f
C518 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 3.81788f
C519 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.01833f
C520 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 16.2949f
C521 top_DAC_0/top_final_switch_0.VOUT[1] a_7625_13005# 0.03215f
C522 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.15103f
C523 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_1896_20320# 0.06418f
C524 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.30111f
C525 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] VDDH 0.01105f
C526 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.11409f
C527 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.VS4 0.01859f
C528 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.VS4 0.0322f
C529 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.03007f
C530 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 0.01088f
C531 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_4717_12507# 0.02171f
C532 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.06256f
C533 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.11409f
C534 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.02207f
C535 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 0.79254f
C536 top_DAC_0/top_final_switch_0.VOUT[3] VDDH 1.66679f
C537 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 VDDH 0.14089f
C538 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.06788f
C539 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_1896_10974# 0.03761f
C540 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.13753f
C541 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 VDDH 0.15149f
C542 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_final_switch_0.VOUT[0] 0.0151f
C543 a_4717_15057# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C544 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.6218f
C545 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 1.48f
C546 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.02665f
C547 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.02537f
C548 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.10472f
C549 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 0.21461f
C550 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 1.27914f
C551 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 0.02715f
C552 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 VDDH 3.66239f
C553 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.06295f
C554 a_9353_12507# VOUT 0.04471f
C555 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_2678_17510# 0.0506f
C556 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 0.16205f
C557 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 0.06082f
C558 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04368f
C559 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.16457f
C560 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 10.4407f
C561 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.1481f
C562 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.09163f
C563 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.29277f
C564 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 1.78725f
C565 a_9353_14150# VOUT 0.06741f
C566 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 VOUT 0.03859f
C567 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.48051f
C568 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 1.57333f
C569 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 16.1091f
C570 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 1.32352f
C571 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.05362f
C572 a_2678_17510# VDDH 0.72716f
C573 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 9.03926f
C574 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH 1.85588f
C575 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.26998f
C576 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.06101f
C577 a_1896_10974# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.02981f
C578 DIN4 DIN5 0.34355f
C579 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.66352f
C580 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.11848f
C581 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.05806f
C582 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 0.03142f
C583 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.09784f
C584 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.15777f
C585 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.20454f
C586 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04695f
C587 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.19835f
C588 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.04859f
C589 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_9901_12507# 0.02171f
C590 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04845f
C591 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.05179f
C592 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.5492f
C593 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09325f
C594 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04841f
C595 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.21128f
C596 top_DAC_0/top_final_switch_0.VOUT[1] a_7625_15057# 0.03805f
C597 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 0.02015f
C598 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.38434f
C599 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_5642_9535# 0.01613f
C600 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.05175f
C601 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.01136f
C602 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 VDDH 0.10974f
C603 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 0.48684f
C604 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_1896_21703# 0.0991f
C605 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05891f
C606 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.VL3 0.06329f
C607 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN a_5642_11461# 0.01003f
C608 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.12689f
C609 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.19158f
C610 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 1.32046f
C611 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.09546f
C612 top_DAC_0/top_final_switch_0.VOUT[4] a_12809_12507# 0.01061f
C613 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.1675f
C614 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 0.11835f
C615 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 1.41253f
C616 a_5642_9535# VDDH 0.79462f
C617 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 3.7974f
C618 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C619 top_DAC_0/top_final_switch_0.VOUT[0] VOUT 6.7893f
C620 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.11127f
C621 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.VS1 0.27984f
C622 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_final_switch_0.VOUT[3] 0.01093f
C623 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.05359f
C624 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04075f
C625 a_9901_14150# VDDH 0.49013f
C626 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_9901_15057# 0.04959f
C627 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.17853f
C628 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.0184f
C629 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 0.08857f
C630 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.1676f
C631 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.28795f
C632 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44471_4828# 0.01759f
C633 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 1.25122f
C634 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.VH2 1.1774f
C635 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 15.7968f
C636 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.09106f
C637 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC VDDH 1.19654f
C638 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 VDDH 1.31557f
C639 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 0.18469f
C640 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.73748f
C641 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 1.5609f
C642 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_1896_10356# 0.02965f
C643 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_37022_20295# 0.01181f
C644 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.06101f
C645 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_9353_14150# 0.04959f
C646 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.02113f
C647 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[4] 0.31502f
C648 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.20712f
C649 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC ROUT2 0.01108f
C650 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] VDDH 0.01046f
C651 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 0.0944f
C652 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.56698f
C653 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.04791f
C654 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] VDDH 1.39235f
C655 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09038f
C656 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.VL2 0.57437f
C657 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.VH2 0.06502f
C658 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 0.63647f
C659 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.48886f
C660 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.32927f
C661 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.01651f
C662 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.05884f
C663 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.05183f
C664 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.33061f
C665 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VOUT 0.67332f
C666 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 1.21733f
C667 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.0119f
C668 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04805f
C669 top_DAC_0/top_final_switch_0.VOUT[1] a_7625_12507# 0.01061f
C670 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.10324f
C671 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 0.03202f
C672 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.12875f
C673 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_final_switch_0.VOUT[1] 0.01299f
C674 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A VDD 0.33616f
C675 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.05983f
C676 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.15447f
C677 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.50346f
C678 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.11848f
C679 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax VOUT 0.0675f
C680 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.05996f
C681 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_final_switch_0.VOUT[3] 0.43345f
C682 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 0.02015f
C683 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] VDDH 2.01688f
C684 a_1636_14353# a_2300_14353# 0.01589f
C685 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04841f
C686 a_7625_13005# a_8173_13005# 0.0103f
C687 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.01149f
C688 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 14.4869f
C689 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.05175f
C690 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_2678_16243# 0.0585f
C691 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.48595f
C692 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.14299f
C693 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B VDD 0.36582f
C694 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 VDDH 0.04638f
C695 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.01806f
C696 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.04736f
C697 top_DAC_0/top_final_switch_0.VOUT[3] VOUT 6.36704f
C698 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_final_switch_0.VOUT[2] 0.01317f
C699 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.01854f
C700 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 1.81409f
C701 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 3.76093f
C702 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.05244f
C703 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.01649f
C704 a_9353_14150# a_9901_14150# 0.0237f
C705 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_final_switch_0.VOUT[2] 0.01082f
C706 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.1308f
C707 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 0.54952f
C708 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.11021f
C709 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.09f
C710 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_11081_15057# 0.04959f
C711 a_2678_16243# VDDH 0.72648f
C712 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.58792f
C713 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.VH2 0.31328f
C714 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.11771f
C715 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.20355f
C716 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.VH3 2.98928f
C717 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.03011f
C718 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.02136f
C719 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.05169f
C720 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 1.22792f
C721 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1896_16243# 0.0747f
C722 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.18985f
C723 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.15123f
C724 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 0.13531f
C725 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 0.30567f
C726 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.02254f
C727 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.19295f
C728 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.04788f
C729 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 0.02199f
C730 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_final_switch_0.VOUT[3] 0.01325f
C731 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 1.2479f
C732 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 VDDH 3.72704f
C733 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.VH2 0.05155f
C734 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 VOUT 0.02759f
C735 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.43649f
C736 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT 3.98706f
C737 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.14754f
C738 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.06718f
C739 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] VDDH 1.30585f
C740 top_DAC_0/top_final_switch_0.VOUT[1] a_7625_14150# 0.01864f
C741 VDD ROUT2 0.6068f
C742 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_5642_8388# 0.10623f
C743 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_1636_13708# 0.02725f
C744 a_4717_14150# VDDH 0.48125f
C745 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.VS4 0.03086f
C746 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.05596f
C747 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.02352f
C748 a_9353_12507# a_9901_12507# 0.0103f
C749 DIN5 DIN6 0.36448f
C750 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.VL2 0.05973f
C751 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.10895f
C752 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.VL2 0.18856f
C753 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.0686f
C754 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.18545f
C755 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 0.03915f
C756 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.10293f
C757 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 0.59845f
C758 a_5642_8388# VDDH 0.72861f
C759 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] VDDH 1.54852f
C760 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_final_switch_0.VOUT[4] 0.01346f
C761 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.04329f
C762 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.01212f
C763 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 VDDH 0.20568f
C764 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_1896_12504# 0.01649f
C765 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.96812f
C766 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_final_switch_0.VOUT[4] 0.11637f
C767 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 2.15145f
C768 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 1.97214f
C769 a_11629_15057# VDDH 0.49751f
C770 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.42123f
C771 a_4978_9535# a_5642_9535# 0.02543f
C772 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.05183f
C773 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.17921f
C774 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.07123f
C775 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[1] 0.39674f
C776 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_17510# 0.06384f
C777 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.05177f
C778 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.09624f
C779 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_final_switch_0.VOUT[4] 0.03086f
C780 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 1.73155f
C781 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.VS4 1.61787f
C782 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.01138f
C783 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 0.31595f
C784 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.02821f
C785 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.11848f
C786 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 15.8859f
C787 a_4717_12507# VOUT 0.039f
C788 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.03652f
C789 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.08314f
C790 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.0483f
C791 a_9901_14150# VOUT 0.0409f
C792 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 0.02121f
C793 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.02873f
C794 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.01647f
C795 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.30067f
C796 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_final_switch_0.VOUT[3] 0.20445f
C797 a_45015_4828# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.02202f
C798 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 VDDH 0.14301f
C799 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.02204f
C800 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 VDDH 0.41945f
C801 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 0.09131f
C802 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.01814f
C803 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.06721f
C804 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 17.3168f
C805 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.0759f
C806 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.63972f
C807 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.05213f
C808 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.02116f
C809 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.08304f
C810 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.VH3 0.26823f
C811 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 VDDH 3.49358f
C812 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.13238f
C813 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 0.11409f
C814 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.18515f
C815 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 1.19856f
C816 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.01172f
C817 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.11409f
C818 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.09704f
C819 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04845f
C820 a_7625_15057# a_8173_15057# 0.0237f
C821 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.56233f
C822 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.0517f
C823 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.VL2 5.30487f
C824 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_38617_19854# 0.01035f
C825 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 1.88113f
C826 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.0119f
C827 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 2.09546f
C828 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.08427f
C829 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 0.15587f
C830 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_5897_15057# 0.04959f
C831 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 1.97838f
C832 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.22399f
C833 a_1636_15118# VDDH 0.554f
C834 a_9901_12507# VOUT 0.03463f
C835 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.05185f
C836 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 0.0191f
C837 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 2.89603f
C838 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_2678_20320# 0.05719f
C839 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.04747f
C840 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.0119f
C841 top_DAC_0/top_rseg_n_dcell_0.VL2 VDDH 0.14809f
C842 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.04842f
C843 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09312f
C844 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.61294f
C845 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 3.39716f
C846 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 2.6115f
C847 a_12809_15057# VDDH 0.48955f
C848 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 VDDH 0.11006f
C849 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.04811f
C850 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.578f
C851 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.02015f
C852 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH 4.26993f
C853 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.33336f
C854 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.02214f
C855 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 1.73307f
C856 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.06066f
C857 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.18941f
C858 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.2455f
C859 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 11.41f
C860 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.1866f
C861 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.05518f
C862 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.11409f
C863 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.12577f
C864 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.60657f
C865 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_9901_14150# 0.04994f
C866 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_final_switch_0.VOUT[2] 5.5062f
C867 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.01643f
C868 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_1636_13352# 0.02725f
C869 a_6445_15057# VDDH 0.49751f
C870 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.31886f
C871 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 1.85017f
C872 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 0.09357f
C873 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 5.80789f
C874 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_final_switch_0.VOUT[1] 0.01731f
C875 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] DIN8 0.01582f
C876 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.VH3 0.05427f
C877 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.05329f
C878 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.20774f
C879 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.03404f
C880 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] VDD 1.24016f
C881 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 17.4112f
C882 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.05999f
C883 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.50988f
C884 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 1.16723f
C885 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_1896_11886# 0.02524f
C886 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.04843f
C887 a_4717_14150# VOUT 0.05095f
C888 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.01753f
C889 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.04843f
C890 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 VDDH 0.0402f
C891 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_16243# 0.07145f
C892 DIN6 DIN7 0.33364f
C893 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.0636f
C894 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 1.97694f
C895 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.VL3 0.68768f
C896 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09024f
C897 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.09063f
C898 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 0.02715f
C899 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.21492f
C900 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 1.36638f
C901 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.59731f
C902 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.05765f
C903 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04846f
C904 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.38958f
C905 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.05174f
C906 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 4.12073f
C907 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 0.07007f
C908 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.12623f
C909 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx a_2678_10974# 0.02385f
C910 a_11629_15057# VOUT 0.01454f
C911 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.01718f
C912 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 0.61284f
C913 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.02948f
C914 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_8173_13005# 0.0208f
C915 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.98866f
C916 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 0.0119f
C917 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.97868f
C918 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.33091f
C919 a_1896_19053# a_2678_19053# 0.02127f
C920 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 0.15742f
C921 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.04946f
C922 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 9.22813f
C923 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.70899f
C924 VDDH VDD 5.24685f
C925 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH 2.43082f
C926 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.08957f
C927 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.43454f
C928 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y VDD 0.28031f
C929 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 VDDH 0.04651f
C930 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 16.6023f
C931 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 1.72824f
C932 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 0.36625f
C933 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.01131f
C934 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.04975f
C935 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.18005f
C936 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.1029f
C937 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 1.93547f
C938 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.22605f
C939 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_7625_12507# 0.0208f
C940 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD 0.23151f
C941 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.06201f
C942 top_DAC_0/top_final_switch_0.VOUT[1] a_8173_14150# 0.01201f
C943 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_37737_19479# 0.02737f
C944 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 2.2876f
C945 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.09759f
C946 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.06145f
C947 a_7625_15057# VDDH 0.49751f
C948 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.26895f
C949 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.05025f
C950 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.09117f
C951 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 0.60003f
C952 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.05769f
C953 a_1636_14353# VDDH 0.53376f
C954 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_final_switch_0.VOUT[4] 0.04554f
C955 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] DIN9 0.17935f
C956 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.12411f
C957 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.06095f
C958 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.5188f
C959 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.02726f
C960 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.06862f
C961 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.03375f
C962 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 1.33058f
C963 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.10107f
C964 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_2678_19053# 0.0593f
C965 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_2300_15118# 0.04824f
C966 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.0494f
C967 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A VDDH 0.90617f
C968 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.08819f
C969 top_DAC_0/top_final_switch_0.VOUT[3] a_11629_15057# 0.01175f
C970 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_final_switch_0.VOUT[0] 0.05663f
C971 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 0.03397f
C972 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 0.02726f
C973 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.0484f
C974 a_12809_14150# VDDH 0.48022f
C975 a_1636_15118# VOUT 0.01189f
C976 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[4] 0.47259f
C977 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_4717_14150# 0.05017f
C978 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.31218f
C979 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.04529f
C980 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.53884f
C981 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.04843f
C982 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 17.1095f
C983 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 1.97444f
C984 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.VS1 0.10469f
C985 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] VDDH 0.01032f
C986 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.21426f
C987 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.02715f
C988 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.02163f
C989 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 1.34308f
C990 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.VL2 0.12688f
C991 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 VDDH 0.0707f
C992 a_12809_15057# VOUT 0.04557f
C993 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 VDDH 0.20563f
C994 a_41907_22057# VDDH 0.31401f
C995 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_12809_12507# 0.01625f
C996 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_4978_11461# 0.06246f
C997 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.17102f
C998 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.44932f
C999 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04847f
C1000 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 11.5953f
C1001 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 0.0119f
C1002 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_1896_12504# 0.02948f
C1003 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.26638f
C1004 top_DAC_0/top_final_switch_0.VOUT[0] a_6445_15057# 0.01175f
C1005 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.12526f
C1006 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.09548f
C1007 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.VH2 0.05868f
C1008 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.01814f
C1009 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.12526f
C1010 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.03535f
C1011 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.18751f
C1012 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.05681f
C1013 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 0.16919f
C1014 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 10.3151f
C1015 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04903f
C1016 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.20199f
C1017 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.09809f
C1018 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.VS1 0.06092f
C1019 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 5.06241f
C1020 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C1021 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 15.5261f
C1022 top_DAC_0/top_final_switch_0.VOUT[2] a_8173_13005# 0.02847f
C1023 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 0.43907f
C1024 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 1.72759f
C1025 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 0.21361f
C1026 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 0.02715f
C1027 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04786f
C1028 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 1.3734f
C1029 a_6445_15057# VOUT 0.01454f
C1030 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.1322f
C1031 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.29779f
C1032 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD VDDH 1.18085f
C1033 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 VDDH 0.20664f
C1034 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 12.9813f
C1035 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 0.1869f
C1036 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04882f
C1037 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_38584_20665# 0.01092f
C1038 a_5642_9535# a_5642_8388# 0.015f
C1039 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.58839f
C1040 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] VDDH 2.61713f
C1041 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.07846f
C1042 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09789f
C1043 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 13.196f
C1044 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.57403f
C1045 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.05777f
C1046 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 10.3939f
C1047 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 0.55355f
C1048 a_7625_13005# VOUT 0.02203f
C1049 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] VDD 1.57937f
C1050 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_final_switch_0.VOUT[3] 0.01843f
C1051 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_5642_10963# 0.01106f
C1052 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_2678_10974# 0.02444f
C1053 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.13739f
C1054 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_41907_22057# 0.02974f
C1055 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 0.64599f
C1056 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_9353_13005# 0.0208f
C1057 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.0979f
C1058 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.0259f
C1059 VDDH DIN0 0.4291f
C1060 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 1.33533f
C1061 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.04787f
C1062 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.02766f
C1063 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.03392f
C1064 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] VDD 0.48049f
C1065 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 17.1369f
C1066 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 VDDH 1.7572f
C1067 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 0.02042f
C1068 DIN7 DIN8 0.33719f
C1069 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.1304f
C1070 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.09239f
C1071 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.20364f
C1072 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD 0.21864f
C1073 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.06751f
C1074 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 1.9603f
C1075 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.07143f
C1076 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.12599f
C1077 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 1.31057f
C1078 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 0.21425f
C1079 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 0.02715f
C1080 a_1896_19053# VDDH 0.722f
C1081 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.09256f
C1082 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.09577f
C1083 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y VDD 0.41365f
C1084 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.09114f
C1085 a_8173_15057# top_DAC_0/top_final_switch_0.VOUT[2] 0.03029f
C1086 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.25378f
C1087 a_7625_14150# VDDH 0.49013f
C1088 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.33109f
C1089 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 VDDH 0.10926f
C1090 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VOUT 0.61926f
C1091 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[1] 0.59493f
C1092 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.1529f
C1093 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.07088f
C1094 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.0119f
C1095 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 1.21429f
C1096 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 2.8803f
C1097 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.08251f
C1098 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.80349f
C1099 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 0.0953f
C1100 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 1.28515f
C1101 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.VS4 0.04912f
C1102 a_12809_13005# VOUT 0.02119f
C1103 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 VDDH 0.09915f
C1104 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C1105 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.VS1 0.04547f
C1106 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.63053f
C1107 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 17.3348f
C1108 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.36098f
C1109 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 0.69015f
C1110 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.0673f
C1111 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_2300_14353# 0.04784f
C1112 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.VH2 0.05944f
C1113 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.VS4 0.01837f
C1114 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.01617f
C1115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A VDDH 0.90804f
C1116 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.01844f
C1117 a_7625_15057# VOUT 0.04641f
C1118 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.72782f
C1119 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] VDDH 0.98177f
C1120 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.0485f
C1121 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.63136f
C1122 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.13332f
C1123 a_1636_14353# VOUT 0.02722f
C1124 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05095f
C1125 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 1.57251f
C1126 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 4.1684f
C1127 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.20918f
C1128 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.22509f
C1129 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.1906f
C1130 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 0.25566f
C1131 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.01812f
C1132 a_4978_11461# a_4978_10963# 0.015f
C1133 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.02834f
C1134 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 1.24832f
C1135 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.11409f
C1136 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VDDH 2.24695f
C1137 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.13705f
C1138 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05297f
C1139 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.05838f
C1140 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 0.54188f
C1141 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.23045f
C1142 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.05383f
C1143 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.35307f
C1144 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.55369f
C1145 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.07189f
C1146 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.02024f
C1147 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] VDDH 1.54537f
C1148 a_12809_14150# VOUT 0.06888f
C1149 a_40525_21457# VDDH 0.35437f
C1150 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.VS4 0.36163f
C1151 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.04942f
C1152 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 0.01397f
C1153 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] VDD 1.81308f
C1154 VDDH DIN1 0.42749f
C1155 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.20641f
C1156 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.VH3 0.05787f
C1157 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04948f
C1158 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_1896_11886# 0.02948f
C1159 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.05173f
C1160 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 0.02839f
C1161 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 0.03446f
C1162 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_final_switch_0.VOUT[2] 0.20339f
C1163 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.09294f
C1164 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 VDDH 0.0686f
C1165 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 VDDH 0.22406f
C1166 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_final_switch_0.VOUT[3] 0.01676f
C1167 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.20862f
C1168 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.08824f
C1169 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.02186f
C1170 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.01649f
C1171 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.09596f
C1172 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.0119f
C1173 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 1.18866f
C1174 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.03135f
C1175 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C1176 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_1896_19053# 0.03145f
C1177 top_DAC_0/top_final_switch_0.VOUT[2] a_9353_13005# 0.03212f
C1178 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.06438f
C1179 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 3.73465f
C1180 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 1.27692f
C1181 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.02715f
C1182 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.2143f
C1183 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 0.02197f
C1184 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 0.05305f
C1185 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.30168f
C1186 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.02047f
C1187 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_final_switch_0.VOUT[0] 0.59734f
C1188 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.VL2 0.56064f
C1189 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.04984f
C1190 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.03108f
C1191 top_DAC_0/top_final_switch_0.VOUT[2] a_9353_15057# 0.03805f
C1192 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.09973f
C1193 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 14.8638f
C1194 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 VDDH 6.21616f
C1195 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 0.55111f
C1196 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.08714f
C1197 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.10418f
C1198 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 1.22987f
C1199 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.96629f
C1200 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 VDDH 0.04942f
C1201 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.0152f
C1202 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.18654f
C1203 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.07012f
C1204 a_7625_12507# VOUT 0.04471f
C1205 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 VDDH 0.11672f
C1206 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 0.06072f
C1207 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 0.1877f
C1208 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD VOUT 0.61932f
C1209 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.09312f
C1210 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.0857f
C1211 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 3.3366f
C1212 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 1.83395f
C1213 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.02167f
C1214 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.05244f
C1215 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_2678_10356# 0.02628f
C1216 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 ROUT2 0.0484f
C1217 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_40525_21457# 0.0755f
C1218 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.VL2 0.05912f
C1219 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.69498f
C1220 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.10358f
C1221 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.06657f
C1222 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.1324f
C1223 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 16.2094f
C1224 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.28898f
C1225 a_1896_17510# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 0.03145f
C1226 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.55748f
C1227 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_final_switch_0.VOUT[2] 0.01423f
C1228 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.15063f
C1229 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 0.52521f
C1230 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.08546f
C1231 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 3.55677f
C1232 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.80785f
C1233 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 1.48649f
C1234 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.04851f
C1235 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.78185f
C1236 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.07481f
C1237 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.02218f
C1238 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.02156f
C1239 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.04751f
C1240 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.16418f
C1241 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 0.1499f
C1242 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.03879f
C1243 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 0.50407f
C1244 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 0.0555f
C1245 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 1.22509f
C1246 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.VH2 0.95191f
C1247 a_1896_17510# VDDH 0.722f
C1248 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.55643f
C1249 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.VS4 0.74491f
C1250 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.09522f
C1251 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.01346f
C1252 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.0486f
C1253 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_8173_12507# 0.02171f
C1254 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.VS4 0.01859f
C1255 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 0.16949f
C1256 VDDH DIN2 0.42749f
C1257 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.09326f
C1258 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_12809_14150# 0.04134f
C1259 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VDDH 1.06161f
C1260 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.13195f
C1261 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.15602f
C1262 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_2678_19053# 0.06357f
C1263 top_DAC_0/top_final_switch_0.VOUT[2] VDDH 1.65987f
C1264 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.13293f
C1265 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.12781f
C1266 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 VDDH 1.62525f
C1267 DIN8 DIN9 0.33674f
C1268 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_2678_22970# 0.07653f
C1269 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV VDDH 1.06415f
C1270 a_12809_12507# VOUT 0.04641f
C1271 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C1272 top_DAC_0/top_rseg_n_dcell_0.VH3 VDDH 0.46642f
C1273 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.0151f
C1274 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 VDDH 0.07f
C1275 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.VL2 0.39896f
C1276 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 VDDH 0.20535f
C1277 a_45015_4828# VDD 0.03791f
C1278 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 2.15445f
C1279 a_7625_14150# VOUT 0.06741f
C1280 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 1.9819f
C1281 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 0.02194f
C1282 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.05318f
C1283 a_1636_13708# VOUT 0.0165f
C1284 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_1896_16243# 0.08441f
C1285 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.06147f
C1286 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC a_38584_20665# 0.02697f
C1287 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.11409f
C1288 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 0.05667f
C1289 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.19276f
C1290 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.0942f
C1291 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] VDD 2.59466f
C1292 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.VL2 0.05356f
C1293 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.10201f
C1294 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[0] 0.40016f
C1295 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 1.26125f
C1296 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.04856f
C1297 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 0.71512f
C1298 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.02197f
C1299 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.0921f
C1300 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.05322f
C1301 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_1896_19053# 0.13749f
C1302 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 0.06038f
C1303 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_final_switch_0.VOUT[4] 0.02878f
C1304 a_11081_14150# a_11629_14150# 0.0237f
C1305 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 0.24855f
C1306 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] DIN8 0.0349f
C1307 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.96636f
C1308 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.35945f
C1309 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_5642_10963# 0.0541f
C1310 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.04992f
C1311 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT 21.3105f
C1312 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 VDDH 2.32429f
C1313 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.12455f
C1314 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C1315 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 17.6537f
C1316 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.04794f
C1317 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04799f
C1318 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09785f
C1319 a_39861_22057# VDDH 0.2924f
C1320 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 18.3073f
C1321 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 VDDH 0.15493f
C1322 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 2.73645f
C1323 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04799f
C1324 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 1.14685f
C1325 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 0.11409f
C1326 top_DAC_0/top_final_switch_0.VOUT[2] a_9353_12507# 0.01061f
C1327 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A 0.01383f
C1328 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 VDDH 0.11236f
C1329 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.54398f
C1330 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 1.73519f
C1331 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 1.88678f
C1332 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.VL3 0.62483f
C1333 VDDH DIN3 0.42749f
C1334 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 1.2633f
C1335 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.11902f
C1336 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 VDDH 0.02285f
C1337 top_DAC_0/top_final_switch_0.VOUT[2] a_9353_14150# 0.01867f
C1338 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] a_45015_4828# 0.02963f
C1339 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.04852f
C1340 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 1.78008f
C1341 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.0119f
C1342 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.05086f
C1343 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.2656f
C1344 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 2.14311f
C1345 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.08427f
C1346 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_final_switch_0.VOUT[2] 0.01031f
C1347 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_39768_20665# 0.03153f
C1348 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_8173_15057# 0.04959f
C1349 a_8173_14150# VDDH 0.49013f
C1350 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx VDDH 0.39611f
C1351 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.VS1 2.74289f
C1352 a_2678_22970# VDDH 0.77537f
C1353 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 1.13576f
C1354 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.7893f
C1355 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.06435f
C1356 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 1.3535f
C1357 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 3.15778f
C1358 a_5897_12507# a_6445_12507# 0.0103f
C1359 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.06701f
C1360 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.11409f
C1361 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 0.06065f
C1362 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] VDD 1.73139f
C1363 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.20093f
C1364 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx a_2678_11886# 0.0175f
C1365 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.17964f
C1366 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.47f
C1367 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.05544f
C1368 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 0.05302f
C1369 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 0.02197f
C1370 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_7625_14150# 0.04959f
C1371 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 VDDH 0.56552f
C1372 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[3] 0.39596f
C1373 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.04809f
C1374 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.5508f
C1375 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09787f
C1376 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.02015f
C1377 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.04787f
C1378 a_39861_22057# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.03219f
C1379 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.46871f
C1380 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.1019f
C1381 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 0.03958f
C1382 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 1.40088f
C1383 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.03966f
C1384 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.15269f
C1385 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_final_switch_0.VOUT[4] 0.19335f
C1386 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 0.0421f
C1387 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 0.69233f
C1388 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.48636f
C1389 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.25263f
C1390 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_final_switch_0.VOUT[2] 0.43345f
C1391 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 1.85343f
C1392 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.09478f
C1393 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.33918f
C1394 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.10422f
C1395 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD a_11629_15057# 0.01033f
C1396 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_2678_21703# 0.01199f
C1397 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.61765f
C1398 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.0591f
C1399 a_4717_15057# VDDH 0.49013f
C1400 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.11409f
C1401 a_9353_13005# a_9901_13005# 0.0103f
C1402 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.VS1 0.07771f
C1403 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.04328f
C1404 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.09934f
C1405 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 0.0119f
C1406 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.02181f
C1407 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 1.24381f
C1408 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_final_switch_0.VOUT[0] 0.01446f
C1409 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.04324f
C1410 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VOUT 0.62599f
C1411 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A VDDH 3.88898f
C1412 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A VDD 0.35622f
C1413 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 11.8244f
C1414 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_final_switch_0.VOUT[1] 0.59768f
C1415 top_DAC_0/top_final_switch_0.VOUT[2] VOUT 6.36553f
C1416 VDDH DIN4 0.42749f
C1417 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04799f
C1418 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.04862f
C1419 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_final_switch_0.VOUT[1] 0.03452f
C1420 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.VL3 0.05812f
C1421 a_9353_15057# a_9901_15057# 0.0237f
C1422 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 1.73225f
C1423 a_1636_13352# VOUT 0.01053f
C1424 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 1.18645f
C1425 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 1.77943f
C1426 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.13628f
C1427 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 VDDH 2.01261f
C1428 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_9353_15057# 0.04959f
C1429 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04811f
C1430 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.03991f
C1431 a_1896_20320# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A 0.07342f
C1432 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 0.17836f
C1433 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 VDDH 0.0706f
C1434 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.05183f
C1435 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 VDDH 0.21415f
C1436 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.10302f
C1437 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.33687f
C1438 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.05772f
C1439 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.57187f
C1440 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.13425f
C1441 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_2678_11886# 0.02366f
C1442 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 4.16288f
C1443 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.0315f
C1444 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.07459f
C1445 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.44293f
C1446 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.VH2 0.06354f
C1447 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_1896_17510# 0.01034f
C1448 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.02948f
C1449 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_final_switch_0.VOUT[2] 0.66459f
C1450 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B VDD 0.25878f
C1451 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.06054f
C1452 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.16544f
C1453 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_38617_19854# 0.02826f
C1454 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.94034f
C1455 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.57206f
C1456 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 0.04904f
C1457 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 0.01848f
C1458 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 1.95031f
C1459 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.65418f
C1460 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 1.27264f
C1461 a_11081_12507# a_11629_12507# 0.0103f
C1462 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 3.83598f
C1463 a_1896_22970# VDDH 0.74102f
C1464 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.02308f
C1465 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.VS4 0.06264f
C1466 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.10009f
C1467 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 VDDH 2.92054f
C1468 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.06891f
C1469 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.18998f
C1470 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 0.10426f
C1471 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_final_switch_0.VOUT[3] 0.5979f
C1472 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.05516f
C1473 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.10104f
C1474 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.12584f
C1475 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_final_switch_0.VOUT[4] 0.11625f
C1476 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.18669f
C1477 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_final_switch_0.VOUT[3] 5.48581f
C1478 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] VDDH 0.01029f
C1479 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_1896_11886# 0.02366f
C1480 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.19149f
C1481 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.09855f
C1482 a_9901_15057# VDDH 0.49792f
C1483 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD a_12809_15057# 0.01033f
C1484 a_2678_21703# VDDH 0.75803f
C1485 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH 1.86798f
C1486 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 VDDH 0.36689f
C1487 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_final_switch_0.VOUT[3] 0.02123f
C1488 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.04797f
C1489 a_1636_15118# a_1636_14353# 0.02286f
C1490 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.48603f
C1491 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B VDD 0.29366f
C1492 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.06107f
C1493 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.03419f
C1494 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.02748f
C1495 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.06886f
C1496 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 1.21986f
C1497 a_8173_12507# VOUT 0.03463f
C1498 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.0119f
C1499 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.10119f
C1500 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 1.3027f
C1501 a_1896_17510# a_2678_17510# 0.02127f
C1502 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 15.2414f
C1503 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04402f
C1504 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A 0.3799f
C1505 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.05186f
C1506 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.10026f
C1507 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 3.4847f
C1508 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.05995f
C1509 a_8173_14150# VOUT 0.0409f
C1510 VDDH DIN5 0.42749f
C1511 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.16197f
C1512 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04361f
C1513 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.12637f
C1514 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx VOUT 0.20902f
C1515 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.19372f
C1516 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.96691f
C1517 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.0433f
C1518 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.09248f
C1519 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.18597f
C1520 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_final_switch_0.VOUT[2] 0.204f
C1521 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 1.73509f
C1522 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.04477f
C1523 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.17902f
C1524 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.20703f
C1525 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 5.28584f
C1526 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 VDDH 0.06984f
C1527 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.05167f
C1528 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 VDDH 0.49734f
C1529 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.01826f
C1530 a_5897_14150# a_6445_14150# 0.0237f
C1531 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.01429f
C1532 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.22726f
C1533 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 0.26016f
C1534 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD 0.21864f
C1535 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 4.05624f
C1536 a_4717_15057# top_DAC_0/top_final_switch_0.VOUT[0] 0.03029f
C1537 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_22970# 0.03145f
C1538 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.33598f
C1539 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.48656f
C1540 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.62948f
C1541 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.10492f
C1542 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 1.89956f
C1543 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.08493f
C1544 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04806f
C1545 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.10242f
C1546 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.66863f
C1547 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 0.04346f
C1548 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.02523f
C1549 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.02615f
C1550 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.09461f
C1551 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 1.47977f
C1552 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.07187f
C1553 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.21451f
C1554 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.02715f
C1555 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 1.34745f
C1556 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.VS4 0.03261f
C1557 top_DAC_0/top_final_switch_0.VOUT[2] a_9901_14150# 0.01204f
C1558 top_DAC_0/top_final_switch_0.VOUT[0] a_4717_13005# 0.02832f
C1559 a_4717_15057# VOUT 0.0236f
C1560 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC a_39768_20665# 0.01079f
C1561 a_11081_15057# VDDH 0.49886f
C1562 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.10032f
C1563 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 4.37057f
C1564 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.17853f
C1565 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] ROUT2 0.01445f
C1566 a_1896_21703# a_2678_21703# 0.02127f
C1567 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.05973f
C1568 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04066f
C1569 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] ROUT2 0.02421f
C1570 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.07155f
C1571 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.09591f
C1572 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A VOUT 0.95598f
C1573 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.10584f
C1574 a_4717_13005# VOUT 0.0131f
C1575 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 0.0119f
C1576 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 1.19056f
C1577 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 2.49981f
C1578 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 VDDH 0.41311f
C1579 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 VDDH 0.11272f
C1580 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.VS4 0.06204f
C1581 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_2678_10974# 0.04394f
C1582 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.VL2 0.06058f
C1583 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 0.05308f
C1584 VDDH DIN6 0.42765f
C1585 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.0203f
C1586 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 1.3376f
C1587 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.01056f
C1588 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.05518f
C1589 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_6445_13005# 0.0208f
C1590 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_37804_20713# 0.0211f
C1591 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.93455f
C1592 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.096f
C1593 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.0497f
C1594 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_8173_14150# 0.04994f
C1595 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 17.0519f
C1596 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 1.23034f
C1597 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.05001f
C1598 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.09116f
C1599 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 1.73087f
C1600 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.0532f
C1601 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.01904f
C1602 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 1.63811f
C1603 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.05244f
C1604 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.09271f
C1605 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.03409f
C1606 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.07652f
C1607 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04706f
C1608 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.02906f
C1609 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.08193f
C1610 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.08272f
C1611 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 1.37192f
C1612 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.05433f
C1613 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 0.09544f
C1614 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A 4.38923f
C1615 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_5897_12507# 0.0208f
C1616 top_DAC_0/top_rseg_n_dcell_0.VS4 VDDH 0.47346f
C1617 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.03386f
C1618 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] VDD 1.04528f
C1619 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.26339f
C1620 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.04783f
C1621 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.59483f
C1622 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.4374f
C1623 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.07818f
C1624 a_2300_15118# a_2300_14353# 0.02286f
C1625 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 0.3076f
C1626 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.59336f
C1627 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.VH3 0.06987f
C1628 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.04329f
C1629 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_1896_16243# 0.0335f
C1630 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.08427f
C1631 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 1.916f
C1632 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD 0.21618f
C1633 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] VDD 1.96314f
C1634 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 0.13356f
C1635 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.VS1 0.05653f
C1636 a_9901_15057# VOUT 0.01454f
C1637 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD 0.2275f
C1638 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_11629_13005# 0.0208f
C1639 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.10038f
C1640 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.8597f
C1641 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.85676f
C1642 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT 26.2719f
C1643 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 1.57642f
C1644 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04807f
C1645 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.05224f
C1646 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.11409f
C1647 a_1896_16243# VDDH 0.72203f
C1648 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.0583f
C1649 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.15973f
C1650 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.45968f
C1651 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 0.17986f
C1652 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.VS1 0.07695f
C1653 a_1896_22970# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 0.09901f
C1654 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.15057f
C1655 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.29614f
C1656 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.05188f
C1657 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] ROUT2 0.0162f
C1658 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.16758f
C1659 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 1.15809f
C1660 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 0.0119f
C1661 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.30979f
C1662 VDDH DIN7 0.42767f
C1663 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_11081_12507# 0.0208f
C1664 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.05451f
C1665 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.98976f
C1666 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 0.01611f
C1667 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.03532f
C1668 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] a_45343_4828# 0.01631f
C1669 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.15088f
C1670 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH 3.43289f
C1671 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.55413f
C1672 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 VDDH 0.07006f
C1673 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.03532f
C1674 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.20881f
C1675 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.19454f
C1676 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 VDDH 0.21507f
C1677 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.61039f
C1678 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04891f
C1679 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.03788f
C1680 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.06014f
C1681 a_5897_15057# VDDH 0.49886f
C1682 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.SH[2] 19.0673f
C1683 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.11989f
C1684 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.VL2 0.06145f
C1685 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.05872f
C1686 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_21703# 0.03151f
C1687 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.01646f
C1688 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 1.64648f
C1689 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.05244f
C1690 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 1.15198f
C1691 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_final_switch_0.VOUT[3] 0.17157f
C1692 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 0.09809f
C1693 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 1.34945f
C1694 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.01851f
C1695 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.72578f
C1696 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.20262f
C1697 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.VL3 0.06558f
C1698 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.07353f
C1699 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.06102f
C1700 top_DAC_0/top_final_switch_0.VOUT[3] a_9901_13005# 0.02844f
C1701 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.158f
C1702 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_2678_10356# 0.02366f
C1703 a_4978_8388# VDDH 0.79433f
C1704 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 0.06214f
C1705 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.09644f
C1706 top_DAC_0/top_final_switch_0.VOUT[0] a_5897_13005# 0.03196f
C1707 a_9901_15057# top_DAC_0/top_final_switch_0.VOUT[3] 0.03029f
C1708 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.VH3 0.05157f
C1709 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44737_4828# 0.02083f
C1710 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.2177f
C1711 VDD DIN0 0.71624f
C1712 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.06117f
C1713 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC a_39768_20389# 0.02668f
C1714 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[3] 0.59534f
C1715 a_11081_14150# VDDH 0.49013f
C1716 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.05244f
C1717 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 1.79741f
C1718 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.5557f
C1719 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 0.09994f
C1720 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 VOUT 0.75441f
C1721 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44737_4828# 0.04364f
C1722 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_rseg_n_dcell_0.VS1 0.0444f
C1723 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.03137f
C1724 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 0.55841f
C1725 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.12773f
C1726 a_5897_13005# VOUT 0.02204f
C1727 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 1.94958f
C1728 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 0.08427f
C1729 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.11848f
C1730 a_11081_15057# VOUT 0.04641f
C1731 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.19767f
C1732 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_2678_10356# 0.04179f
C1733 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.VS4 0.03256f
C1734 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.03391f
C1735 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.VS1 0.06127f
C1736 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_7625_13005# 0.0208f
C1737 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.0433f
C1738 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx a_2678_16243# 0.08404f
C1739 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 VDDH 0.04526f
C1740 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.15598f
C1741 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 11.1111f
C1742 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 VDDH 0.33228f
C1743 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 0.04864f
C1744 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 0.60342f
C1745 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.35106f
C1746 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.12736f
C1747 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.04929f
C1748 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.22369f
C1749 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.10571f
C1750 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.13214f
C1751 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.02163f
C1752 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.02218f
C1753 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.04735f
C1754 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04809f
C1755 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 1.19314f
C1756 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.11409f
C1757 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C VDD 0.33516f
C1758 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.02213f
C1759 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.VH2 0.07957f
C1760 VDDH DIN8 0.4277f
C1761 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.20205f
C1762 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.17101f
C1763 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 2.66628f
C1764 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.05552f
C1765 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.VS4 0.01859f
C1766 VDDH ROUT1 29.7603f
C1767 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_final_switch_0.VOUT[4] 0.07919f
C1768 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.VH2 0.05876f
C1769 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.07524f
C1770 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 1.96808f
C1771 a_37595_19462# a_37737_19479# 0.04234f
C1772 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.03534f
C1773 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 1.68068f
C1774 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.05244f
C1775 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 17.521f
C1776 a_11081_13005# VOUT 0.02203f
C1777 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 VDDH 0.07378f
C1778 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] VDDH 1.07221f
C1779 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.09502f
C1780 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 0.09454f
C1781 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.05769f
C1782 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 1.32022f
C1783 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.09811f
C1784 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.05628f
C1785 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] VDDH 0.99488f
C1786 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04883f
C1787 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 2.1375f
C1788 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_final_switch_0.VOUT[2] 0.01788f
C1789 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09746f
C1790 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.04978f
C1791 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_12809_13005# 0.01625f
C1792 top_DAC_0/top_final_switch_0.VOUT[3] a_11081_15057# 0.03805f
C1793 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD VDDH 0.74385f
C1794 VDD DIN1 0.66672f
C1795 top_DAC_0/top_rseg_n_dcell_0.VL3 VDDH 0.57817f
C1796 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.VL2 0.34015f
C1797 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.05086f
C1798 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] DIN6 0.03492f
C1799 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.SH[3] 16.9983f
C1800 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.69667f
C1801 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.02197f
C1802 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.13238f
C1803 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 2.17542f
C1804 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.05305f
C1805 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 7.26391f
C1806 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 0.03176f
C1807 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.06435f
C1808 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.10029f
C1809 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.82681f
C1810 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.07333f
C1811 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A VDD 1.0555f
C1812 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 0.20097f
C1813 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.01028f
C1814 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.06643f
C1815 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.08427f
C1816 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 2.0142f
C1817 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.22976f
C1818 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.09785f
C1819 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.09942f
C1820 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.11032f
C1821 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_final_switch_0.VOUT[0] 0.08765f
C1822 top_DAC_0/top_final_switch_0.VOUT[1] a_8173_15057# 0.01175f
C1823 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.3192f
C1824 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.73909f
C1825 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_final_switch_0.VOUT[4] 0.02498f
C1826 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_2300_13708# 0.03745f
C1827 a_5897_14150# VDDH 0.49013f
C1828 top_DAC_0/top_final_switch_0.VOUT[0] a_5897_15057# 0.03805f
C1829 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.01144f
C1830 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A VDDH 0.82663f
C1831 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 0.57986f
C1832 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.04811f
C1833 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.22293f
C1834 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.04333f
C1835 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.02124f
C1836 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.05591f
C1837 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 0.1278f
C1838 top_DAC_0/top_final_switch_0.VOUT[3] a_11081_13005# 0.03209f
C1839 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 VDDH 0.14505f
C1840 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.23003f
C1841 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 VDDH 0.11246f
C1842 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.02388f
C1843 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VOUT 0.44339f
C1844 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.2354f
C1845 top_DAC_0/top_rseg_n_dcell_0.SH[2] VDDH 0.63542f
C1846 VDDH DIN9 0.40422f
C1847 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_rseg_n_dcell_0.VS4 0.01859f
C1848 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD 0.21631f
C1849 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.0119f
C1850 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.12879f
C1851 top_DAC_0/top_final_switch_0.VOUT[0] a_5897_12507# 0.01061f
C1852 a_5897_15057# VOUT 0.04644f
C1853 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 0.0847f
C1854 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 2.29207f
C1855 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 ROUT1 0.01978f
C1856 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.11409f
C1857 top_DAC_0/top_final_switch_0.VOUT[4] VDDH 2.1005f
C1858 a_4978_9535# a_4978_8388# 0.015f
C1859 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.VS4 0.06276f
C1860 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.21449f
C1861 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.VH2 0.14076f
C1862 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.61812f
C1863 a_39768_20665# a_39768_20389# 0.02286f
C1864 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.28496f
C1865 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.02737f
C1866 a_5897_12507# VOUT 0.04473f
C1867 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 0.05245f
C1868 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 1.8445f
C1869 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.04809f
C1870 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.64115f
C1871 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.05622f
C1872 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.08198f
C1873 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.02015f
C1874 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.04929f
C1875 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 0.09809f
C1876 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 1.29067f
C1877 a_11081_14150# VOUT 0.06741f
C1878 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.05174f
C1879 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09272f
C1880 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.92259f
C1881 VDD DIN2 0.66783f
C1882 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.68733f
C1883 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] VDDH 0.89706f
C1884 a_45343_4828# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.01335f
C1885 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.24317f
C1886 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 4.14638f
C1887 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 VDDH 2.7521f
C1888 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.10646f
C1889 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_final_switch_0.VOUT[1] 0.20372f
C1890 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.29339f
C1891 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.09612f
C1892 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] VDDH 0.01064f
C1893 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.01148f
C1894 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.19471f
C1895 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.01383f
C1896 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.07239f
C1897 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 VDDH 0.16077f
C1898 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.10246f
C1899 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.01125f
C1900 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.12989f
C1901 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.10185f
C1902 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_6445_12507# 0.02171f
C1903 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.16754f
C1904 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.05224f
C1905 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 1.85532f
C1906 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.3835f
C1907 a_39861_22496# ROUT2 0.13835f
C1908 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.03539f
C1909 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.05972f
C1910 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.09312f
C1911 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 0.18788f
C1912 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.VS1 0.07172f
C1913 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04931f
C1914 a_2300_15118# VDDH 0.54014f
C1915 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.02165f
C1916 a_11081_12507# VOUT 0.04471f
C1917 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 0.54711f
C1918 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 0.04809f
C1919 DIN0 DIN1 0.32901f
C1920 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.06525f
C1921 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B VDD 0.4727f
C1922 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] DIN6 0.01584f
C1923 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.SH[4] 16.3155f
C1924 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1636_15118# 0.03043f
C1925 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 0.09709f
C1926 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 4.14551f
C1927 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.0386f
C1928 top_DAC_0/top_final_switch_0.VOUT[3] a_11081_14150# 0.01871f
C1929 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.06657f
C1930 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.08257f
C1931 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_final_switch_0.VOUT[0] 0.01642f
C1932 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C1933 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 VDDH 0.11563f
C1934 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_11629_15057# 0.04959f
C1935 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_final_switch_0.VOUT[0] 0.0398f
C1936 a_11629_14150# VDDH 0.49013f
C1937 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.02339f
C1938 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 0.16825f
C1939 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.01514f
C1940 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx a_1896_10974# 0.02584f
C1941 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.04839f
C1942 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.53572f
C1943 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.05787f
C1944 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.VH2 0.05427f
C1945 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_final_switch_0.VOUT[1] 0.01422f
C1946 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.10148f
C1947 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.09623f
C1948 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] ROUT2 0.06337f
C1949 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.38211f
C1950 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.10002f
C1951 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD VOUT 0.6262f
C1952 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A VDD 0.59039f
C1953 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.15687f
C1954 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_2678_20320# 0.01554f
C1955 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_11629_12507# 0.02171f
C1956 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.10472f
C1957 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.0981f
C1958 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 1.25806f
C1959 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 0.02201f
C1960 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 0.04735f
C1961 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.17104f
C1962 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.02147f
C1963 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C1964 VDD DIN3 0.67007f
C1965 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.0249f
C1966 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_11081_14150# 0.04959f
C1967 top_DAC_0/top_rseg_n_dcell_0.SH[4] VDDH 1.34727f
C1968 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 1.95068f
C1969 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 1.27523f
C1970 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 6.01491f
C1971 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_2300_13352# 0.03772f
C1972 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] VDDH 2.0654f
C1973 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B VDDH 2.1824f
C1974 top_DAC_0/top_final_switch_0.VOUT[1] VDDH 1.66034f
C1975 top_DAC_0/top_final_switch_0.VOUT[0] a_5897_14150# 0.01852f
C1976 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.04287f
C1977 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04845f
C1978 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.24146f
C1979 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 0.31985f
C1980 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN a_5642_9535# 0.01975f
C1981 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 17.3149f
C1982 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.08235f
C1983 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 0.03135f
C1984 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.04827f
C1985 top_DAC_0/top_final_switch_0.VOUT[3] a_11081_12507# 0.01061f
C1986 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 0.14746f
C1987 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 1.90588f
C1988 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.09304f
C1989 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.01808f
C1990 a_5897_14150# VOUT 0.06743f
C1991 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.VS1 0.0717f
C1992 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.10742f
C1993 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.VS4 0.01905f
C1994 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.01642f
C1995 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.07698f
C1996 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 7.06738f
C1997 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_final_switch_0.VOUT[4] 0.44592f
C1998 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 VDDH 0.04651f
C1999 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 VDDH 0.33162f
C2000 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.VL2 0.1484f
C2001 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05095f
C2002 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 VDDH 0.1547f
C2003 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.01034f
C2004 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.4555f
C2005 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.06121f
C2006 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.0672f
C2007 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.02775f
C2008 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.03397f
C2009 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 VOUT 0.02946f
C2010 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.VH3 0.13103f
C2011 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 1.26639f
C2012 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 0.10213f
C2013 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.04851f
C2014 a_5897_13005# a_6445_13005# 0.0103f
C2015 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 3.43068f
C2016 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 0.06052f
C2017 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.03545f
C2018 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 0.51079f
C2019 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 0.0481f
C2020 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] VDDH 0.88394f
C2021 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05296f
C2022 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx a_1896_10356# 0.05988f
C2023 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] DIN7 0.17937f
C2024 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_4978_10963# 0.01297f
C2025 top_DAC_0/top_final_switch_0.VOUT[4] VOUT 8.15099f
C2026 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.05823f
C2027 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.10018f
C2028 a_11081_15057# a_11629_15057# 0.0237f
C2029 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_final_switch_0.VOUT[3] 0.01686f
C2030 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.16603f
C2031 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_12809_15057# 0.04134f
C2032 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 16.8926f
C2033 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.06658f
C2034 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.09162f
C2035 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.01148f
C2036 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.17953f
C2037 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.09189f
C2038 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 1.15664f
C2039 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.01119f
C2040 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.0483f
C2041 a_2678_20320# VDDH 0.73328f
C2042 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09743f
C2043 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.96691f
C2044 VDD DIN4 0.67214f
C2045 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 0.02214f
C2046 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.14454f
C2047 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.04748f
C2048 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 0.02179f
C2049 DIN9 GND 2.58682f
C2050 DIN8 GND 2.24158f
C2051 DIN7 GND 2.21448f
C2052 DIN6 GND 2.18502f
C2053 DIN5 GND 2.16664f
C2054 DIN4 GND 2.15816f
C2055 DIN3 GND 2.13965f
C2056 DIN2 GND 2.11716f
C2057 DIN1 GND 2.1019f
C2058 DIN0 GND 2.34399f
C2059 VOUT GND 42.23114f
C2060 ROUT2 GND 14.28184f
C2061 ROUT1 GND 16.95354f
C2062 VDD GND 0.15684p
C2063 VDDH GND 0.7762p
C2064 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B GND 0.39231f
C2065 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y GND 0.3768f
C2066 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A GND 0.68099f
C2067 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y GND 0.70838f
C2068 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C GND 0.3332f
C2069 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B GND 0.32574f
C2070 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B GND 0.31137f
C2071 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A GND 0.25769f
C2072 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A GND 0.32968f
C2073 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y GND 0.45293f
C2074 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C GND 0.41678f
C2075 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B GND 0.42992f
C2076 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y GND 0.33977f
C2077 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A GND 0.73456f
C2078 a_45343_4828# GND 0.02142f $ **FLOATING
C2079 a_44471_4828# GND 0.02172f $ **FLOATING
C2080 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B GND 0.44413f
C2081 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A GND 0.49956f
C2082 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 GND 1.58565f
C2083 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 GND 1.01698f
C2084 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 GND 0.83396f
C2085 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 GND 0.84338f
C2086 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 GND 0.72928f
C2087 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 GND 0.81839f
C2088 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 GND 1.60815f
C2089 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 GND 1.05072f
C2090 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 GND 0.85279f
C2091 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 GND 0.85992f
C2092 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 GND 0.74171f
C2093 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 GND 0.83636f
C2094 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 GND 1.64361f
C2095 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 GND 1.10159f
C2096 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 GND 0.88377f
C2097 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 GND 0.74063f
C2098 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 GND 0.77336f
C2099 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 GND 0.88264f
C2100 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 GND 2.61761f
C2101 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 GND 1.84052f
C2102 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 GND 1.36319f
C2103 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 GND 1.54449f
C2104 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 GND 1.34744f
C2105 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 GND 2.56072f
C2106 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 GND 1.89955f
C2107 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 GND 0.92879f
C2108 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 GND 1.14314f
C2109 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 GND 0.8323f
C2110 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 GND 0.71956f
C2111 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 GND 0.79316f
C2112 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 GND 1.88785f
C2113 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 GND 0.87481f
C2114 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 GND 1.12833f
C2115 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 GND 0.79452f
C2116 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 GND 0.69232f
C2117 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 GND 0.75887f
C2118 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 GND 1.8686f
C2119 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 GND 0.85431f
C2120 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 GND 1.11076f
C2121 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 GND 0.77008f
C2122 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 GND 0.66926f
C2123 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 GND 0.73878f
C2124 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 GND 2.28785f
C2125 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 GND 0.84039f
C2126 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 GND 1.16435f
C2127 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 GND 0.77204f
C2128 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 GND 0.71421f
C2129 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 GND 0.72923f
C2130 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A GND 0.9729f
C2131 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 GND 1.00383f
C2132 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 GND 0.94283f
C2133 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 GND 0.92717f
C2134 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 GND 0.86196f
C2135 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 GND 1.47451f
C2136 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 GND 2.4135f
C2137 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 GND 3.29904f
C2138 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 GND 0.999f
C2139 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 GND 0.9622f
C2140 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 GND 0.95203f
C2141 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 GND 0.93445f
C2142 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 GND 1.12363f
C2143 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 GND 2.48462f
C2144 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 GND 3.37108f
C2145 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 GND 1.03387f
C2146 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 GND 0.98141f
C2147 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 GND 0.97038f
C2148 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 GND 0.95434f
C2149 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 GND 1.13854f
C2150 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 GND 2.48866f
C2151 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 GND 3.44747f
C2152 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 GND 1.10941f
C2153 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 GND 1.06449f
C2154 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 GND 1.50227f
C2155 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 GND 1.05333f
C2156 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 GND 1.44211f
C2157 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 GND 2.61871f
C2158 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 GND 4.12386f
C2159 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 GND 0.98593f
C2160 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 GND 1.48196f
C2161 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 GND 0.92766f
C2162 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 GND 2.04138f
C2163 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 GND 2.40878f
C2164 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 GND 3.28652f
C2165 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 GND 0.83546f
C2166 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 GND 0.83142f
C2167 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 GND 1.31433f
C2168 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 GND 0.8334f
C2169 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 GND 1.49005f
C2170 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 GND 2.32599f
C2171 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 GND 3.09657f
C2172 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 GND 0.79398f
C2173 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 GND 0.79447f
C2174 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 GND 1.27612f
C2175 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 GND 0.80491f
C2176 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 GND 1.44901f
C2177 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 GND 2.29709f
C2178 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 GND 3.04183f
C2179 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 GND 0.76536f
C2180 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 GND 0.79117f
C2181 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 GND 1.26691f
C2182 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 GND 0.79436f
C2183 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 GND 1.44302f
C2184 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 GND 2.29524f
C2185 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 GND 3.03441f
C2186 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A GND 0.77271f
C2187 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] GND 4.20597f
C2188 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] GND 8.05747f
C2189 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] GND 4.29275f
C2190 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] GND 3.2508f
C2191 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A GND 0.76913f
C2192 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A GND 0.77224f
C2193 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 GND 1.4175f
C2194 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 GND 1.32581f
C2195 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 GND 1.37474f
C2196 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GND 2.6963f
C2197 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GND 3.30161f
C2198 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND 5.16186f
C2199 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND 42.83636f
C2200 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND 8.84505f
C2201 a_5642_8388# GND 0.11496f $ **FLOATING
C2202 a_4978_8388# GND 0.10989f $ **FLOATING
C2203 a_5642_9535# GND 0.11145f $ **FLOATING
C2204 a_4978_9535# GND 0.10301f $ **FLOATING
C2205 a_5642_10963# GND 0.35967f $ **FLOATING
C2206 a_4978_10963# GND 0.36693f $ **FLOATING
C2207 a_5642_11461# GND 0.38872f $ **FLOATING
C2208 a_4978_11461# GND 0.34413f $ **FLOATING
C2209 a_2678_10356# GND 0.3141f $ **FLOATING
C2210 a_1896_10356# GND 0.31627f $ **FLOATING
C2211 a_2678_10974# GND 0.31147f $ **FLOATING
C2212 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 GND 32.24118f
C2213 a_1896_10974# GND 0.31363f $ **FLOATING
C2214 top_DAC_0/top_rseg_n_dcell_0.VS4 GND 1.44778f
C2215 top_DAC_0/top_rseg_n_dcell_0.SH[4] GND 31.09953f
C2216 top_DAC_0/top_rseg_n_dcell_0.SH[3] GND 32.83591f
C2217 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 GND 9.87811f
C2218 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 GND 9.79582f
C2219 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 GND 10.80865f
C2220 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 GND 9.54184f
C2221 top_DAC_0/top_rseg_n_dcell_0.VS1 GND 7.91312f
C2222 top_DAC_0/top_rseg_n_dcell_0.SH[2] GND 36.92257f
C2223 top_DAC_0/top_rseg_n_dcell_0.SH[1] GND 26.97365f
C2224 a_12809_12507# GND 0.23775f $ **FLOATING
C2225 a_11629_12507# GND 0.2248f $ **FLOATING
C2226 a_12809_13005# GND 0.23111f $ **FLOATING
C2227 a_11629_13005# GND 0.2208f $ **FLOATING
C2228 a_11081_12507# GND 0.22626f $ **FLOATING
C2229 a_9901_12507# GND 0.22553f $ **FLOATING
C2230 a_11081_13005# GND 0.2208f $ **FLOATING
C2231 a_9901_13005# GND 0.2208f $ **FLOATING
C2232 a_9353_12507# GND 0.22485f $ **FLOATING
C2233 a_8173_12507# GND 0.22611f $ **FLOATING
C2234 a_9353_13005# GND 0.2208f $ **FLOATING
C2235 a_8173_13005# GND 0.2208f $ **FLOATING
C2236 a_7625_12507# GND 0.22504f $ **FLOATING
C2237 a_6445_12507# GND 0.22721f $ **FLOATING
C2238 a_7625_13005# GND 0.2208f $ **FLOATING
C2239 a_6445_13005# GND 0.2208f $ **FLOATING
C2240 a_5897_12507# GND 0.22396f $ **FLOATING
C2241 a_4717_12507# GND 0.23225f $ **FLOATING
C2242 a_5897_13005# GND 0.22049f $ **FLOATING
C2243 a_4717_13005# GND 0.23057f $ **FLOATING
C2244 a_2678_11886# GND 0.31079f $ **FLOATING
C2245 a_1896_11886# GND 0.31296f $ **FLOATING
C2246 a_2678_12504# GND 0.31285f $ **FLOATING
C2247 a_1896_12504# GND 0.31297f $ **FLOATING
C2248 a_12809_14150# GND 0.03735f $ **FLOATING
C2249 a_12809_15057# GND 0.03468f $ **FLOATING
C2250 top_DAC_0/top_final_switch_0.VOUT[4] GND 7.39747f
C2251 top_DAC_0/top_final_switch_0.VOUT[3] GND 6.06922f
C2252 top_DAC_0/top_final_switch_0.VOUT[2] GND 5.72707f
C2253 top_DAC_0/top_final_switch_0.VOUT[1] GND 5.82584f
C2254 a_4717_14150# GND 0.03708f $ **FLOATING
C2255 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB GND 4.94893f
C2256 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA GND 11.89824f
C2257 top_DAC_0/top_final_switch_0.VOUT[0] GND 6.28621f
C2258 a_4717_15057# GND 0.03501f $ **FLOATING
C2259 a_2300_13352# GND 0.27287f $ **FLOATING
C2260 a_1636_13352# GND 0.27787f $ **FLOATING
C2261 a_2300_13708# GND 0.26729f $ **FLOATING
C2262 a_1636_13708# GND 0.26729f $ **FLOATING
C2263 a_2300_14353# GND 0.06968f $ **FLOATING
C2264 a_1636_14353# GND 0.06968f $ **FLOATING
C2265 a_2300_15118# GND 0.06696f $ **FLOATING
C2266 a_1636_15118# GND 0.06696f $ **FLOATING
C2267 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.79418f
C2268 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.67704f
C2269 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.643f
C2270 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.61395f
C2271 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.65617f
C2272 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] GND 10.40641f
C2273 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.67288f
C2274 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.64256f
C2275 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] GND 9.02532f
C2276 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.61568f
C2277 top_DAC_0/top_rseg_n_dcell_0.VL2 GND 4.45416f
C2278 top_DAC_0/top_rseg_n_dcell_0.VH2 GND 4.55966f
C2279 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] GND 18.48214f
C2280 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 GND 6.70388f
C2281 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] GND 15.81766f
C2282 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 GND 17.84785f
C2283 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] GND 15.60426f
C2284 top_DAC_0/top_rseg_n_dcell_0.VH3 GND 3.11056f
C2285 top_DAC_0/top_rseg_n_dcell_0.VL3 GND 3.18256f
C2286 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 GND 14.78577f
C2287 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 GND 13.01433f
C2288 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] GND 17.41479f
C2289 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] GND 17.13611f
C2290 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] GND 18.52176f
C2291 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] GND 20.01692f
C2292 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 GND 18.02337f
C2293 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] GND 16.36461f
C2294 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] GND 15.5843f
C2295 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.61845f
C2296 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] GND 7.27954f
C2297 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.66383f
C2298 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] GND 7.07277f
C2299 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.63305f
C2300 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] GND 7.21126f
C2301 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] GND 8.73283f
C2302 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.75299f
C2303 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] GND 15.57737f
C2304 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] GND 15.5338f
C2305 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] GND 15.68769f
C2306 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] GND 50.2481f
C2307 a_39883_19098# GND 0.21843f $ **FLOATING
C2308 a_37277_19098# GND 0.24267f $ **FLOATING
C2309 a_39883_19479# GND 0.20382f $ **FLOATING
C2310 a_37737_19479# GND 0.18912f $ **FLOATING
C2311 a_39883_19854# GND 0.20634f $ **FLOATING
C2312 a_38617_19854# GND 0.21532f $ **FLOATING
C2313 a_37595_19462# GND 0.15668f $ **FLOATING
C2314 a_36813_19462# GND 0.19962f $ **FLOATING
C2315 a_37595_19760# GND 0.19172f $ **FLOATING
C2316 a_36813_19760# GND 0.19708f $ **FLOATING
C2317 a_39768_20389# GND 0.17117f $ **FLOATING
C2318 a_38584_20389# GND 0.17006f $ **FLOATING
C2319 a_39768_20665# GND 0.17317f $ **FLOATING
C2320 a_38584_20665# GND 0.17331f $ **FLOATING
C2321 a_37804_20295# GND 0.18145f $ **FLOATING
C2322 a_37022_20295# GND 0.17721f $ **FLOATING
C2323 a_37804_20713# GND 0.18276f $ **FLOATING
C2324 a_37022_20713# GND 0.17864f $ **FLOATING
C2325 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD GND 0.89224f
C2326 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD GND 0.97215f
C2327 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD GND 0.75334f
C2328 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD GND 1.35643f
C2329 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 GND 5.23006f
C2330 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD GND 1.83958f
C2331 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN GND 44.39035f
C2332 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] GND 17.68056f
C2333 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] GND 17.46266f
C2334 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] GND 18.87729f
C2335 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] GND 17.2396f
C2336 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] GND 17.84095f
C2337 a_40525_21457# GND 0.05335f $ **FLOATING
C2338 a_39861_21457# GND 0.01074f $ **FLOATING
C2339 a_41907_22057# GND 0.01121f $ **FLOATING
C2340 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV GND 11.21902f
C2341 a_44067_22496# GND 0.18164f $ **FLOATING
C2342 a_39861_22496# GND 0.0387f $ **FLOATING
C2343 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV GND 19.55606f
C2344 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC GND 4.69893f
C2345 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC GND 11.75439f
C2346 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 GND 0.2652f
C2347 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 GND 0.28781f
C2348 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 GND 2.93597f
C2349 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 GND 3.21084f
C2350 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 GND 2.10079f
C2351 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 GND 9.78667f
C2352 a_2678_16243# GND 0.03553f $ **FLOATING
C2353 a_1896_16243# GND 0.04167f $ **FLOATING
C2354 a_2678_17510# GND 0.03283f $ **FLOATING
C2355 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B GND 6.69444f
C2356 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx GND 10.82046f
C2357 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 GND 6.04689f
C2358 a_1896_17510# GND 0.04167f $ **FLOATING
C2359 a_2678_19053# GND 0.03256f $ **FLOATING
C2360 a_1896_19053# GND 0.04167f $ **FLOATING
C2361 a_2678_20320# GND 0.03256f $ **FLOATING
C2362 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A GND 2.76149f
C2363 a_1896_20320# GND 0.04167f $ **FLOATING
C2364 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 GND 16.97545f
C2365 a_2678_21703# GND 0.03256f $ **FLOATING
C2366 a_1896_21703# GND 0.04167f $ **FLOATING
C2367 a_2678_22970# GND 0.03813f $ **FLOATING
C2368 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND 4.61337f
C2369 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND 9.31942f
C2370 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax GND 2.76712f
C2371 a_1896_22970# GND 0.04724f $ **FLOATING
C2372 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.t2 GND 0.0447f
C2373 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.t1 GND 0.19887f
C2374 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.n0 GND 4.85619f
C2375 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5.t0 GND 0.20023f
C2376 ROUT2.t1 GND 0.02488f
C2377 ROUT2.t2 GND 1.41742f
C2378 ROUT2.t4 GND 2.04267f
C2379 ROUT2.t5 GND 2.33027f
C2380 ROUT2.t0 GND 1.70501f
C2381 ROUT2.n0 GND 1.47089f
C2382 ROUT2.n1 GND 0.21478f
C2383 ROUT2.t3 GND 0.02473f
C2384 ROUT2.n2 GND 0.02835f
C2385 ROUT2.n3 GND 0.09357f
C2386 a_19276_8950.t2 GND 0.07488f
C2387 a_19276_8950.t1 GND 0.07606f
C2388 a_19276_8950.n0 GND 5.28272f
C2389 a_19276_8950.t0 GND 0.06634f
C2390 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t1 GND 0.39374f
C2391 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t3 GND 0.19462f
C2392 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t2 GND 0.21619f
C2393 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n0 GND 1.60492f
C2394 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t0 GND 0.20263f
C2395 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n1 GND 3.37677f
C2396 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.t2 GND 0.20596f
C2397 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.t1 GND 0.22743f
C2398 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.n0 GND 4.83206f
C2399 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41.t0 GND 0.03454f
C2400 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t2 GND 0.01292f
C2401 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t1 GND 0.09788f
C2402 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t0 GND 0.10105f
C2403 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.n0 GND 1.62825f
C2404 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.t2 GND 0.04657f
C2405 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.t0 GND 0.13984f
C2406 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.t1 GND 0.13973f
C2407 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41.n0 GND 2.57846f
C2408 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t2 GND 0.02279f
C2409 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t1 GND 0.1333f
C2410 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t0 GND 0.39583f
C2411 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.n0 GND 2.7632f
C2412 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.t2 GND 0.19941f
C2413 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.t1 GND 0.02987f
C2414 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.n0 GND 4.06638f
C2415 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38.t0 GND 0.20435f
C2416 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t1 GND 0.13031f
C2417 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y GND 0.31167f
C2418 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t2 GND 0.30126f
C2419 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[4] GND 5.44042f
C2420 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[4] GND 0.68417f
C2421 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 GND 0.21176f
C2422 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t0 GND 0.09569f
C2423 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 GND 0.02473f
C2424 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t2 GND 0.02752f
C2425 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t1 GND 0.15141f
C2426 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t0 GND 0.17047f
C2427 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.n0 GND 2.83038f
C2428 a_21099_20174.t2 GND 0.19205f
C2429 a_21099_20174.t3 GND 0.07964f
C2430 a_21099_20174.n0 GND 5.71483f
C2431 a_21099_20174.t1 GND 0.0575f
C2432 a_21099_20174.n1 GND 4.4887f
C2433 a_21099_20174.t0 GND 0.1673f
C2434 a_22479_20174.t2 GND 0.1868f
C2435 a_22479_20174.t3 GND 0.07658f
C2436 a_22479_20174.n0 GND 5.49565f
C2437 a_22479_20174.t1 GND 0.07075f
C2438 a_22479_20174.n1 GND 4.99847f
C2439 a_22479_20174.t0 GND 0.17175f
C2440 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t1 GND 0.02245f
C2441 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t0 GND 0.13087f
C2442 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t2 GND 0.40073f
C2443 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.n0 GND 2.77278f
C2444 a_14607_6250.t3 GND 0.08343f
C2445 a_14607_6250.t2 GND 0.08172f
C2446 a_14607_6250.t4 GND 0.06448f
C2447 a_14607_6250.n0 GND 3.71167f
C2448 a_14607_6250.t1 GND 0.0952f
C2449 a_14607_6250.n1 GND 4.09447f
C2450 a_14607_6250.n2 GND 4.80455f
C2451 a_14607_6250.t0 GND 0.06448f
C2452 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t2 GND 0.01506f
C2453 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t1 GND 0.09156f
C2454 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t0 GND 0.08868f
C2455 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.n0 GND 1.45797f
C2456 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.t1 GND 0.09894f
C2457 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.t2 GND 0.01383f
C2458 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.n0 GND 1.89904f
C2459 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26.t0 GND 0.08819f
C2460 a_24209_18133.t3 GND 0.03955f
C2461 a_24209_18133.t2 GND 0.03423f
C2462 a_24209_18133.n0 GND 1.24539f
C2463 a_24209_18133.t1 GND 0.03423f
C2464 a_24209_18133.n1 GND 0.78371f
C2465 a_24209_18133.t4 GND 0.03423f
C2466 a_24209_18133.n2 GND 1.28824f
C2467 a_24209_18133.t0 GND 0.04042f
C2468 a_19000_8950.t2 GND 0.07342f
C2469 a_19000_8950.t1 GND 0.07455f
C2470 a_19000_8950.n0 GND 5.18539f
C2471 a_19000_8950.t0 GND 0.06664f
C2472 a_13779_6250.t3 GND 0.04948f
C2473 a_13779_6250.t2 GND 0.04849f
C2474 a_13779_6250.t4 GND 0.039f
C2475 a_13779_6250.n0 GND 2.19006f
C2476 a_13779_6250.t1 GND 0.05645f
C2477 a_13779_6250.n1 GND 2.38608f
C2478 a_13779_6250.n2 GND 2.59144f
C2479 a_13779_6250.t0 GND 0.039f
C2480 a_33910_8950.t1 GND 0.09187f
C2481 a_33910_8950.t2 GND 0.10902f
C2482 a_33910_8950.n0 GND 5.42682f
C2483 a_33910_8950.t0 GND 0.0723f
C2484 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t2 GND 0.01248f
C2485 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t1 GND 0.09062f
C2486 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t0 GND 0.08856f
C2487 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.n0 GND 1.58095f
C2488 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t1 GND 0.01438f
C2489 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t2 GND 0.0778f
C2490 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t0 GND 0.08737f
C2491 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.n0 GND 1.43709f
C2492 a_15905_7686.t3 GND 0.07983f
C2493 a_15905_7686.t1 GND 0.08121f
C2494 a_15905_7686.n0 GND 3.82467f
C2495 a_15905_7686.t2 GND 0.09398f
C2496 a_15905_7686.t4 GND 0.07505f
C2497 a_15905_7686.n1 GND 5.374f
C2498 a_15905_7686.n2 GND 2.89621f
C2499 a_15905_7686.t0 GND 0.07505f
C2500 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t1 GND 0.01506f
C2501 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t2 GND 0.08796f
C2502 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t0 GND 0.0907f
C2503 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.n0 GND 1.45497f
C2504 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.t2 GND 0.10272f
C2505 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.t1 GND 0.01601f
C2506 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.n0 GND 2.08049f
C2507 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39.t0 GND 0.10078f
C2508 a_34580_8950.t1 GND 0.10677f
C2509 a_34580_8950.t2 GND 0.12828f
C2510 a_34580_8950.n0 GND 6.09613f
C2511 a_34580_8950.t0 GND 0.06882f
C2512 a_31318_7686.t1 GND 0.10563f
C2513 a_31318_7686.t3 GND 0.08474f
C2514 a_31318_7686.n0 GND 3.77304f
C2515 a_31318_7686.t4 GND 0.08064f
C2516 a_31318_7686.n1 GND 2.70857f
C2517 a_31318_7686.t2 GND 0.14779f
C2518 a_31318_7686.n2 GND 5.91896f
C2519 a_31318_7686.t0 GND 0.08064f
C2520 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t2 GND 0.01583f
C2521 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t1 GND 0.08108f
C2522 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t0 GND 0.09013f
C2523 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.n0 GND 1.56677f
C2524 a_16181_7686.t3 GND 0.08006f
C2525 a_16181_7686.t1 GND 0.07704f
C2526 a_16181_7686.n0 GND 3.67426f
C2527 a_16181_7686.t2 GND 0.09319f
C2528 a_16181_7686.t4 GND 0.07394f
C2529 a_16181_7686.n1 GND 5.40641f
C2530 a_16181_7686.n2 GND 2.82116f
C2531 a_16181_7686.t0 GND 0.07394f
C2532 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.t1 GND 0.16127f
C2533 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.t2 GND 0.63594f
C2534 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.n0 GND 4.57733f
C2535 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40.t0 GND 0.02546f
C2536 a_22755_20174.t3 GND 0.16937f
C2537 a_22755_20174.t4 GND 0.06934f
C2538 a_22755_20174.n0 GND 4.88352f
C2539 a_22755_20174.t2 GND 0.06731f
C2540 a_22755_20174.n1 GND 0.88718f
C2541 a_22755_20174.t1 GND 0.06731f
C2542 a_22755_20174.n2 GND 4.60037f
C2543 a_22755_20174.t0 GND 0.15559f
C2544 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t0 GND 0.05654f
C2545 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t1 GND 0.05718f
C2546 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n0 GND 1.04424f
C2547 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t3 GND 0.05624f
C2548 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t2 GND 0.0538f
C2549 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n1 GND 0.81076f
C2550 a_15317_6250.t3 GND 0.09555f
C2551 a_15317_6250.t2 GND 0.09358f
C2552 a_15317_6250.t4 GND 0.07299f
C2553 a_15317_6250.n0 GND 5.4004f
C2554 a_15317_6250.t1 GND 0.0965f
C2555 a_15317_6250.n1 GND 4.00369f
C2556 a_15317_6250.n2 GND 4.6643f
C2557 a_15317_6250.t0 GND 0.07299f
C2558 a_15041_6250.t3 GND 0.08408f
C2559 a_15041_6250.t2 GND 0.08235f
C2560 a_15041_6250.t4 GND 0.0646f
C2561 a_15041_6250.n0 GND 4.76416f
C2562 a_15041_6250.t1 GND 0.08975f
C2563 a_15041_6250.n1 GND 3.79219f
C2564 a_15041_6250.n2 GND 3.95828f
C2565 a_15041_6250.t0 GND 0.0646f
C2566 a_19670_8950.t2 GND 0.0805f
C2567 a_19670_8950.t1 GND 0.08183f
C2568 a_19670_8950.n0 GND 5.8709f
C2569 a_19670_8950.t0 GND 0.06677f
C2570 a_27896_6250.t1 GND 0.13945f
C2571 a_27896_6250.t4 GND 0.0817f
C2572 a_27896_6250.n0 GND 5.49877f
C2573 a_27896_6250.t3 GND 0.17983f
C2574 a_27896_6250.n1 GND 4.84462f
C2575 a_27896_6250.t2 GND 0.17181f
C2576 a_27896_6250.n2 GND 5.30212f
C2577 a_27896_6250.t0 GND 0.0817f
C2578 a_15593_6250.t3 GND 0.09595f
C2579 a_15593_6250.t2 GND 0.09395f
C2580 a_15593_6250.t4 GND 0.07288f
C2581 a_15593_6250.n0 GND 5.40773f
C2582 a_15593_6250.t1 GND 0.09172f
C2583 a_15593_6250.n1 GND 3.72117f
C2584 a_15593_6250.n2 GND 4.84372f
C2585 a_15593_6250.t0 GND 0.07288f
C2586 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t0 GND 0.08474f
C2587 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n0 GND 0.03475f
C2588 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n1 GND 0.0748f
C2589 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n2 GND 0.04966f
C2590 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t1 GND 0.08119f
C2591 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n3 GND 0.01025f
C2592 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t4 GND 0.16835f
C2593 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t8 GND 0.16754f
C2594 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n4 GND 0.52525f
C2595 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t11 GND 0.16754f
C2596 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n5 GND 0.26303f
C2597 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t3 GND 0.16754f
C2598 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n6 GND 0.26303f
C2599 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t7 GND 0.16754f
C2600 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n7 GND 0.26303f
C2601 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t16 GND 0.16754f
C2602 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n8 GND 0.26303f
C2603 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t12 GND 0.16754f
C2604 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n9 GND 0.26303f
C2605 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t6 GND 0.16568f
C2606 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t9 GND 0.16835f
C2607 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t17 GND 0.16835f
C2608 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t14 GND 0.16754f
C2609 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n10 GND 0.52525f
C2610 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t13 GND 0.16754f
C2611 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n11 GND 0.26303f
C2612 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t10 GND 0.16754f
C2613 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n12 GND 0.26303f
C2614 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t15 GND 0.16754f
C2615 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n13 GND 0.26303f
C2616 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t5 GND 0.16754f
C2617 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n14 GND 0.26303f
C2618 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n15 GND 0.43732f
C2619 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.t2 GND 0.16568f
C2620 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n16 GND 0.42527f
C2621 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n17 GND 0.19515f
C2622 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n18 GND 15.7048f
C2623 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2.n19 GND 0.08218f
C2624 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t0 GND 0.01441f
C2625 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t1 GND 0.07654f
C2626 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t2 GND 0.08569f
C2627 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.n0 GND 1.43498f
C2628 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t1 GND 0.02728f
C2629 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t2 GND 0.16768f
C2630 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t0 GND 0.1501f
C2631 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.n0 GND 2.84284f
C2632 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t3 GND 0.03817f
C2633 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t2 GND 0.03817f
C2634 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 GND 0.08382f
C2635 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y GND 0.1918f
C2636 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 GND 0.03616f
C2637 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.A GND 0.01088f
C2638 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t7 GND 0.06318f
C2639 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t4 GND 0.03945f
C2640 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 GND 0.12027f
C2641 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 GND 0.07308f
C2642 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.A GND 0.01088f
C2643 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t8 GND 0.06318f
C2644 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t6 GND 0.03945f
C2645 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 GND 0.12027f
C2646 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 GND 0.03223f
C2647 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 GND 0.66246f
C2648 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[0] GND 2.72474f
C2649 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t5 GND 0.23963f
C2650 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 GND 11.603f
C2651 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 GND 1.68418f
C2652 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t1 GND 0.02481f
C2653 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t0 GND 0.02481f
C2654 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 GND 0.05916f
C2655 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 GND 0.11622f
C2656 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t3 GND 0.04311f
C2657 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t2 GND 0.04311f
C2658 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 GND 0.09469f
C2659 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y GND 0.21666f
C2660 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 GND 0.04085f
C2661 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t4 GND 0.76823f
C2662 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 GND 16.1392f
C2663 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t1 GND 0.02802f
C2664 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t0 GND 0.02802f
C2665 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 GND 0.06682f
C2666 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 GND 0.13128f
C2667 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.t2 GND 0.03678f
C2668 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.t0 GND 0.12308f
C2669 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.t1 GND 0.36729f
C2670 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40.n0 GND 2.56969f
C2671 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t1 GND 0.16796f
C2672 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t2 GND 0.63095f
C2673 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.n0 GND 4.13463f
C2674 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t3 GND 0.02217f
C2675 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.n1 GND 1.41681f
C2676 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8.t0 GND 0.02748f
C2677 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.t2 GND 0.10458f
C2678 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.t1 GND 0.01471f
C2679 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.n0 GND 2.07892f
C2680 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43.t0 GND 0.10179f
C2681 a_20222_8950.t2 GND 0.08054f
C2682 a_20222_8950.t1 GND 0.08241f
C2683 a_20222_8950.n0 GND 5.87337f
C2684 a_20222_8950.t0 GND 0.06369f
C2685 a_17167_7686.t3 GND 0.08487f
C2686 a_17167_7686.t1 GND 0.07389f
C2687 a_17167_7686.n0 GND 4.0948f
C2688 a_17167_7686.t2 GND 0.09304f
C2689 a_17167_7686.t4 GND 0.07249f
C2690 a_17167_7686.n1 GND 5.60801f
C2691 a_17167_7686.n2 GND 2.60041f
C2692 a_17167_7686.t0 GND 0.07249f
C2693 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t0 GND -0.50828f
C2694 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t1 GND -3.67942f
C2695 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t3 GND -2.37382f
C2696 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t2 GND -2.36382f
C2697 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n0 GND -3.97308f
C2698 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t4 GND -2.36382f
C2699 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n1 GND -3.49244f
C2700 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n2 GND -5.38322f
C2701 a_17443_7686.t3 GND 0.04297f
C2702 a_17443_7686.t1 GND 0.0365f
C2703 a_17443_7686.n0 GND 2.11432f
C2704 a_17443_7686.t2 GND 0.04624f
C2705 a_17443_7686.t4 GND 0.03583f
C2706 a_17443_7686.n1 GND 2.81877f
C2707 a_17443_7686.n2 GND 1.26954f
C2708 a_17443_7686.t0 GND 0.03583f
C2709 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t1 GND 0.01499f
C2710 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t2 GND 0.09144f
C2711 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t0 GND 0.08878f
C2712 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.n0 GND 1.46182f
C2713 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t2 GND 0.01209f
C2714 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t1 GND 0.08753f
C2715 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t0 GND 0.08547f
C2716 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.n0 GND 1.50136f
C2717 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.t0 GND 0.03636f
C2718 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.t2 GND 0.12209f
C2719 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.t1 GND 0.36895f
C2720 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24.n0 GND 2.57743f
C2721 a_29158_6250.t1 GND 0.14531f
C2722 a_29158_6250.t4 GND 0.08367f
C2723 a_29158_6250.n0 GND 4.77562f
C2724 a_29158_6250.t3 GND 0.14572f
C2725 a_29158_6250.n1 GND 4.0453f
C2726 a_29158_6250.t2 GND 0.17762f
C2727 a_29158_6250.n2 GND 6.44309f
C2728 a_29158_6250.t0 GND 0.08367f
C2729 a_15869_6250.t3 GND 0.04927f
C2730 a_15869_6250.t2 GND 0.04824f
C2731 a_15869_6250.t4 GND 0.03722f
C2732 a_15869_6250.n0 GND 2.76876f
C2733 a_15869_6250.t1 GND 0.04443f
C2734 a_15869_6250.n1 GND 1.74851f
C2735 a_15869_6250.n2 GND 2.56635f
C2736 a_15869_6250.t0 GND 0.03722f
C2737 a_20498_8950.t2 GND 0.04106f
C2738 a_20498_8950.t1 GND 0.04203f
C2739 a_20498_8950.n0 GND 2.9852f
C2740 a_20498_8950.t0 GND 0.03172f
C2741 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t2 GND 0.01294f
C2742 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t1 GND 0.10145f
C2743 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t0 GND 0.09797f
C2744 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.n0 GND 1.62712f
C2745 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.t2 GND 0.02493f
C2746 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.t1 GND 0.09805f
C2747 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.n0 GND 2.57844f
C2748 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7.t0 GND 0.09858f
C2749 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.t2 GND 0.02096f
C2750 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.t1 GND 0.52014f
C2751 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.n0 GND 4.09913f
C2752 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8.t0 GND 0.15978f
C2753 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.t1 GND 0.23806f
C2754 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.t2 GND 0.03472f
C2755 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.n0 GND 4.61553f
C2756 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25.t0 GND 0.21169f
C2757 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.t2 GND 0.0256f
C2758 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.t1 GND 0.59039f
C2759 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.n0 GND 4.42116f
C2760 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24.t0 GND 0.16286f
C2761 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.t2 GND 0.09067f
C2762 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.t1 GND 0.10022f
C2763 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.n0 GND 2.09413f
C2764 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42.t0 GND 0.01498f
C2765 a_20547_20174.t2 GND 0.12781f
C2766 a_20547_20174.t1 GND 0.05892f
C2767 a_20547_20174.n0 GND 4.03512f
C2768 a_20547_20174.t3 GND 0.06702f
C2769 a_20547_20174.n1 GND 5.04796f
C2770 a_20547_20174.t0 GND 0.16318f
C2771 a_22469_18133.t3 GND 0.06328f
C2772 a_22469_18133.t5 GND 0.0616f
C2773 a_22469_18133.n0 GND 1.91453f
C2774 a_22469_18133.t2 GND 0.06202f
C2775 a_22469_18133.n1 GND 1.68038f
C2776 a_22469_18133.t1 GND 0.06202f
C2777 a_22469_18133.n2 GND 1.49729f
C2778 a_22469_18133.t4 GND 0.06202f
C2779 a_22469_18133.n3 GND 2.52226f
C2780 a_22469_18133.t0 GND 0.07458f
C2781 a_4415_23194.t0 GND 0.23302f
C2782 a_4415_23194.t4 GND 8.33848f
C2783 a_4415_23194.t7 GND 6.5048f
C2784 a_4415_23194.n0 GND 3.76697f
C2785 a_4415_23194.t6 GND 8.33848f
C2786 a_4415_23194.t2 GND 6.5048f
C2787 a_4415_23194.n1 GND 3.96448f
C2788 a_4415_23194.t3 GND 0.0891f
C2789 a_4415_23194.t5 GND 0.30089f
C2790 a_4415_23194.n2 GND 2.48064f
C2791 a_4415_23194.n3 GND 0.57795f
C2792 a_4415_23194.n4 GND 0.53655f
C2793 a_4415_23194.n5 GND 2.67475f
C2794 a_4415_23194.t1 GND 0.0891f
C2795 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.t2 GND 0.20441f
C2796 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.t1 GND 0.03593f
C2797 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.n0 GND 5.13537f
C2798 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9.t0 GND 0.22429f
C2799 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.t2 GND 0.09859f
C2800 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.t1 GND 0.01938f
C2801 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.n0 GND 2.39212f
C2802 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10.t0 GND 0.08991f
C2803 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t5 GND 0.1888f
C2804 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[4] GND 3.43312f
C2805 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[4] GND 0.36483f
C2806 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.Y GND 0.04408f
C2807 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t1 GND 0.0216f
C2808 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 GND 0.06165f
C2809 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 GND 0.04788f
C2810 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t2 GND 0.01404f
C2811 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t0 GND 0.01404f
C2812 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 GND 0.06081f
C2813 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 GND 0.09879f
C2814 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 GND 0.30007f
C2815 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t4 GND 0.02235f
C2816 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t3 GND 0.03579f
C2817 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 GND 0.06697f
C2818 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n6 GND 0.01729f
C2819 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t1 GND 0.06405f
C2820 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t2 GND 0.14686f
C2821 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[3] GND 2.03364f
C2822 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[3] GND 0.20139f
C2823 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_0.Y GND 0.08421f
C2824 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 GND 0.12812f
C2825 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t0 GND 0.04173f
C2826 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.t2 GND 0.01499f
C2827 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.t1 GND 0.08471f
C2828 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.n0 GND 2.01508f
C2829 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6.t0 GND 0.08522f
C2830 a_23031_20174.t2 GND 0.15567f
C2831 a_23031_20174.t1 GND 0.07037f
C2832 a_23031_20174.n0 GND 4.70467f
C2833 a_23031_20174.t3 GND 0.06564f
C2834 a_23031_20174.n1 GND 4.64301f
C2835 a_23031_20174.t0 GND 0.16064f
C2836 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t10 GND 0.3978f
C2837 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t11 GND 0.10005f
C2838 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n0 GND 0.45496f
C2839 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t9 GND 0.10005f
C2840 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n1 GND 0.25833f
C2841 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t8 GND 0.39701f
C2842 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t1 GND 0.11669f
C2843 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t4 GND 0.11669f
C2844 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n2 GND 1.17006f
C2845 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t0 GND 0.11669f
C2846 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t5 GND 0.11669f
C2847 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n3 GND 0.48525f
C2848 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n4 GND 1.72063f
C2849 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t3 GND 0.11669f
C2850 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t6 GND 0.11669f
C2851 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n5 GND 1.17107f
C2852 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t7 GND 0.11669f
C2853 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t2 GND 0.11669f
C2854 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n6 GND 0.48425f
C2855 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n7 GND 1.8498f
C2856 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n8 GND 3.18521f
C2857 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t13 GND 0.40061f
C2858 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t15 GND 0.3992f
C2859 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n9 GND 0.64417f
C2860 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t12 GND 0.40061f
C2861 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.t14 GND 0.3992f
C2862 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n10 GND 0.63961f
C2863 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n11 GND 3.47383f
C2864 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2.n12 GND 0.27271f
C2865 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.t1 GND 0.03836f
C2866 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.t2 GND 0.19594f
C2867 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.n0 GND 4.27168f
C2868 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3.t0 GND 0.19402f
C2869 a_24411_20174.t2 GND 0.17057f
C2870 a_24411_20174.t3 GND 0.06972f
C2871 a_24411_20174.n0 GND 4.89637f
C2872 a_24411_20174.t1 GND 0.16728f
C2873 a_24411_20174.n1 GND 5.40937f
C2874 a_24411_20174.t0 GND 0.0867f
C2875 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t2 GND 0.0125f
C2876 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t1 GND 0.08878f
C2877 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t0 GND 0.0907f
C2878 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.n0 GND 1.58019f
C2879 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t0 GND 0.09594f
C2880 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n0 GND 0.03934f
C2881 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n1 GND 0.08468f
C2882 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n2 GND 0.05622f
C2883 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t1 GND 0.09191f
C2884 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n3 GND 0.01161f
C2885 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t3 GND 0.18837f
C2886 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t6 GND 0.19059f
C2887 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n4 GND 0.90969f
C2888 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t5 GND 0.1906f
C2889 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n5 GND 0.42796f
C2890 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t2 GND 0.18758f
C2891 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n6 GND 1.95827f
C2892 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n7 GND 8.68209f
C2893 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t4 GND 0.18096f
C2894 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.t7 GND 0.17847f
C2895 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n8 GND 1.96854f
C2896 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n9 GND 11.2325f
C2897 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1.n10 GND 0.06052f
C2898 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t0 GND 0.19229f
C2899 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t2 GND 0.22982f
C2900 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t3 GND 0.21285f
C2901 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n0 GND 2.94206f
C2902 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n1 GND 1.71712f
C2903 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t1 GND 0.20585f
C2904 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.t2 GND 0.0362f
C2905 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.t1 GND 0.20214f
C2906 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.n0 GND 4.25884f
C2907 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9.t0 GND 0.20281f
C2908 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.t1 GND -0.0437f
C2909 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.n0 GND -0.90533f
C2910 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10.t0 GND -0.04356f
C2911 a_23049_18133.t5 GND 0.06059f
C2912 a_23049_18133.t1 GND 0.05908f
C2913 a_23049_18133.n0 GND 1.66289f
C2914 a_23049_18133.t3 GND 0.05948f
C2915 a_23049_18133.n1 GND 1.49069f
C2916 a_23049_18133.t2 GND 0.05948f
C2917 a_23049_18133.n2 GND 1.41357f
C2918 a_23049_18133.t4 GND 0.05948f
C2919 a_23049_18133.n3 GND 2.3636f
C2920 a_23049_18133.t0 GND 0.07113f
C2921 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.t2 GND 0.10286f
C2922 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.t1 GND 0.01467f
C2923 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.n0 GND 2.07652f
C2924 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44.t0 GND 0.10595f
C2925 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.t1 GND 0.01522f
C2926 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.t2 GND 0.09452f
C2927 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.n0 GND 1.89603f
C2928 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11.t0 GND 0.09423f
C2929 a_23583_20174.t2 GND 0.13926f
C2930 a_23583_20174.t1 GND 0.17307f
C2931 a_23583_20174.t3 GND 0.07081f
C2932 a_23583_20174.n0 GND 5.33077f
C2933 a_23583_20174.n1 GND 5.29359f
C2934 a_23583_20174.t0 GND 0.0925f
C2935 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t0 GND 0.37557f
C2936 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t3 GND 0.19527f
C2937 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t2 GND 0.19937f
C2938 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n0 GND 1.75815f
C2939 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n1 GND 2.71685f
C2940 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t1 GND 0.19137f
C2941 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n2 GND 0.35177f
C2942 a_34186_8950.t1 GND 0.10046f
C2943 a_34186_8950.t2 GND 0.11818f
C2944 a_34186_8950.n0 GND 5.80655f
C2945 a_34186_8950.t0 GND 0.07481f
C2946 a_28172_6250.t1 GND 0.12364f
C2947 a_28172_6250.t4 GND 0.07206f
C2948 a_28172_6250.n0 GND 4.94854f
C2949 a_28172_6250.t3 GND 0.15859f
C2950 a_28172_6250.n1 GND 4.24803f
C2951 a_28172_6250.t2 GND 0.15202f
C2952 a_28172_6250.n2 GND 4.62506f
C2953 a_28172_6250.t0 GND 0.07206f
C2954 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t3 GND 0.27743f
C2955 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t4 GND 0.28945f
C2956 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t8 GND 0.88849f
C2957 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t6 GND 0.87989f
C2958 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n0 GND 1.08085f
C2959 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t7 GND 0.87989f
C2960 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t9 GND 0.88849f
C2961 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n1 GND 0.72036f
C2962 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n2 GND 0.58652f
C2963 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n3 GND 1.07239f
C2964 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n4 GND 0.80072f
C2965 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t2 GND 0.37408f
C2966 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n5 GND 1.36783f
C2967 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t1 GND 0.28834f
C2968 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n6 GND 1.18764f
C2969 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t5 GND 0.08754f
C2970 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.t0 GND 0.09368f
C2971 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax.n7 GND 0.93685f
C2972 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t2 GND 0.20388f
C2973 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t3 GND 0.19134f
C2974 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n0 GND 1.5154f
C2975 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t0 GND 0.1968f
C2976 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n1 GND 0.75134f
C2977 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t1 GND 0.39307f
C2978 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t1 GND 0.07548f
C2979 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t3 GND 0.07543f
C2980 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n0 GND 0.1418f
C2981 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t5 GND 0.07543f
C2982 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t4 GND 0.28512f
C2983 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t7 GND 0.2877f
C2984 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t10 GND 0.28677f
C2985 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n1 GND 0.35847f
C2986 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t13 GND 0.28766f
C2987 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t6 GND 0.28677f
C2988 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n2 GND 0.35058f
C2989 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n3 GND 0.08769f
C2990 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n4 GND 0.15103f
C2991 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t2 GND 0.28512f
C2992 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t12 GND 0.28766f
C2993 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t8 GND 0.28677f
C2994 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n5 GND 0.35058f
C2995 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t9 GND 0.2877f
C2996 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t11 GND 0.28677f
C2997 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n6 GND 0.35847f
C2998 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n7 GND 0.08769f
C2999 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n8 GND 0.15103f
C3000 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n9 GND 0.1243f
C3001 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n10 GND 0.13769f
C3002 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n11 GND 0.35047f
C3003 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n12 GND 0.26235f
C3004 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t0 GND 0.07543f
C3005 a_19552_8950.t2 GND 0.08071f
C3006 a_19552_8950.t1 GND 0.08167f
C3007 a_19552_8950.n0 GND 5.66782f
C3008 a_19552_8950.t0 GND 0.0698f
C3009 ROUT1.t4 GND 6.96884f
C3010 ROUT1.t2 GND 5.43635f
C3011 ROUT1.n0 GND 3.31329f
C3012 ROUT1.t3 GND 0.07446f
C3013 ROUT1.t1 GND 0.2508f
C3014 ROUT1.n1 GND 2.0531f
C3015 ROUT1.n2 GND 0.43339f
C3016 ROUT1.t0 GND 6.96884f
C3017 ROUT1.t5 GND 5.43635f
C3018 ROUT1.n3 GND 3.14493f
C3019 ROUT1.n4 GND 0.37532f
C3020 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.t1 GND 0.10104f
C3021 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.t2 GND 0.01339f
C3022 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.n0 GND 1.8875f
C3023 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28.t0 GND 0.09807f
C3024 a_33358_8950.t1 GND 0.04502f
C3025 a_33358_8950.t2 GND 0.05347f
C3026 a_33358_8950.n0 GND 2.76188f
C3027 a_33358_8950.t0 GND 0.03963f
C3028 a_27344_6250.t1 GND 0.06897f
C3029 a_27344_6250.t4 GND 0.04091f
C3030 a_27344_6250.n0 GND 2.62657f
C3031 a_27344_6250.t3 GND 0.08929f
C3032 a_27344_6250.n1 GND 2.43648f
C3033 a_27344_6250.t2 GND 0.08534f
C3034 a_27344_6250.n2 GND 2.71152f
C3035 a_27344_6250.t0 GND 0.04091f
C3036 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.t2 GND 0.01445f
C3037 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.t1 GND 0.10131f
C3038 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.n0 GND 1.97942f
C3039 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27.t0 GND 0.10483f
C3040 a_22203_20174.t2 GND 0.17024f
C3041 a_22203_20174.t3 GND 0.07006f
C3042 a_22203_20174.n0 GND 5.08543f
C3043 a_22203_20174.t1 GND 0.05862f
C3044 a_22203_20174.n1 GND 4.26715f
C3045 a_22203_20174.t0 GND 0.14851f
C3046 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t2 GND 0.0223f
C3047 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t0 GND 0.12906f
C3048 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t1 GND 0.42098f
C3049 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.n0 GND 2.85982f
C3050 a_15353_7686.t3 GND 0.03957f
C3051 a_15353_7686.t1 GND 0.04498f
C3052 a_15353_7686.n0 GND 2.05844f
C3053 a_15353_7686.t2 GND 0.04733f
C3054 a_15353_7686.t4 GND 0.03831f
C3055 a_15353_7686.n1 GND 2.62168f
C3056 a_15353_7686.n2 GND 1.51138f
C3057 a_15353_7686.t0 GND 0.03831f
C3058 a_16891_7686.t3 GND 0.08331f
C3059 a_16891_7686.t1 GND 0.09293f
C3060 a_16891_7686.t4 GND 0.07283f
C3061 a_16891_7686.n0 GND 5.53481f
C3062 a_16891_7686.t2 GND 0.07283f
C3063 a_16891_7686.n1 GND 2.64424f
C3064 a_16891_7686.n2 GND 3.92477f
C3065 a_16891_7686.t0 GND 0.07429f
C3066 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t0 GND 0.10561f
C3067 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n0 GND 0.0433f
C3068 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n1 GND 0.09321f
C3069 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n2 GND 0.06188f
C3070 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t1 GND 0.10117f
C3071 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n3 GND 0.01278f
C3072 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t3 GND 0.20879f
C3073 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n4 GND 0.27086f
C3074 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t2 GND 0.20979f
C3075 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n5 GND 0.545f
C3076 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].t4 GND 0.20647f
C3077 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n6 GND 15.6438f
C3078 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4].n7 GND 0.06662f
C3079 top_DAC_0/top_rseg_n_dcell_0.VS1.n0 GND 0.04824f
C3080 top_DAC_0/top_rseg_n_dcell_0.VS1.n1 GND 0.02742f
C3081 top_DAC_0/top_rseg_n_dcell_0.VS1.n2 GND 0.02742f
C3082 top_DAC_0/top_rseg_n_dcell_0.VS1.n3 GND 0.0273f
C3083 top_DAC_0/top_rseg_n_dcell_0.VS1.n4 GND 1.23966f
C3084 top_DAC_0/top_rseg_n_dcell_0.SH[1].t0 GND 0.06573f
C3085 top_DAC_0/top_rseg_n_dcell_0.SH[1].n0 GND 0.02695f
C3086 top_DAC_0/top_rseg_n_dcell_0.SH[1].n1 GND 0.05801f
C3087 top_DAC_0/top_rseg_n_dcell_0.SH[1].n2 GND 0.03851f
C3088 top_DAC_0/top_rseg_n_dcell_0.SH[1].t1 GND 0.06297f
C3089 top_DAC_0/top_rseg_n_dcell_0.SH[1].t2 GND 0.12277f
C3090 top_DAC_0/top_rseg_n_dcell_0.SH[1].t5 GND 0.12226f
C3091 top_DAC_0/top_rseg_n_dcell_0.SH[1].n4 GND 0.24246f
C3092 top_DAC_0/top_rseg_n_dcell_0.SH[1].t3 GND 0.12226f
C3093 top_DAC_0/top_rseg_n_dcell_0.SH[1].n5 GND 0.13493f
C3094 top_DAC_0/top_rseg_n_dcell_0.SH[1].t6 GND 0.12226f
C3095 top_DAC_0/top_rseg_n_dcell_0.SH[1].n6 GND 0.13493f
C3096 top_DAC_0/top_rseg_n_dcell_0.SH[1].t4 GND 0.12226f
C3097 top_DAC_0/top_rseg_n_dcell_0.SH[1].n7 GND 0.14433f
C3098 top_DAC_0/top_rseg_n_dcell_0.SH[1].n8 GND 0.0446f
C3099 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.t1 GND 0.04645f
C3100 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.t2 GND 0.14921f
C3101 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.t0 GND 0.13937f
C3102 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25.n0 GND 2.57872f
C3103 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t0 GND 0.09761f
C3104 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n0 GND 0.04002f
C3105 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n1 GND 0.08615f
C3106 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n2 GND 0.0572f
C3107 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t1 GND 0.09351f
C3108 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n3 GND 0.01181f
C3109 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t10 GND 0.19391f
C3110 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t2 GND 0.19298f
C3111 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n4 GND 0.605f
C3112 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t7 GND 0.19298f
C3113 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n5 GND 0.30296f
C3114 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t4 GND 0.19298f
C3115 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n6 GND 0.30296f
C3116 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t6 GND 0.19298f
C3117 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n7 GND 0.30296f
C3118 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t9 GND 0.19298f
C3119 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n8 GND 0.30296f
C3120 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t5 GND 0.19298f
C3121 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n9 GND 0.30296f
C3122 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t8 GND 0.19298f
C3123 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n10 GND 0.30296f
C3124 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].t3 GND 0.19298f
C3125 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n11 GND 0.24595f
C3126 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n12 GND 15.8955f
C3127 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6].n13 GND 0.06157f
C3128 top_DAC_0/top_rseg_n_dcell_0.SH[4].t0 GND 0.10988f
C3129 top_DAC_0/top_rseg_n_dcell_0.SH[4].n0 GND 0.04505f
C3130 top_DAC_0/top_rseg_n_dcell_0.SH[4].n1 GND 0.09698f
C3131 top_DAC_0/top_rseg_n_dcell_0.SH[4].n2 GND 0.06438f
C3132 top_DAC_0/top_rseg_n_dcell_0.SH[4].t1 GND 0.10526f
C3133 top_DAC_0/top_rseg_n_dcell_0.SH[4].n3 GND 0.0133f
C3134 top_DAC_0/top_rseg_n_dcell_0.SH[4].t5 GND 0.21566f
C3135 top_DAC_0/top_rseg_n_dcell_0.SH[4].t3 GND 0.21482f
C3136 top_DAC_0/top_rseg_n_dcell_0.SH[4].n4 GND 0.41293f
C3137 top_DAC_0/top_rseg_n_dcell_0.SH[4].t6 GND 0.21482f
C3138 top_DAC_0/top_rseg_n_dcell_0.SH[4].n5 GND 0.22937f
C3139 top_DAC_0/top_rseg_n_dcell_0.SH[4].t4 GND 0.21482f
C3140 top_DAC_0/top_rseg_n_dcell_0.SH[4].n6 GND 0.22937f
C3141 top_DAC_0/top_rseg_n_dcell_0.SH[4].t2 GND 0.21482f
C3142 top_DAC_0/top_rseg_n_dcell_0.SH[4].n7 GND 0.24931f
C3143 top_DAC_0/top_rseg_n_dcell_0.SH[4].n8 GND 0.07456f
C3144 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t1 GND 0.21159f
C3145 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t2 GND 0.22082f
C3146 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t3 GND 0.21829f
C3147 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n0 GND 2.05618f
C3148 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n1 GND 0.68941f
C3149 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t0 GND 0.43691f
C3150 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t3 GND 0.04207f
C3151 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t0 GND 0.15904f
C3152 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t5 GND 0.0423f
C3153 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t4 GND 0.04183f
C3154 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n0 GND 0.16659f
C3155 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t9 GND 0.15996f
C3156 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n1 GND 0.18631f
C3157 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t13 GND 0.15996f
C3158 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n2 GND 0.10596f
C3159 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t6 GND 0.16046f
C3160 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t8 GND 0.15996f
C3161 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n3 GND 0.19556f
C3162 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n4 GND 0.04891f
C3163 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n5 GND 0.08386f
C3164 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t2 GND 0.15904f
C3165 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t12 GND 0.16048f
C3166 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t7 GND 0.15996f
C3167 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n6 GND 0.19996f
C3168 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t10 GND 0.16046f
C3169 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t11 GND 0.15996f
C3170 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n7 GND 0.19556f
C3171 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n8 GND 0.04891f
C3172 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n9 GND 0.08386f
C3173 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n10 GND 0.06653f
C3174 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t1 GND 0.04207f
C3175 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n11 GND 0.14113f
C3176 top_DAC_0/top_rseg_n_dcell_0.VH3.t4 GND 0.0194f
C3177 top_DAC_0/top_rseg_n_dcell_0.VH3.t3 GND 0.02035f
C3178 top_DAC_0/top_rseg_n_dcell_0.VH3.n1 GND 1.19499f
C3179 top_DAC_0/top_rseg_n_dcell_0.VH3.t1 GND 0.01939f
C3180 top_DAC_0/top_rseg_n_dcell_0.VH3.t2 GND 0.01934f
C3181 top_DAC_0/top_rseg_n_dcell_0.VH3.n2 GND 0.11763f
C3182 top_DAC_0/top_rseg_n_dcell_0.VH3.t0 GND 0.01934f
C3183 top_DAC_0/top_rseg_n_dcell_0.VH3.n3 GND 0.13268f
C3184 a_8051_10107.t12 GND 0.01041f
C3185 a_8051_10107.t15 GND 0.01041f
C3186 a_8051_10107.t0 GND 0.01041f
C3187 a_8051_10107.n0 GND 0.02413f
C3188 a_8051_10107.t2 GND 0.01041f
C3189 a_8051_10107.t13 GND 0.01041f
C3190 a_8051_10107.n1 GND 0.02413f
C3191 a_8051_10107.n2 GND 0.17752f
C3192 a_8051_10107.t6 GND 0.02333f
C3193 a_8051_10107.t10 GND 0.02333f
C3194 a_8051_10107.n3 GND 0.35392f
C3195 a_8051_10107.n4 GND 0.34189f
C3196 a_8051_10107.t4 GND 0.0233f
C3197 a_8051_10107.n5 GND 0.09101f
C3198 a_8051_10107.t5 GND 0.0233f
C3199 a_8051_10107.n6 GND 0.09101f
C3200 a_8051_10107.n7 GND 0.08577f
C3201 a_8051_10107.t8 GND 0.02333f
C3202 a_8051_10107.t11 GND 0.02333f
C3203 a_8051_10107.n8 GND 0.21448f
C3204 a_8051_10107.t7 GND 0.02333f
C3205 a_8051_10107.t9 GND 0.02333f
C3206 a_8051_10107.n9 GND 0.29964f
C3207 a_8051_10107.n10 GND 0.38663f
C3208 a_8051_10107.n11 GND 0.63923f
C3209 a_8051_10107.n12 GND 0.07503f
C3210 a_8051_10107.t14 GND 0.01041f
C3211 a_8051_10107.t1 GND 0.01041f
C3212 a_8051_10107.n13 GND 0.02413f
C3213 a_8051_10107.n14 GND 0.17752f
C3214 a_8051_10107.n15 GND 0.02413f
C3215 a_8051_10107.t3 GND 0.01041f
C3216 a_28882_6250.t1 GND 0.14276f
C3217 a_28882_6250.t4 GND 0.08249f
C3218 a_28882_6250.n0 GND 4.59159f
C3219 a_28882_6250.t3 GND 0.15799f
C3220 a_28882_6250.n1 GND 4.32313f
C3221 a_28882_6250.t2 GND 0.17484f
C3222 a_28882_6250.n2 GND 6.44471f
C3223 a_28882_6250.t0 GND 0.08249f
C3224 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t0 GND 0.08516f
C3225 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n0 GND 0.03492f
C3226 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n1 GND 0.07516f
C3227 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n2 GND 0.0499f
C3228 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t1 GND 0.08158f
C3229 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n3 GND 0.0103f
C3230 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t3 GND 0.16917f
C3231 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t12 GND 0.16836f
C3232 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n4 GND 0.52781f
C3233 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t2 GND 0.16836f
C3234 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n5 GND 0.26431f
C3235 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t6 GND 0.16836f
C3236 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n6 GND 0.26431f
C3237 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t14 GND 0.16836f
C3238 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n7 GND 0.26431f
C3239 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t16 GND 0.16836f
C3240 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n8 GND 0.26431f
C3241 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t11 GND 0.16836f
C3242 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n9 GND 0.26431f
C3243 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t13 GND 0.16649f
C3244 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t4 GND 0.16917f
C3245 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t5 GND 0.16969f
C3246 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t17 GND 0.16882f
C3247 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n10 GND 0.57115f
C3248 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t15 GND 0.16882f
C3249 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n11 GND 0.28601f
C3250 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t7 GND 0.16882f
C3251 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n12 GND 0.28601f
C3252 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t10 GND 0.16882f
C3253 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n13 GND 0.28601f
C3254 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t9 GND 0.16882f
C3255 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n14 GND 0.28601f
C3256 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n15 GND 0.43945f
C3257 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.t8 GND 0.16649f
C3258 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n16 GND 0.42862f
C3259 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n17 GND 0.20782f
C3260 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n18 GND 13.6678f
C3261 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n19 GND 13.4839f
C3262 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1.n20 GND 0.06924f
C3263 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t2 GND 0.02428f
C3264 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t3 GND 0.02428f
C3265 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 GND 0.0579f
C3266 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y GND 0.18773f
C3267 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 GND 0.11375f
C3268 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t7 GND 0.05811f
C3269 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t11 GND 0.03424f
C3270 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t6 GND 0.05811f
C3271 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t10 GND 0.03424f
C3272 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 GND 0.0975f
C3273 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 GND 0.14465f
C3274 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 GND 0.04362f
C3275 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t9 GND 0.06176f
C3276 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t5 GND 0.03854f
C3277 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 GND 0.12163f
C3278 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.B GND 0.01494f
C3279 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 GND 0.05564f
C3280 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t12 GND 0.06176f
C3281 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t8 GND 0.03854f
C3282 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 GND 0.12159f
C3283 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.B GND 0.01532f
C3284 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 GND 0.04107f
C3285 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 GND 0.63673f
C3286 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[0] GND 2.63598f
C3287 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t4 GND 0.23379f
C3288 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 GND 10.3706f
C3289 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 GND 2.64516f
C3290 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 GND 0.02673f
C3291 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 GND 0.03539f
C3292 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t0 GND 0.03736f
C3293 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t1 GND 0.03736f
C3294 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 GND 0.08204f
C3295 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.t2 GND 0.01319f
C3296 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.t0 GND 0.03696f
C3297 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.t1 GND 0.0369f
C3298 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10.n0 GND 0.66059f
C3299 a_30332_7686.t1 GND 0.0892f
C3300 a_30332_7686.t3 GND 0.09588f
C3301 a_30332_7686.n0 GND 3.63616f
C3302 a_30332_7686.t4 GND 0.07875f
C3303 a_30332_7686.n1 GND 2.9429f
C3304 a_30332_7686.t2 GND 0.14222f
C3305 a_30332_7686.n2 GND 5.73614f
C3306 a_30332_7686.t0 GND 0.07875f
C3307 a_21651_20174.t2 GND 0.21223f
C3308 a_21651_20174.t3 GND 0.08827f
C3309 a_21651_20174.n0 GND 6.60332f
C3310 a_21651_20174.t1 GND 0.0607f
C3311 a_21651_20174.n1 GND 4.57762f
C3312 a_21651_20174.t0 GND 0.15786f
C3313 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t0 GND 0.01293f
C3314 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t2 GND 0.10101f
C3315 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t1 GND 0.09801f
C3316 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.n0 GND 1.62769f
C3317 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.t1 GND 0.0341f
C3318 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.t0 GND 0.12376f
C3319 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.t2 GND 0.36301f
C3320 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8.n0 GND 2.62716f
C3321 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t1 GND 0.06182f
C3322 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t4 GND 0.21263f
C3323 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[3] GND 3.59225f
C3324 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[3] GND 0.2209f
C3325 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t3 GND 0.04704f
C3326 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t5 GND 0.02938f
C3327 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 GND 0.08811f
C3328 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 GND 0.02491f
C3329 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 GND 0.32297f
C3330 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 GND 0.16531f
C3331 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y GND 0.14996f
C3332 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 GND 0.02367f
C3333 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t2 GND 0.02839f
C3334 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t0 GND 0.02839f
C3335 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 GND 0.08229f
C3336 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 GND 0.01239f
C3337 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t3 GND 0.01854f
C3338 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t7 GND 0.01854f
C3339 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n0 GND 0.04373f
C3340 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t9 GND 0.01854f
C3341 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t1 GND 0.01854f
C3342 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n1 GND 0.04396f
C3343 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t0 GND 0.01854f
C3344 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t8 GND 0.01854f
C3345 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n2 GND 0.04396f
C3346 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n3 GND 0.25242f
C3347 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t4 GND 0.07589f
C3348 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t5 GND 0.0695f
C3349 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n4 GND 1.46047f
C3350 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n5 GND 0.06518f
C3351 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t6 GND 0.01854f
C3352 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t2 GND 0.01854f
C3353 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n6 GND 0.04396f
C3354 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n7 GND 0.13765f
C3355 a_14672_18696.t2 GND 0.0346f
C3356 a_14672_18696.t1 GND 0.03023f
C3357 a_14672_18696.t3 GND 0.02819f
C3358 a_14672_18696.n0 GND 0.98182f
C3359 a_14672_18696.n1 GND 1.49663f
C3360 a_14672_18696.t0 GND 0.02853f
C3361 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.t1 GND 0.11065f
C3362 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.t2 GND 0.10704f
C3363 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.n0 GND 2.06692f
C3364 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37.t0 GND 0.0154f
C3365 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.t1 GND 0.04652f
C3366 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.t0 GND 0.13968f
C3367 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.t2 GND 0.13957f
C3368 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57.n0 GND 2.57959f
C3369 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.t2 GND 0.09431f
C3370 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.t1 GND 0.0907f
C3371 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.n0 GND 1.89944f
C3372 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5.t0 GND 0.01555f
C3373 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t18 GND 0.07931f
C3374 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t23 GND 0.07931f
C3375 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n0 GND 0.18708f
C3376 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t20 GND 0.07931f
C3377 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t17 GND 0.07931f
C3378 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n1 GND 0.18806f
C3379 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t22 GND 0.07931f
C3380 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t19 GND 0.07931f
C3381 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n2 GND 0.18806f
C3382 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t16 GND 0.07931f
C3383 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t21 GND 0.07931f
C3384 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n3 GND 0.18806f
C3385 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n4 GND 1.07994f
C3386 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t14 GND 0.19984f
C3387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t12 GND 0.176f
C3388 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t2 GND 0.176f
C3389 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n5 GND 0.72684f
C3390 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n6 GND 2.09379f
C3391 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t9 GND 0.176f
C3392 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t0 GND 0.176f
C3393 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n7 GND 0.72829f
C3394 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n8 GND 1.44342f
C3395 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t7 GND 0.176f
C3396 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t11 GND 0.176f
C3397 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n9 GND 0.72829f
C3398 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n10 GND 0.60469f
C3399 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t1 GND 0.18546f
C3400 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n11 GND 0.5189f
C3401 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t15 GND 0.19033f
C3402 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t4 GND 0.176f
C3403 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t13 GND 0.176f
C3404 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n12 GND 0.72829f
C3405 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n13 GND 1.0751f
C3406 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t6 GND 0.176f
C3407 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t8 GND 0.176f
C3408 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n14 GND 0.72829f
C3409 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n15 GND 1.44342f
C3410 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t5 GND 0.176f
C3411 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t10 GND 0.176f
C3412 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n16 GND 0.72684f
C3413 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n17 GND 1.42725f
C3414 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t3 GND 0.18546f
C3415 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n18 GND 0.69316f
C3416 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n19 GND 1.65076f
C3417 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n20 GND 0.36304f
C3418 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n21 GND 0.58892f
C3419 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t4 GND 0.09798f
C3420 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t7 GND 0.09517f
C3421 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n0 GND 1.57121f
C3422 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t5 GND 0.09798f
C3423 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t3 GND 0.09517f
C3424 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n1 GND 0.98853f
C3425 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n2 GND 0.81058f
C3426 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t1 GND 0.09798f
C3427 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t0 GND 0.09517f
C3428 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n3 GND 1.25415f
C3429 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t2 GND 0.09798f
C3430 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t6 GND 0.09517f
C3431 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n4 GND 1.30559f
C3432 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n5 GND 0.68388f
C3433 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n6 GND 1.49193f
C3434 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t10 GND 0.09131f
C3435 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t9 GND 0.09131f
C3436 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n7 GND 0.60876f
C3437 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t15 GND 0.09131f
C3438 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t11 GND 0.09131f
C3439 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n8 GND 0.63869f
C3440 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n9 GND 1.68727f
C3441 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t13 GND 0.09131f
C3442 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t12 GND 0.09131f
C3443 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n10 GND 0.81419f
C3444 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t8 GND 0.09131f
C3445 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t14 GND 0.09131f
C3446 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n11 GND 0.48631f
C3447 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n12 GND 1.56335f
C3448 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n13 GND 1.03015f
C3449 a_14055_6250.t4 GND 0.09741f
C3450 a_14055_6250.t3 GND 0.09544f
C3451 a_14055_6250.t1 GND 0.07626f
C3452 a_14055_6250.n0 GND 4.32003f
C3453 a_14055_6250.t2 GND 0.11145f
C3454 a_14055_6250.n1 GND 4.74566f
C3455 a_14055_6250.n2 GND 5.27749f
C3456 a_14055_6250.t0 GND 0.07626f
C3457 a_20823_20174.t3 GND 0.15734f
C3458 a_20823_20174.t1 GND 0.05584f
C3459 a_20823_20174.n0 GND 4.21706f
C3460 a_20823_20174.t2 GND 0.05584f
C3461 a_20823_20174.n1 GND 0.59217f
C3462 a_20823_20174.t4 GND 0.07011f
C3463 a_20823_20174.n2 GND 4.88166f
C3464 a_20823_20174.t0 GND 0.16998f
C3465 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t2 GND 0.01248f
C3466 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t1 GND 0.09426f
C3467 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t0 GND 0.09768f
C3468 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.n0 GND 1.54809f
C3469 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t0 GND 0.07332f
C3470 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n0 GND 0.03006f
C3471 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n1 GND 0.06471f
C3472 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n2 GND 0.04296f
C3473 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t1 GND 0.07024f
C3474 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t2 GND 0.15352f
C3475 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t3 GND 0.14496f
C3476 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n4 GND 0.17762f
C3477 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t11 GND 0.14496f
C3478 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n5 GND 0.22757f
C3479 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t7 GND 0.14496f
C3480 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n6 GND 0.22757f
C3481 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t4 GND 0.14496f
C3482 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n7 GND 0.22757f
C3483 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t14 GND 0.14496f
C3484 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n8 GND 0.22757f
C3485 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t17 GND 0.14496f
C3486 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n9 GND 0.22757f
C3487 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t13 GND 0.14565f
C3488 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n10 GND 0.37838f
C3489 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t10 GND 0.14335f
C3490 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n11 GND 2.00631f
C3491 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n12 GND 2.11515f
C3492 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t8 GND 0.14565f
C3493 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n13 GND 0.33941f
C3494 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t20 GND 0.14335f
C3495 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n14 GND 2.10313f
C3496 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n15 GND 7.38065f
C3497 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t6 GND 0.13868f
C3498 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t9 GND 0.13798f
C3499 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n16 GND 0.44941f
C3500 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t5 GND 0.13798f
C3501 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n17 GND 0.22506f
C3502 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t16 GND 0.13798f
C3503 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n18 GND 0.22506f
C3504 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t19 GND 0.13798f
C3505 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n19 GND 0.22506f
C3506 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t18 GND 0.13815f
C3507 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t15 GND 0.13798f
C3508 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n20 GND 0.20036f
C3509 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n21 GND 0.1515f
C3510 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.t12 GND 0.13639f
C3511 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n22 GND 2.01789f
C3512 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n23 GND 8.92053f
C3513 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3.n24 GND 0.04625f
C3514 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t1 GND 0.07769f
C3515 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t2 GND 0.03615f
C3516 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t4 GND 0.02256f
C3517 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n0 GND 0.07188f
C3518 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t5 GND 0.0362f
C3519 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t3 GND 0.0226f
C3520 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n1 GND 0.06891f
C3521 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n2 GND 0.02012f
C3522 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n3 GND 4.68779f
C3523 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n4 GND 0.107f
C3524 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n5 GND 0.02567f
C3525 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t0 GND 0.05407f
C3526 a_30608_7686.t1 GND 0.0933f
C3527 a_30608_7686.t2 GND 0.08812f
C3528 a_30608_7686.n0 GND 3.52034f
C3529 a_30608_7686.t4 GND 0.07942f
C3530 a_30608_7686.n1 GND 2.88984f
C3531 a_30608_7686.t3 GND 0.14424f
C3532 a_30608_7686.n2 GND 5.80531f
C3533 a_30608_7686.t0 GND 0.07942f
C3534 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t18 GND 0.39601f
C3535 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t1 GND 0.08658f
C3536 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t0 GND 0.10174f
C3537 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n0 GND 0.56019f
C3538 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n1 GND 0.44593f
C3539 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t3 GND 0.40442f
C3540 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t15 GND 0.40271f
C3541 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n2 GND 0.89528f
C3542 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n3 GND 0.66573f
C3543 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t6 GND 0.12379f
C3544 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t14 GND 0.12172f
C3545 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n4 GND 6.7007f
C3546 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t19 GND 0.12376f
C3547 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t20 GND 0.12314f
C3548 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n5 GND 0.40108f
C3549 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t21 GND 0.12314f
C3550 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n6 GND 0.20085f
C3551 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t24 GND 0.12314f
C3552 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n7 GND 0.20085f
C3553 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t2 GND 0.12314f
C3554 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n8 GND 0.20085f
C3555 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t5 GND 0.12314f
C3556 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n9 GND 0.20085f
C3557 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t23 GND 0.12314f
C3558 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n10 GND 0.20085f
C3559 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t11 GND 0.12172f
C3560 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t22 GND 0.12376f
C3561 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t8 GND 0.12418f
C3562 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t13 GND 0.1235f
C3563 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n11 GND 0.43438f
C3564 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t12 GND 0.1235f
C3565 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n12 GND 0.21753f
C3566 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t9 GND 0.1235f
C3567 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n13 GND 0.21753f
C3568 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t7 GND 0.1235f
C3569 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n14 GND 0.21753f
C3570 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t4 GND 0.1235f
C3571 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n15 GND 0.21753f
C3572 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n16 GND 0.33544f
C3573 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t10 GND 0.12172f
C3574 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n17 GND 0.41895f
C3575 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n18 GND 0.42347f
C3576 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n19 GND 0.09724f
C3577 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n20 GND 11.1294f
C3578 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t16 GND 0.22885f
C3579 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].t17 GND 0.12695f
C3580 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n21 GND 0.19942f
C3581 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n22 GND 0.03481f
C3582 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2].n23 GND 0.27626f
C3583 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.t1 GND 0.08527f
C3584 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.t2 GND 0.08305f
C3585 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.n0 GND 1.91518f
C3586 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7.t0 GND 0.01651f
C3587 a_34856_8950.t1 GND 0.10872f
C3588 a_34856_8950.t2 GND 0.13049f
C3589 a_34856_8950.n0 GND 6.09434f
C3590 a_34856_8950.t0 GND 0.06644f
C3591 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t3 GND 0.038f
C3592 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t2 GND 0.038f
C3593 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 GND 0.08345f
C3594 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y GND 0.19095f
C3595 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 GND 0.036f
C3596 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t4 GND 0.70975f
C3597 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 GND 14.2799f
C3598 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t0 GND 0.0247f
C3599 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t1 GND 0.0247f
C3600 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 GND 0.05889f
C3601 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 GND 0.1157f
C3602 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t2 GND 0.0261f
C3603 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t3 GND 0.0261f
C3604 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 GND 0.06224f
C3605 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y GND 0.20181f
C3606 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 GND 0.12228f
C3607 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t6 GND 0.06247f
C3608 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t4 GND 0.03681f
C3609 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t5 GND 0.06247f
C3610 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t7 GND 0.03681f
C3611 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 GND 0.10482f
C3612 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 GND 0.1555f
C3613 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.A GND 0.01041f
C3614 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 GND 0.04689f
C3615 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t8 GND 0.57365f
C3616 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 GND 15.4363f
C3617 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 GND 0.02873f
C3618 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 GND 0.03805f
C3619 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t0 GND 0.04016f
C3620 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t1 GND 0.04016f
C3621 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 GND 0.0882f
C3622 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t3 GND 0.13497f
C3623 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t4 GND 0.18291f
C3624 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n0 GND 0.62616f
C3625 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t2 GND 0.04322f
C3626 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t12 GND 0.16799f
C3627 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t6 GND 0.16762f
C3628 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n1 GND 0.19518f
C3629 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t7 GND 0.16762f
C3630 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n2 GND 0.09252f
C3631 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t15 GND 0.16799f
C3632 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t14 GND 0.16762f
C3633 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n3 GND 0.19518f
C3634 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t8 GND 0.16762f
C3635 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n4 GND 0.09252f
C3636 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n5 GND 0.08905f
C3637 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t13 GND 0.16799f
C3638 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t9 GND 0.16762f
C3639 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n6 GND 0.19518f
C3640 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t10 GND 0.16762f
C3641 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n7 GND 0.09252f
C3642 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t17 GND 0.16799f
C3643 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t16 GND 0.16762f
C3644 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n8 GND 0.19518f
C3645 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t11 GND 0.16762f
C3646 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n9 GND 0.09252f
C3647 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n10 GND 0.21323f
C3648 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t1 GND 0.04581f
C3649 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t0 GND 0.04261f
C3650 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n11 GND 0.29976f
C3651 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n12 GND 0.21959f
C3652 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n13 GND 0.28569f
C3653 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.t5 GND 0.06288f
C3654 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx.n14 GND 0.51077f
C3655 a_29434_6250.t1 GND 0.07592f
C3656 a_29434_6250.t4 GND 0.04358f
C3657 a_29434_6250.n0 GND 2.54446f
C3658 a_29434_6250.t3 GND 0.06837f
C3659 a_29434_6250.n1 GND 1.92423f
C3660 a_29434_6250.t2 GND 0.09262f
C3661 a_29434_6250.n2 GND 3.30724f
C3662 a_29434_6250.t0 GND 0.04358f
C3663 a_35132_8950.t1 GND 0.05535f
C3664 a_35132_8950.t2 GND 0.06636f
C3665 a_35132_8950.n0 GND 3.04622f
C3666 a_35132_8950.t0 GND 0.03208f
C3667 top_DAC_0/top_final_switch_0.VOUT[2].t3 GND 0.01008f
C3668 top_DAC_0/top_final_switch_0.VOUT[2].t2 GND 0.01008f
C3669 top_DAC_0/top_final_switch_0.VOUT[2].n0 GND 0.02294f
C3670 top_DAC_0/top_final_switch_0.VOUT[2].t0 GND 0.01008f
C3671 top_DAC_0/top_final_switch_0.VOUT[2].t1 GND 0.01008f
C3672 top_DAC_0/top_final_switch_0.VOUT[2].n1 GND 0.02395f
C3673 top_DAC_0/top_final_switch_0.VOUT[2].n2 GND 1.36615f
C3674 top_DAC_0/top_final_switch_0.VOUT[2].t8 GND 0.93759f
C3675 top_DAC_0/top_final_switch_0.VOUT[2].t9 GND 0.93174f
C3676 top_DAC_0/top_final_switch_0.VOUT[2].n3 GND 1.55465f
C3677 top_DAC_0/top_final_switch_0.VOUT[2].t6 GND 0.93236f
C3678 top_DAC_0/top_final_switch_0.VOUT[2].t11 GND 0.93066f
C3679 top_DAC_0/top_final_switch_0.VOUT[2].n4 GND 1.20046f
C3680 top_DAC_0/top_final_switch_0.VOUT[2].n5 GND 0.82741f
C3681 top_DAC_0/top_final_switch_0.VOUT[2].t4 GND 0.38306f
C3682 top_DAC_0/top_final_switch_0.VOUT[2].t10 GND 0.38121f
C3683 top_DAC_0/top_final_switch_0.VOUT[2].n6 GND 1.01242f
C3684 top_DAC_0/top_final_switch_0.VOUT[2].t5 GND 0.38937f
C3685 top_DAC_0/top_final_switch_0.VOUT[2].t7 GND 0.38279f
C3686 top_DAC_0/top_final_switch_0.VOUT[2].n7 GND 1.1277f
C3687 top_DAC_0/top_final_switch_0.VOUT[2].n8 GND 0.54763f
C3688 top_DAC_0/top_final_switch_0.VOUT[2].n9 GND 1.78948f
C3689 top_DAC_0/top_final_switch_0.VOUT[2].n10 GND 0.2511f
C3690 a_23859_20174.t2 GND 0.06748f
C3691 a_23859_20174.t1 GND 0.08959f
C3692 a_23859_20174.t3 GND 0.03679f
C3693 a_23859_20174.n0 GND 2.82037f
C3694 a_23859_20174.n1 GND 2.83277f
C3695 a_23859_20174.t0 GND 0.053f
C3696 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t10 GND 0.57173f
C3697 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t12 GND 0.57394f
C3698 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t14 GND 0.57311f
C3699 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n0 GND 0.57028f
C3700 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t13 GND 0.57394f
C3701 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t15 GND 0.57311f
C3702 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n1 GND 0.5671f
C3703 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n2 GND 1.86177f
C3704 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n3 GND 2.60622f
C3705 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t11 GND 0.17341f
C3706 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n4 GND 0.23921f
C3707 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t0 GND 0.02203f
C3708 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t2 GND 0.02203f
C3709 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n5 GND 0.45415f
C3710 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n6 GND 0.47964f
C3711 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t1 GND 0.02201f
C3712 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n7 GND 0.07372f
C3713 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t5 GND 0.02201f
C3714 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n8 GND 0.07372f
C3715 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n9 GND 0.32363f
C3716 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t4 GND 0.02203f
C3717 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t3 GND 0.02203f
C3718 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n10 GND 0.45415f
C3719 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n11 GND 0.47964f
C3720 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t6 GND 0.02201f
C3721 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n12 GND 0.07372f
C3722 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t7 GND 0.02201f
C3723 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n13 GND 0.07372f
C3724 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n14 GND 0.19305f
C3725 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n15 GND 0.64379f
C3726 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n16 GND 0.22337f
C3727 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t9 GND 0.17341f
C3728 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.n17 GND 0.2098f
C3729 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1.t8 GND 0.57148f
C3730 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t2 GND 0.15112f
C3731 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n0 GND 0.31314f
C3732 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t3 GND 0.03061f
C3733 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n1 GND 0.09861f
C3734 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t15 GND 0.19802f
C3735 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n3 GND 0.13878f
C3736 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t11 GND 0.19802f
C3737 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n4 GND 0.14564f
C3738 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t6 GND 0.19802f
C3739 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n5 GND 0.14564f
C3740 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t9 GND 0.19802f
C3741 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n6 GND 0.10675f
C3742 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t16 GND 0.19802f
C3743 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n7 GND 0.10675f
C3744 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t10 GND 0.19802f
C3745 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n8 GND 0.14564f
C3746 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t13 GND 0.19802f
C3747 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n9 GND 0.14564f
C3748 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t7 GND 0.19802f
C3749 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n10 GND 0.14408f
C3750 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t8 GND 0.19802f
C3751 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n11 GND 0.10675f
C3752 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t17 GND 0.19802f
C3753 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n12 GND 0.14564f
C3754 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t14 GND 0.19802f
C3755 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n13 GND 0.14564f
C3756 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t12 GND 0.19802f
C3757 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n14 GND 0.10859f
C3758 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n15 GND 0.39639f
C3759 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n16 GND 0.8517f
C3760 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t1 GND 0.03061f
C3761 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n17 GND 0.08691f
C3762 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t0 GND 0.15112f
C3763 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n18 GND 0.11384f
C3764 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n19 GND 0.67032f
C3765 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t4 GND 0.09915f
C3766 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n20 GND 0.53323f
C3767 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t5 GND 0.09577f
C3768 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n21 GND 0.14399f
C3769 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t2 GND 0.09331f
C3770 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t4 GND 0.09112f
C3771 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n0 GND 1.44549f
C3772 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t7 GND 0.09331f
C3773 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t3 GND 0.09112f
C3774 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n1 GND 1.29109f
C3775 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n2 GND 1.38567f
C3776 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t5 GND 0.09331f
C3777 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t6 GND 0.09112f
C3778 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n3 GND 1.13504f
C3779 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t1 GND 0.09331f
C3780 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t0 GND 0.09112f
C3781 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n4 GND 1.60154f
C3782 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n5 GND 1.29052f
C3783 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n6 GND 1.36983f
C3784 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t10 GND 0.08941f
C3785 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t9 GND 0.08941f
C3786 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n7 GND 0.62001f
C3787 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t12 GND 0.08941f
C3788 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t15 GND 0.08941f
C3789 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n8 GND 0.95504f
C3790 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n9 GND 2.44269f
C3791 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t13 GND 0.08941f
C3792 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t8 GND 0.08941f
C3793 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n10 GND 0.83514f
C3794 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t14 GND 0.08941f
C3795 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t11 GND 0.08941f
C3796 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n11 GND 0.7235f
C3797 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n12 GND 2.41198f
C3798 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n13 GND 0.91107f
C3799 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t3 GND 0.04627f
C3800 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t12 GND 0.04627f
C3801 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n0 GND 0.10915f
C3802 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t15 GND 0.04627f
C3803 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t0 GND 0.04627f
C3804 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n1 GND 0.10972f
C3805 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t2 GND 0.04627f
C3806 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t13 GND 0.04627f
C3807 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n2 GND 0.10972f
C3808 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n3 GND 0.63006f
C3809 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t5 GND 0.10271f
C3810 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t6 GND 0.10271f
C3811 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n4 GND 0.61687f
C3812 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t7 GND 0.10271f
C3813 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t10 GND 0.10271f
C3814 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n5 GND 0.42623f
C3815 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n6 GND 0.92706f
C3816 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t9 GND 0.10271f
C3817 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t11 GND 0.10271f
C3818 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n7 GND 0.61598f
C3819 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t8 GND 0.10271f
C3820 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t4 GND 0.10271f
C3821 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n8 GND 0.42711f
C3822 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n9 GND 0.68929f
C3823 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n10 GND 1.50345f
C3824 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n11 GND 0.20317f
C3825 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t14 GND 0.04627f
C3826 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t1 GND 0.04627f
C3827 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n12 GND 0.10972f
C3828 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n13 GND 0.34359f
C3829 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t9 GND 0.04528f
C3830 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t8 GND 0.04528f
C3831 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n0 GND 0.09481f
C3832 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t11 GND 0.17013f
C3833 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t19 GND 0.04528f
C3834 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t22 GND 0.04528f
C3835 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n1 GND 0.09481f
C3836 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t21 GND 0.17013f
C3837 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t12 GND 0.04528f
C3838 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t23 GND 0.04528f
C3839 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n2 GND 0.09481f
C3840 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t13 GND 0.17013f
C3841 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t15 GND 0.04528f
C3842 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t17 GND 0.04528f
C3843 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n3 GND 0.09481f
C3844 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t18 GND 0.17013f
C3845 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t27 GND 0.04528f
C3846 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t24 GND 0.04528f
C3847 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n4 GND 0.09481f
C3848 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t26 GND 0.21091f
C3849 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n5 GND 0.81416f
C3850 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n6 GND 0.10911f
C3851 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t25 GND 0.17019f
C3852 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n7 GND 0.40872f
C3853 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n8 GND 0.53208f
C3854 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n9 GND 0.4693f
C3855 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n10 GND 0.10911f
C3856 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t16 GND 0.17019f
C3857 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n11 GND 0.40872f
C3858 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n12 GND 0.53208f
C3859 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n13 GND 0.4693f
C3860 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n14 GND 0.10911f
C3861 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t14 GND 0.17019f
C3862 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n15 GND 0.40872f
C3863 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n16 GND 0.53208f
C3864 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n17 GND 0.4693f
C3865 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n18 GND 0.10911f
C3866 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t20 GND 0.17019f
C3867 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n19 GND 0.40872f
C3868 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n20 GND 0.53208f
C3869 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n21 GND 0.4683f
C3870 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n22 GND 0.10549f
C3871 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t10 GND 0.17019f
C3872 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n23 GND 1.07705f
C3873 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t4 GND 0.10478f
C3874 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n24 GND 1.33842f
C3875 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t2 GND 0.02415f
C3876 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t6 GND 0.02415f
C3877 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n25 GND 0.05228f
C3878 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t3 GND 0.02415f
C3879 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t7 GND 0.02415f
C3880 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n26 GND 0.0573f
C3881 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t0 GND 0.02415f
C3882 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t1 GND 0.02415f
C3883 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n27 GND 0.05228f
C3884 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n28 GND 0.6261f
C3885 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n29 GND 0.56497f
C3886 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t5 GND 0.10957f
C3887 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n30 GND 0.84934f
C3888 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t2 GND 0.02214f
C3889 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t9 GND 0.02214f
C3890 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n0 GND 0.05223f
C3891 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t8 GND 0.02214f
C3892 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t1 GND 0.02214f
C3893 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n1 GND 0.0525f
C3894 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t7 GND 0.02214f
C3895 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t0 GND 0.02214f
C3896 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n2 GND 0.0525f
C3897 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t3 GND 0.02214f
C3898 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t6 GND 0.02214f
C3899 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n3 GND 0.0525f
C3900 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n4 GND 0.3015f
C3901 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t4 GND 0.07201f
C3902 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t5 GND 0.06819f
C3903 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n5 GND 1.29541f
C3904 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n6 GND 0.07426f
C3905 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n7 GND 0.16442f
C3906 a_28606_6250.t1 GND 0.12539f
C3907 a_28606_6250.t4 GND 0.07275f
C3908 a_28606_6250.n0 GND 3.93804f
C3909 a_28606_6250.t3 GND 0.15297f
C3910 a_28606_6250.n1 GND 4.11942f
C3911 a_28606_6250.t2 GND 0.15386f
C3912 a_28606_6250.n2 GND 5.76483f
C3913 a_28606_6250.t0 GND 0.07275f
C3914 a_34304_8950.t1 GND 0.10705f
C3915 a_34304_8950.t2 GND 0.12718f
C3916 a_34304_8950.n0 GND 6.19294f
C3917 a_34304_8950.t0 GND 0.07284f
C3918 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y GND 0.56561f
C3919 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t0 GND 0.10003f
C3920 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n0 GND 0.04101f
C3921 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n1 GND 0.08829f
C3922 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n2 GND 0.05861f
C3923 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t1 GND 0.09583f
C3924 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n3 GND 0.0121f
C3925 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t5 GND 0.19162f
C3926 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t4 GND 0.19796f
C3927 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n4 GND 0.77307f
C3928 top_DAC_0/top_final_switch_0.bb[0] GND 1.02307f
C3929 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t3 GND 0.27685f
C3930 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n5 GND 10.3749f
C3931 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.bb[0] GND 0.20519f
C3932 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t7 GND 0.18607f
C3933 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n6 GND 1.91143f
C3934 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n7 GND 12.3818f
C3935 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.bb[0] GND 3.51124f
C3936 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUTB GND 0.35266f
C3937 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t2 GND 0.34983f
C3938 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.t6 GND 0.19406f
C3939 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n8 GND 0.30484f
C3940 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n9 GND 0.06065f
C3941 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.A GND 0.15634f
C3942 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0.n10 GND 0.08695f
C3943 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t0 GND 0.02265f
C3944 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t1 GND 0.13251f
C3945 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t2 GND 0.39729f
C3946 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.n0 GND 2.76756f
C3947 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t0 GND 0.02742f
C3948 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t1 GND 0.15083f
C3949 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t2 GND 0.16899f
C3950 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.n0 GND 2.83612f
C3951 a_24687_20174.t2 GND 0.16517f
C3952 a_24687_20174.t3 GND 0.06747f
C3953 a_24687_20174.n0 GND 5.15358f
C3954 a_24687_20174.t1 GND 0.07601f
C3955 a_24687_20174.n1 GND 4.60987f
C3956 a_24687_20174.t0 GND 0.12791f
C3957 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t2 GND 0.04119f
C3958 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t5 GND 0.03353f
C3959 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t8 GND 0.02094f
C3960 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n0 GND 0.06383f
C3961 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n1 GND 0.03879f
C3962 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t9 GND 0.03353f
C3963 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t7 GND 0.02094f
C3964 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n2 GND 0.06383f
C3965 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n3 GND 0.01711f
C3966 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n4 GND 0.35016f
C3967 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n5 GND 4.38855f
C3968 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n6 GND 0.18482f
C3969 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t3 GND 0.02026f
C3970 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t1 GND 0.02026f
C3971 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n7 GND 0.04503f
C3972 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t0 GND 0.07496f
C3973 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t4 GND 0.02096f
C3974 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t6 GND 0.03356f
C3975 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n8 GND 0.06289f
C3976 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n9 GND 0.05268f
C3977 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n10 GND 0.14872f
C3978 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n11 GND 0.12975f
C3979 a_33634_8950.t1 GND 0.09175f
C3980 a_33634_8950.t2 GND 0.10894f
C3981 a_33634_8950.n0 GND 5.52296f
C3982 a_33634_8950.t0 GND 0.07635f
C3983 a_27620_6250.t1 GND 0.13813f
C3984 a_27620_6250.t4 GND 0.0814f
C3985 a_27620_6250.n0 GND 5.35733f
C3986 a_27620_6250.t3 GND 0.17912f
C3987 a_27620_6250.n1 GND 4.85263f
C3988 a_27620_6250.t2 GND 0.17054f
C3989 a_27620_6250.n2 GND 5.33946f
C3990 a_27620_6250.t0 GND 0.0814f
C3991 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t0 GND 0.07325f
C3992 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n0 GND 0.03003f
C3993 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n1 GND 0.06465f
C3994 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n2 GND 0.04292f
C3995 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t1 GND 0.07018f
C3996 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t11 GND 0.14953f
C3997 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t12 GND 0.14551f
C3998 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n4 GND 0.33771f
C3999 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t8 GND 0.14321f
C4000 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n5 GND 2.12021f
C4001 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n6 GND 3.80472f
C4002 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t15 GND 0.14551f
C4003 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t9 GND 0.14482f
C4004 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n7 GND 0.45402f
C4005 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t5 GND 0.14482f
C4006 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n8 GND 0.22736f
C4007 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t17 GND 0.14482f
C4008 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n9 GND 0.18513f
C4009 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t13 GND 0.14482f
C4010 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n10 GND 0.22736f
C4011 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t19 GND 0.14482f
C4012 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n11 GND 0.22736f
C4013 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t18 GND 0.14482f
C4014 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n12 GND 0.22736f
C4015 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n13 GND 0.15135f
C4016 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t14 GND 0.14321f
C4017 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n14 GND 1.97681f
C4018 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n15 GND 5.21044f
C4019 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t4 GND 0.13854f
C4020 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t16 GND 0.13785f
C4021 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n16 GND 0.44898f
C4022 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t20 GND 0.13785f
C4023 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n17 GND 0.16315f
C4024 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t3 GND 0.13785f
C4025 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n18 GND 0.21086f
C4026 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t7 GND 0.13785f
C4027 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n19 GND 0.22484f
C4028 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t22 GND 0.13785f
C4029 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n20 GND 0.22484f
C4030 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t6 GND 0.13854f
C4031 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n21 GND 0.37549f
C4032 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t2 GND 0.13626f
C4033 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n22 GND 1.9804f
C4034 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n23 GND 7.73135f
C4035 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t21 GND 0.25618f
C4036 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.t10 GND 0.14211f
C4037 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n24 GND 0.22323f
C4038 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n25 GND 0.04441f
C4039 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3.n26 GND 0.06367f
C4040 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t0 GND 0.07426f
C4041 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t3 GND 0.04735f
C4042 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t5 GND 0.02955f
C4043 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n0 GND 0.09326f
C4044 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n1 GND 0.04267f
C4045 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t4 GND 0.04735f
C4046 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t2 GND 0.02955f
C4047 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n2 GND 0.09323f
C4048 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n3 GND 0.03149f
C4049 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n4 GND 0.48165f
C4050 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n5 GND 5.99489f
C4051 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n6 GND 0.25011f
C4052 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t1 GND 0.10587f
C4053 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n7 GND 0.02569f
C4054 a_16615_7686.t4 GND 0.0819f
C4055 a_16615_7686.t1 GND 0.07479f
C4056 a_16615_7686.n0 GND 3.75672f
C4057 a_16615_7686.t2 GND 0.09282f
C4058 a_16615_7686.t3 GND 0.07318f
C4059 a_16615_7686.n1 GND 5.4585f
C4060 a_16615_7686.n2 GND 2.6889f
C4061 a_16615_7686.t0 GND 0.07318f
C4062 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t2 GND 0.01662f
C4063 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t1 GND 0.09696f
C4064 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t0 GND 0.09405f
C4065 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.n0 GND 1.57947f
C4066 a_21375_20174.t2 GND 0.11548f
C4067 a_21375_20174.t3 GND 0.04818f
C4068 a_21375_20174.n0 GND 3.58176f
C4069 a_21375_20174.t1 GND 0.03156f
C4070 a_21375_20174.n1 GND 2.4369f
C4071 a_21375_20174.t0 GND 0.08612f
C4072 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t6 GND 0.18452f
C4073 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t3 GND 0.18452f
C4074 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n0 GND 1.4305f
C4075 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t13 GND 0.20184f
C4076 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t8 GND 0.19673f
C4077 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n1 GND 1.70817f
C4078 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t12 GND 0.20184f
C4079 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t9 GND 0.19632f
C4080 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n2 GND 1.73221f
C4081 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n3 GND 1.43567f
C4082 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t11 GND 0.20184f
C4083 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t14 GND 0.19632f
C4084 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n4 GND 1.47934f
C4085 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t15 GND 0.20184f
C4086 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t10 GND 0.19673f
C4087 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n5 GND 1.96104f
C4088 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n6 GND 1.32744f
C4089 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n7 GND 1.31284f
C4090 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t5 GND 0.18452f
C4091 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t0 GND 0.18452f
C4092 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n8 GND 1.22182f
C4093 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t2 GND 0.18452f
C4094 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t4 GND 0.18452f
C4095 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n9 GND 1.25158f
C4096 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n10 GND 2.22498f
C4097 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n11 GND 1.1146f
C4098 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n12 GND 2.27113f
C4099 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t1 GND 0.18452f
C4100 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n13 GND 1.05912f
C4101 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t7 GND 0.18452f
C4102 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.t2 GND 0.07822f
C4103 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.t1 GND 0.08851f
C4104 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.n0 GND 1.81943f
C4105 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11.t0 GND 0.01384f
C4106 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.t2 GND 0.10511f
C4107 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.t1 GND 0.10221f
C4108 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.n0 GND 2.37213f
C4109 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12.t0 GND 0.02055f
C4110 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t0 GND 0.09866f
C4111 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n0 GND 0.04045f
C4112 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n1 GND 0.08708f
C4113 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n2 GND 0.05782f
C4114 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t1 GND 0.09452f
C4115 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n3 GND 0.01194f
C4116 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t2 GND 0.19507f
C4117 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n4 GND 0.25416f
C4118 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t5 GND 0.19507f
C4119 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n5 GND 0.30624f
C4120 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t4 GND 0.196f
C4121 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t6 GND 0.19507f
C4122 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n6 GND 0.61154f
C4123 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n7 GND 0.20386f
C4124 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].t3 GND 0.1929f
C4125 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n8 GND 13.9648f
C4126 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5].n9 GND 0.06224f
C4127 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t3 GND 0.01968f
C4128 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t1 GND 0.01968f
C4129 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n0 GND 0.04693f
C4130 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n1 GND 0.09219f
C4131 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t12 GND 0.0471f
C4132 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t9 GND 0.02775f
C4133 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t11 GND 0.0471f
C4134 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t8 GND 0.02775f
C4135 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n2 GND 0.07902f
C4136 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n3 GND 0.11723f
C4137 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n4 GND 0.03535f
C4138 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t6 GND 0.03129f
C4139 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t5 GND 0.05012f
C4140 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n5 GND 0.09554f
C4141 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n6 GND 0.15506f
C4142 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n7 GND 0.75373f
C4143 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t10 GND 0.03124f
C4144 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t7 GND 0.05005f
C4145 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n8 GND 0.09952f
C4146 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t4 GND 0.03129f
C4147 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t13 GND 0.05012f
C4148 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n9 GND 0.0954f
C4149 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n10 GND 0.01346f
C4150 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n11 GND 0.34761f
C4151 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n12 GND 8.72639f
C4152 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n13 GND 6.93802f
C4153 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n14 GND 0.02166f
C4154 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n15 GND 0.02868f
C4155 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t0 GND 0.03028f
C4156 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t2 GND 0.03028f
C4157 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n16 GND 0.06649f
C4158 a_31594_7686.t1 GND 0.11133f
C4159 a_31594_7686.t2 GND 0.08541f
C4160 a_31594_7686.n0 GND 3.94271f
C4161 a_31594_7686.t4 GND 0.08147f
C4162 a_31594_7686.n1 GND 2.66272f
C4163 a_31594_7686.t3 GND 0.14987f
C4164 a_31594_7686.n2 GND 5.98504f
C4165 a_31594_7686.t0 GND 0.08147f
C4166 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t2 GND 0.02716f
C4167 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t1 GND 0.16449f
C4168 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t0 GND 0.1492f
C4169 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.n0 GND 2.95161f
C4170 a_15629_7686.t4 GND 0.07971f
C4171 a_15629_7686.t2 GND 0.0947f
C4172 a_15629_7686.t1 GND 0.07612f
C4173 a_15629_7686.n0 GND 5.33217f
C4174 a_15629_7686.t3 GND 0.07612f
C4175 a_15629_7686.n1 GND 2.97065f
C4176 a_15629_7686.n2 GND 3.98477f
C4177 a_15629_7686.t0 GND 0.08576f
C4178 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t0 GND 0.08409f
C4179 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n0 GND 0.03448f
C4180 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n1 GND 0.07422f
C4181 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n2 GND 0.04927f
C4182 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t1 GND 0.08056f
C4183 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n3 GND 0.01018f
C4184 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t6 GND 0.16704f
C4185 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t8 GND 0.16625f
C4186 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n4 GND 0.52118f
C4187 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t9 GND 0.16625f
C4188 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n5 GND 0.26099f
C4189 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t3 GND 0.16625f
C4190 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n6 GND 0.26099f
C4191 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t13 GND 0.16625f
C4192 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n7 GND 0.26099f
C4193 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t17 GND 0.16625f
C4194 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n8 GND 0.26099f
C4195 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t2 GND 0.16625f
C4196 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n9 GND 0.26099f
C4197 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t4 GND 0.16625f
C4198 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n10 GND 0.2138f
C4199 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t12 GND 0.16704f
C4200 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t7 GND 0.16625f
C4201 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n11 GND 0.52118f
C4202 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t5 GND 0.16625f
C4203 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n12 GND 0.26099f
C4204 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t11 GND 0.16625f
C4205 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n13 GND 0.21681f
C4206 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t14 GND 0.16704f
C4207 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t10 GND 0.16625f
C4208 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n14 GND 0.52118f
C4209 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t16 GND 0.16625f
C4210 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n15 GND 0.26099f
C4211 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.t15 GND 0.16625f
C4212 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n16 GND 0.21681f
C4213 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n17 GND 0.2093f
C4214 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n18 GND 16.7136f
C4215 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3.n19 GND 0.07943f
C4216 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t1 GND 0.01441f
C4217 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t2 GND 0.08695f
C4218 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t0 GND 0.07745f
C4219 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.n0 GND 1.43576f
C4220 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t2 GND 0.04142f
C4221 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t3 GND 0.04142f
C4222 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 GND 0.09096f
C4223 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y GND 0.20814f
C4224 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 GND 0.03924f
C4225 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t6 GND 0.06443f
C4226 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t8 GND 0.03797f
C4227 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t5 GND 0.06443f
C4228 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t7 GND 0.03797f
C4229 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 GND 0.1081f
C4230 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 GND 0.16037f
C4231 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.A GND 0.01074f
C4232 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 GND 0.04836f
C4233 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t4 GND 0.55071f
C4234 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 GND 15.822f
C4235 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 GND 0.02963f
C4236 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t1 GND 0.02692f
C4237 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t0 GND 0.02692f
C4238 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 GND 0.06419f
C4239 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 GND 0.12611f
C4240 a_15224_18696.t2 GND 0.03715f
C4241 a_15224_18696.t1 GND 0.02918f
C4242 a_15224_18696.n0 GND 2.00335f
C4243 a_15224_18696.t0 GND 0.03032f
C4244 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.t1 GND 0.11479f
C4245 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.t2 GND 0.11222f
C4246 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.n0 GND 2.55165f
C4247 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6.t0 GND 0.02134f
C4248 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t0 GND 0.0937f
C4249 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n0 GND 0.03842f
C4250 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n1 GND 0.0827f
C4251 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n2 GND 0.05491f
C4252 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t1 GND 0.08977f
C4253 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n3 GND 0.01134f
C4254 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t8 GND 0.18615f
C4255 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t3 GND 0.18526f
C4256 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n4 GND 0.58079f
C4257 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t2 GND 0.18526f
C4258 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n5 GND 0.29084f
C4259 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t9 GND 0.18526f
C4260 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n6 GND 0.29084f
C4261 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t4 GND 0.18526f
C4262 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n7 GND 0.29084f
C4263 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t7 GND 0.18526f
C4264 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n8 GND 0.29084f
C4265 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t11 GND 0.18526f
C4266 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n9 GND 0.29084f
C4267 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t5 GND 0.18526f
C4268 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n10 GND 0.29022f
C4269 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t10 GND 0.18526f
C4270 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n11 GND 0.19865f
C4271 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n12 GND 16.0287f
C4272 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t12 GND 0.3277f
C4273 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].t6 GND 0.18179f
C4274 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n13 GND 0.28556f
C4275 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n14 GND 0.05681f
C4276 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6].n15 GND 0.08145f
C4277 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t2 GND 0.03385f
C4278 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t1 GND 0.03293f
C4279 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n0 GND 0.67533f
C4280 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t3 GND 0.03385f
C4281 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t0 GND 0.03293f
C4282 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n1 GND 0.52074f
C4283 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n2 GND 0.64975f
C4284 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t5 GND 0.02952f
C4285 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t6 GND 0.02948f
C4286 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n3 GND 0.2736f
C4287 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t4 GND 0.02952f
C4288 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t7 GND 0.02948f
C4289 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n4 GND 0.29926f
C4290 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n5 GND 0.58174f
C4291 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t1 GND 0.03811f
C4292 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t2 GND 0.03811f
C4293 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 GND 0.08371f
C4294 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y GND 0.19154f
C4295 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 GND 0.03611f
C4296 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t4 GND 0.05929f
C4297 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t8 GND 0.03494f
C4298 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t10 GND 0.05929f
C4299 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t5 GND 0.03494f
C4300 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 GND 0.09948f
C4301 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 GND 0.14758f
C4302 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 GND 0.04451f
C4303 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t6 GND 0.06301f
C4304 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t11 GND 0.03932f
C4305 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 GND 0.12528f
C4306 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.A GND 0.02173f
C4307 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t12 GND 0.06309f
C4308 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t9 GND 0.03939f
C4309 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 GND 0.1201f
C4310 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 GND 0.03507f
C4311 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.B GND 0.1019f
C4312 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[1] GND 2.24751f
C4313 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t7 GND 0.23705f
C4314 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 GND 9.91961f
C4315 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 GND 3.7575f
C4316 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 GND 0.02727f
C4317 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t3 GND 0.02477f
C4318 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t0 GND 0.02477f
C4319 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 GND 0.05907f
C4320 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 GND 0.11606f
C4321 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t2 GND 0.35314f
C4322 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t5 GND 0.33746f
C4323 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n0 GND 1.70865f
C4324 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t1 GND 0.16146f
C4325 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t0 GND 0.10648f
C4326 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n1 GND 0.80542f
C4327 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t4 GND 0.16156f
C4328 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n2 GND 1.08214f
C4329 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t3 GND 0.15721f
C4330 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n3 GND 0.91022f
C4331 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t6 GND 0.29044f
C4332 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t7 GND 0.2897f
C4333 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n4 GND 0.31239f
C4334 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t8 GND 0.29044f
C4335 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.t9 GND 0.2897f
C4336 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n5 GND 0.31239f
C4337 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n6 GND 0.20457f
C4338 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B.n7 GND 0.55947f
C4339 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t27 GND 0.03427f
C4340 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t24 GND 0.03427f
C4341 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n0 GND 0.07176f
C4342 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t26 GND 0.13193f
C4343 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n1 GND 0.64193f
C4344 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t25 GND 0.12877f
C4345 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t3 GND 0.12877f
C4346 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t1 GND 0.12877f
C4347 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t21 GND 0.12877f
C4348 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t7 GND 0.03427f
C4349 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t19 GND 0.03427f
C4350 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n2 GND 0.07176f
C4351 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t20 GND 0.12877f
C4352 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t14 GND 0.12877f
C4353 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t11 GND 0.03427f
C4354 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t13 GND 0.03427f
C4355 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n3 GND 0.07176f
C4356 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t12 GND 0.12877f
C4357 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t17 GND 0.12877f
C4358 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t15 GND 0.03427f
C4359 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t18 GND 0.03427f
C4360 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n4 GND 0.07176f
C4361 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t16 GND 0.12877f
C4362 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t37 GND 0.85385f
C4363 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t43 GND 0.63023f
C4364 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n5 GND 0.75417f
C4365 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t36 GND 0.85385f
C4366 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t29 GND 0.63023f
C4367 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n6 GND 0.75417f
C4368 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n7 GND 0.15618f
C4369 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t40 GND 0.85385f
C4370 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t45 GND 0.63023f
C4371 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n8 GND 0.75417f
C4372 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t38 GND 0.85385f
C4373 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t32 GND 0.63023f
C4374 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n9 GND 0.75417f
C4375 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n10 GND 0.12956f
C4376 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n11 GND 0.56592f
C4377 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t33 GND 0.85385f
C4378 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t39 GND 0.63023f
C4379 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n12 GND 0.75417f
C4380 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t31 GND 0.85385f
C4381 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t44 GND 0.63023f
C4382 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n13 GND 0.75417f
C4383 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n14 GND 0.12956f
C4384 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n15 GND 0.38268f
C4385 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t30 GND 0.85385f
C4386 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t35 GND 0.63023f
C4387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n16 GND 0.75417f
C4388 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t28 GND 0.85385f
C4389 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t42 GND 0.63023f
C4390 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n17 GND 0.75417f
C4391 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n18 GND 0.12956f
C4392 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n19 GND 0.38268f
C4393 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t47 GND 0.85385f
C4394 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t34 GND 0.63023f
C4395 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n20 GND 0.75417f
C4396 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t46 GND 0.85385f
C4397 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t41 GND 0.63023f
C4398 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n21 GND 0.75417f
C4399 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n22 GND 0.12956f
C4400 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n23 GND 3.60018f
C4401 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t8 GND 0.08229f
C4402 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t6 GND 0.01828f
C4403 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t5 GND 0.01828f
C4404 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n24 GND 0.03957f
C4405 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t10 GND 0.01828f
C4406 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t4 GND 0.01828f
C4407 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n25 GND 0.03957f
C4408 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t22 GND 0.01828f
C4409 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t23 GND 0.01828f
C4410 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n26 GND 0.07447f
C4411 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n27 GND 0.44489f
C4412 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n28 GND 0.41803f
C4413 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t9 GND 0.0784f
C4414 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n29 GND 0.64686f
C4415 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n30 GND 0.40201f
C4416 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n31 GND 2.25602f
C4417 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n32 GND 0.66179f
C4418 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n33 GND 0.36474f
C4419 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n34 GND 0.3912f
C4420 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n35 GND 0.31649f
C4421 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n36 GND 0.36474f
C4422 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n37 GND 0.3912f
C4423 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n38 GND 0.31649f
C4424 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n39 GND 0.36474f
C4425 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n40 GND 0.3912f
C4426 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n41 GND 0.31649f
C4427 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t0 GND 0.03427f
C4428 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t2 GND 0.03427f
C4429 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n42 GND 0.07176f
C4430 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n43 GND 0.36474f
C4431 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n44 GND 0.39119f
C4432 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n45 GND 0.31649f
C4433 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t0 GND 0.09613f
C4434 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n0 GND 0.03941f
C4435 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n1 GND 0.08484f
C4436 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n2 GND 0.05633f
C4437 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t1 GND 0.09209f
C4438 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n3 GND 0.01163f
C4439 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t5 GND 0.18415f
C4440 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t4 GND 0.19024f
C4441 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n4 GND 0.74208f
C4442 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t6 GND 0.19005f
C4443 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n5 GND 0.39697f
C4444 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t9 GND 0.18793f
C4445 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n6 GND 1.94518f
C4446 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n7 GND 8.90143f
C4447 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t2 GND 0.18151f
C4448 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t8 GND 0.17881f
C4449 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n8 GND 1.92539f
C4450 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n9 GND 11.3951f
C4451 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t3 GND 0.33618f
C4452 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.t7 GND 0.18649f
C4453 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n10 GND 0.29294f
C4454 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n11 GND 0.05828f
C4455 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1.n12 GND 0.08356f
C4456 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t6 GND 0.23142f
C4457 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t13 GND 0.24661f
C4458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t1 GND 0.23142f
C4459 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t5 GND 0.23142f
C4460 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n0 GND 1.02719f
C4461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n1 GND 1.33348f
C4462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t2 GND 0.23136f
C4463 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t12 GND 0.23136f
C4464 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n2 GND 0.73738f
C4465 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n3 GND 1.24044f
C4466 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t16 GND 0.26105f
C4467 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t18 GND 0.2503f
C4468 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n4 GND 1.89151f
C4469 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t24 GND 0.2503f
C4470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n5 GND 1.59785f
C4471 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t22 GND 0.23352f
C4472 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t20 GND 0.2335f
C4473 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n6 GND 1.21388f
C4474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t17 GND 0.2503f
C4475 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n7 GND 1.2622f
C4476 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t31 GND 0.2503f
C4477 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n8 GND 1.05359f
C4478 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t29 GND 0.2503f
C4479 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n9 GND 1.01045f
C4480 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n10 GND 1.13336f
C4481 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t30 GND 0.2335f
C4482 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t27 GND 0.23352f
C4483 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n11 GND 1.21388f
C4484 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t25 GND 0.2503f
C4485 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n12 GND 1.2622f
C4486 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t23 GND 0.2503f
C4487 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n13 GND 1.05359f
C4488 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t26 GND 0.2503f
C4489 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n14 GND 1.32752f
C4490 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t21 GND 0.26105f
C4491 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t28 GND 0.2503f
C4492 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n15 GND 1.89151f
C4493 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t19 GND 0.2503f
C4494 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n16 GND 1.28078f
C4495 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n17 GND 1.12088f
C4496 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n18 GND 1.17777f
C4497 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t7 GND 0.2583f
C4498 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t9 GND 0.23142f
C4499 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t0 GND 0.23142f
C4500 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n19 GND 1.02719f
C4501 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n20 GND 2.29133f
C4502 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t4 GND 0.24661f
C4503 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t8 GND 0.23142f
C4504 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t3 GND 0.23142f
C4505 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n21 GND 1.02719f
C4506 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n22 GND 1.33348f
C4507 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t11 GND 0.23136f
C4508 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t14 GND 0.23136f
C4509 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n23 GND 0.73738f
C4510 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n24 GND 0.92337f
C4511 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n25 GND 1.35167f
C4512 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n26 GND 1.52381f
C4513 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n27 GND 1.40802f
C4514 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t10 GND 0.2583f
C4515 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n28 GND 1.97426f
C4516 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n29 GND 1.02719f
C4517 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t15 GND 0.23142f
C4518 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t10 GND 0.13816f
C4519 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n0 GND 0.17342f
C4520 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t19 GND 0.13816f
C4521 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n1 GND 0.22536f
C4522 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t8 GND 0.13816f
C4523 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n2 GND 0.22536f
C4524 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t21 GND 0.13816f
C4525 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n3 GND 0.22536f
C4526 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t14 GND 0.13816f
C4527 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n4 GND 0.22536f
C4528 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t15 GND 0.13887f
C4529 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t4 GND 0.13816f
C4530 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n5 GND 0.45002f
C4531 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t12 GND 0.13816f
C4532 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n6 GND 0.22536f
C4533 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t3 GND 0.13816f
C4534 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n7 GND 0.22536f
C4535 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t5 GND 0.13816f
C4536 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n8 GND 0.22536f
C4537 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t17 GND 0.13816f
C4538 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n9 GND 0.22536f
C4539 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t7 GND 0.13816f
C4540 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n10 GND 0.22536f
C4541 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t11 GND 0.13816f
C4542 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n11 GND 0.22536f
C4543 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t18 GND 0.13816f
C4544 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n12 GND 0.22536f
C4545 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t9 GND 0.13816f
C4546 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n13 GND 0.22536f
C4547 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t16 GND 0.13816f
C4548 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n14 GND 0.22536f
C4549 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n15 GND 0.1517f
C4550 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t6 GND 0.13657f
C4551 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n16 GND 15.1085f
C4552 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t0 GND 0.11443f
C4553 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t1 GND 0.09714f
C4554 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n17 GND 0.94738f
C4555 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t20 GND 0.45357f
C4556 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t13 GND 0.4517f
C4557 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n18 GND 0.74878f
C4558 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].t2 GND 0.4517f
C4559 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n19 GND 0.38634f
C4560 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0].n20 GND 0.7067f
C4561 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t0 GND 0.05778f
C4562 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t1 GND 0.05865f
C4563 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n0 GND 1.04124f
C4564 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t3 GND 0.05535f
C4565 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t2 GND 0.054f
C4566 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n1 GND 0.78821f
C4567 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t2 GND 0.04008f
C4568 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t3 GND 0.04008f
C4569 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n0 GND 0.08803f
C4570 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n1 GND 0.03797f
C4571 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t10 GND 0.06645f
C4572 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t16 GND 0.04151f
C4573 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n2 GND 0.12322f
C4574 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t11 GND 0.06618f
C4575 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t4 GND 0.04129f
C4576 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n3 GND 0.13445f
C4577 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n4 GND 0.15582f
C4578 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t8 GND 0.04136f
C4579 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t6 GND 0.06626f
C4580 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n5 GND 0.13065f
C4581 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n6 GND 0.08905f
C4582 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n7 GND 0.49955f
C4583 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n8 GND 0.84298f
C4584 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t17 GND 0.04136f
C4585 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t13 GND 0.06626f
C4586 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n9 GND 0.13038f
C4587 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n10 GND 0.08233f
C4588 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n11 GND 0.58676f
C4589 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t7 GND 0.06626f
C4590 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t12 GND 0.04136f
C4591 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n12 GND 0.13038f
C4592 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n13 GND 0.05851f
C4593 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t9 GND 0.06626f
C4594 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t15 GND 0.04136f
C4595 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n14 GND 0.13175f
C4596 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t14 GND 0.06635f
C4597 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t5 GND 0.04143f
C4598 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n15 GND 0.1263f
C4599 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n16 GND 0.0229f
C4600 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n17 GND 0.03311f
C4601 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n18 GND 0.46233f
C4602 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n19 GND 11.365f
C4603 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n20 GND 7.93634f
C4604 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t0 GND 0.02605f
C4605 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t1 GND 0.02605f
C4606 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n21 GND 0.06212f
C4607 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n22 GND 0.12205f
C4608 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.t1 GND 0.09383f
C4609 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.t2 GND 0.01431f
C4610 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.n0 GND 1.89096f
C4611 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21.t0 GND 0.1009f
C4612 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.t1 GND 0.09527f
C4613 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.t2 GND 0.0165f
C4614 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.n0 GND 2.09304f
C4615 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22.t0 GND 0.0952f
C4616 a_24135_20174.t2 GND 0.15093f
C4617 a_24135_20174.t1 GND 0.17697f
C4618 a_24135_20174.t3 GND 0.07252f
C4619 a_24135_20174.n0 GND 5.33538f
C4620 a_24135_20174.n1 GND 5.6647f
C4621 a_24135_20174.t0 GND 0.0995f
C4622 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t1 GND 0.0257f
C4623 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t2 GND 0.0257f
C4624 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 GND 0.06128f
C4625 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y GND 0.19868f
C4626 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 GND 0.12038f
C4627 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t8 GND 0.06536f
C4628 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t5 GND 0.04079f
C4629 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 GND 0.12995f
C4630 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.B GND 0.05637f
C4631 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.A GND 0.02254f
C4632 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t6 GND 0.06545f
C4633 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t4 GND 0.04086f
C4634 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 GND 0.12458f
C4635 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 GND 0.02451f
C4636 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 GND 0.06185f
C4637 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[1] GND 2.34134f
C4638 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t7 GND 0.24665f
C4639 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 GND 11.5282f
C4640 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 GND 2.61648f
C4641 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 GND 0.03746f
C4642 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t3 GND 0.03954f
C4643 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t0 GND 0.03954f
C4644 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 GND 0.08683f
C4645 a_18724_8950.t2 GND 0.03722f
C4646 a_18724_8950.t1 GND 0.0341f
C4647 a_18724_8950.n0 GND 2.59201f
C4648 a_18724_8950.t0 GND 0.03667f
C4649 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t0 GND 0.09004f
C4650 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n0 GND 0.03692f
C4651 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n1 GND 0.07947f
C4652 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n2 GND 0.05276f
C4653 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t1 GND 0.08626f
C4654 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n3 GND 0.0109f
C4655 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t11 GND 0.17679f
C4656 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t7 GND 0.17887f
C4657 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n4 GND 0.85354f
C4658 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t4 GND 0.17802f
C4659 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n5 GND 0.21173f
C4660 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t10 GND 0.17802f
C4661 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n6 GND 0.27947f
C4662 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t2 GND 0.17887f
C4663 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n7 GND 0.46467f
C4664 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t8 GND 0.17604f
C4665 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n8 GND 1.92907f
C4666 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n9 GND 9.26347f
C4667 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t6 GND 0.1703f
C4668 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t3 GND 0.16944f
C4669 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n10 GND 0.49865f
C4670 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t5 GND 0.1703f
C4671 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n11 GND 0.4218f
C4672 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.t9 GND 0.16749f
C4673 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n12 GND 1.91752f
C4674 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n13 GND 9.84727f
C4675 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2.n14 GND 0.0568f
C4676 top_DAC_0/top_final_switch_0.VOUT[3].t3 GND 0.01004f
C4677 top_DAC_0/top_final_switch_0.VOUT[3].t2 GND 0.01004f
C4678 top_DAC_0/top_final_switch_0.VOUT[3].n0 GND 0.02286f
C4679 top_DAC_0/top_final_switch_0.VOUT[3].t0 GND 0.01004f
C4680 top_DAC_0/top_final_switch_0.VOUT[3].t1 GND 0.01004f
C4681 top_DAC_0/top_final_switch_0.VOUT[3].n1 GND 0.02386f
C4682 top_DAC_0/top_final_switch_0.VOUT[3].n2 GND 1.36118f
C4683 top_DAC_0/top_final_switch_0.VOUT[3].t9 GND 0.93418f
C4684 top_DAC_0/top_final_switch_0.VOUT[3].t5 GND 0.92835f
C4685 top_DAC_0/top_final_switch_0.VOUT[3].n3 GND 1.549f
C4686 top_DAC_0/top_final_switch_0.VOUT[3].t8 GND 0.92897f
C4687 top_DAC_0/top_final_switch_0.VOUT[3].t11 GND 0.92728f
C4688 top_DAC_0/top_final_switch_0.VOUT[3].n4 GND 1.19609f
C4689 top_DAC_0/top_final_switch_0.VOUT[3].n5 GND 0.80264f
C4690 top_DAC_0/top_final_switch_0.VOUT[3].t6 GND 0.38166f
C4691 top_DAC_0/top_final_switch_0.VOUT[3].t10 GND 0.37983f
C4692 top_DAC_0/top_final_switch_0.VOUT[3].n6 GND 1.00874f
C4693 top_DAC_0/top_final_switch_0.VOUT[3].t7 GND 0.38796f
C4694 top_DAC_0/top_final_switch_0.VOUT[3].t4 GND 0.3814f
C4695 top_DAC_0/top_final_switch_0.VOUT[3].n7 GND 1.1236f
C4696 top_DAC_0/top_final_switch_0.VOUT[3].n8 GND 0.56741f
C4697 top_DAC_0/top_final_switch_0.VOUT[3].n9 GND 1.52514f
C4698 top_DAC_0/top_final_switch_0.VOUT[3].n10 GND 0.27046f
C4699 top_DAC_0/top_rseg_n_dcell_0.SH[2].t1 GND 0.11219f
C4700 top_DAC_0/top_rseg_n_dcell_0.SH[2].n0 GND 0.046f
C4701 top_DAC_0/top_rseg_n_dcell_0.SH[2].n1 GND 0.09903f
C4702 top_DAC_0/top_rseg_n_dcell_0.SH[2].n2 GND 0.06574f
C4703 top_DAC_0/top_rseg_n_dcell_0.SH[2].t4 GND 0.20956f
C4704 top_DAC_0/top_rseg_n_dcell_0.SH[2].t2 GND 0.2087f
C4705 top_DAC_0/top_rseg_n_dcell_0.SH[2].n3 GND 0.41388f
C4706 top_DAC_0/top_rseg_n_dcell_0.SH[2].t5 GND 0.2087f
C4707 top_DAC_0/top_rseg_n_dcell_0.SH[2].n4 GND 0.23032f
C4708 top_DAC_0/top_rseg_n_dcell_0.SH[2].t3 GND 0.2087f
C4709 top_DAC_0/top_rseg_n_dcell_0.SH[2].n5 GND 0.23032f
C4710 top_DAC_0/top_rseg_n_dcell_0.SH[2].t6 GND 0.2087f
C4711 top_DAC_0/top_rseg_n_dcell_0.SH[2].n6 GND 0.24637f
C4712 top_DAC_0/top_rseg_n_dcell_0.SH[2].n7 GND 0.07614f
C4713 top_DAC_0/top_rseg_n_dcell_0.SH[2].t0 GND 0.10749f
C4714 top_DAC_0/top_rseg_n_dcell_0.SH[2].n8 GND 0.0556f
C4715 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n0 GND 0.01746f
C4716 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n1 GND 0.09034f
C4717 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n2 GND 0.0829f
C4718 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n3 GND 0.08269f
C4719 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t56 GND 0.15492f
C4720 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t42 GND 0.15358f
C4721 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n4 GND 0.38143f
C4722 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t28 GND 0.15358f
C4723 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n5 GND 0.19139f
C4724 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t8 GND 0.15358f
C4725 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n6 GND 0.19139f
C4726 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t61 GND 0.15358f
C4727 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n7 GND 0.19139f
C4728 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t20 GND 0.15358f
C4729 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n8 GND 0.19139f
C4730 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t22 GND 0.15358f
C4731 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n9 GND 0.19139f
C4732 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t45 GND 0.15358f
C4733 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n10 GND 0.19139f
C4734 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t23 GND 0.15358f
C4735 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n11 GND 0.19139f
C4736 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t14 GND 0.15358f
C4737 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n12 GND 0.19139f
C4738 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t65 GND 0.15358f
C4739 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n13 GND 0.1661f
C4740 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t27 GND 0.15492f
C4741 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t35 GND 0.15358f
C4742 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n14 GND 0.38143f
C4743 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t54 GND 0.15358f
C4744 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n15 GND 0.19139f
C4745 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t12 GND 0.15358f
C4746 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n16 GND 0.19139f
C4747 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t41 GND 0.15358f
C4748 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n17 GND 0.16326f
C4749 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n18 GND 0.06574f
C4750 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t59 GND 0.15567f
C4751 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t44 GND 0.15358f
C4752 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n19 GND 0.4875f
C4753 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t21 GND 0.15358f
C4754 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n20 GND 0.19139f
C4755 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t10 GND 0.15358f
C4756 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n21 GND 0.19139f
C4757 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t38 GND 0.15358f
C4758 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n22 GND 0.19139f
C4759 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t39 GND 0.15358f
C4760 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n23 GND 0.19139f
C4761 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t64 GND 0.15358f
C4762 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n24 GND 0.19139f
C4763 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t40 GND 0.15358f
C4764 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n25 GND 0.19139f
C4765 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t26 GND 0.15358f
C4766 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n26 GND 0.19139f
C4767 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t15 GND 0.15358f
C4768 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n27 GND 0.1661f
C4769 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t52 GND 0.31403f
C4770 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t7 GND 0.31286f
C4771 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n28 GND 0.49793f
C4772 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t47 GND 0.31403f
C4773 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t4 GND 0.31286f
C4774 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n29 GND 0.5037f
C4775 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n30 GND 0.53799f
C4776 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t49 GND 0.15358f
C4777 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n31 GND 0.94496f
C4778 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t6 GND 0.15358f
C4779 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n32 GND 0.19139f
C4780 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t25 GND 0.15358f
C4781 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n33 GND 0.19139f
C4782 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t55 GND 0.15358f
C4783 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n34 GND 0.16326f
C4784 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n35 GND 0.05341f
C4785 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n36 GND 0.33285f
C4786 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t16 GND 0.15567f
C4787 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t67 GND 0.15358f
C4788 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n37 GND 0.4875f
C4789 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t43 GND 0.15358f
C4790 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n38 GND 0.19139f
C4791 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t30 GND 0.15358f
C4792 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n39 GND 0.19139f
C4793 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t58 GND 0.15358f
C4794 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n40 GND 0.19139f
C4795 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t60 GND 0.15358f
C4796 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n41 GND 0.19139f
C4797 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t17 GND 0.15358f
C4798 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n42 GND 0.19139f
C4799 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t63 GND 0.15358f
C4800 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n43 GND 0.19139f
C4801 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t48 GND 0.15358f
C4802 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n44 GND 0.19139f
C4803 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t32 GND 0.15358f
C4804 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n45 GND 0.1661f
C4805 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t5 GND 0.15567f
C4806 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t24 GND 0.15358f
C4807 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n46 GND 0.4875f
C4808 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t46 GND 0.15358f
C4809 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n47 GND 0.19139f
C4810 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t13 GND 0.15358f
C4811 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n48 GND 0.16326f
C4812 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n49 GND 0.05341f
C4813 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n50 GND 0.23704f
C4814 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t36 GND 0.15492f
C4815 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t37 GND 0.15358f
C4816 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n51 GND 0.38143f
C4817 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t62 GND 0.15358f
C4818 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n52 GND 0.19139f
C4819 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t18 GND 0.15358f
C4820 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n53 GND 0.19139f
C4821 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t19 GND 0.15358f
C4822 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n54 GND 0.19139f
C4823 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t57 GND 0.15358f
C4824 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n55 GND 0.19139f
C4825 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t66 GND 0.15358f
C4826 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n56 GND 0.19139f
C4827 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t29 GND 0.15358f
C4828 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n57 GND 0.19139f
C4829 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t51 GND 0.15358f
C4830 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n58 GND 0.19139f
C4831 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t53 GND 0.15358f
C4832 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n59 GND 0.19139f
C4833 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t11 GND 0.15358f
C4834 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n60 GND 0.1661f
C4835 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t33 GND 0.15492f
C4836 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t31 GND 0.15358f
C4837 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n61 GND 0.38143f
C4838 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t9 GND 0.15358f
C4839 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n62 GND 0.19139f
C4840 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t50 GND 0.15358f
C4841 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n63 GND 0.19139f
C4842 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t34 GND 0.15358f
C4843 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n64 GND 0.16326f
C4844 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n65 GND 0.05341f
C4845 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n66 GND 0.5305f
C4846 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n67 GND 0.01746f
C4847 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n68 GND 0.19226f
C4848 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n69 GND 0.08269f
C4849 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n70 GND 0.07458f
C4850 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n71 GND 0.53524f
C4851 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n72 GND 0.07796f
C4852 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n73 GND 0.08192f
C4853 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t24 GND 2.8674f
C4854 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t22 GND 1.93769f
C4855 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n0 GND 1.77419f
C4856 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t23 GND 0.02043f
C4857 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t21 GND 0.09009f
C4858 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t13 GND 0.06067f
C4859 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t5 GND 0.06067f
C4860 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n1 GND 0.31327f
C4861 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t4 GND 0.06067f
C4862 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t8 GND 0.06067f
C4863 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n2 GND 0.2523f
C4864 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n3 GND 0.37106f
C4865 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t6 GND 0.06067f
C4866 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t12 GND 0.06067f
C4867 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n4 GND 0.2523f
C4868 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n5 GND 0.2835f
C4869 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t7 GND 0.06067f
C4870 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t14 GND 0.06067f
C4871 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n6 GND 0.2523f
C4872 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n7 GND 0.2835f
C4873 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t15 GND 0.06067f
C4874 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t0 GND 0.06067f
C4875 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n8 GND 0.23066f
C4876 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n9 GND 0.38691f
C4877 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t16 GND 0.06067f
C4878 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t1 GND 0.06067f
C4879 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n10 GND 0.29163f
C4880 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t3 GND 0.06067f
C4881 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t2 GND 0.06067f
C4882 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n11 GND 0.2523f
C4883 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n12 GND 0.37106f
C4884 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t10 GND 0.06067f
C4885 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t9 GND 0.06067f
C4886 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n13 GND 0.2523f
C4887 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n14 GND 0.2835f
C4888 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t11 GND 0.06067f
C4889 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t19 GND 0.06067f
C4890 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n15 GND 0.2523f
C4891 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n16 GND 0.2835f
C4892 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t18 GND 0.06067f
C4893 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t17 GND 0.06067f
C4894 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n17 GND 0.2523f
C4895 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n18 GND 0.39811f
C4896 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n19 GND 4.90173f
C4897 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n20 GND 2.44538f
C4898 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n21 GND 0.2183f
C4899 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n22 GND 0.28717f
C4900 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t20 GND 2.8674f
C4901 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t25 GND 1.93769f
C4902 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n23 GND 1.76738f
C4903 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n24 GND 0.20492f
C4904 top_DAC_0/top_rseg_n_dcell_0.VL2.t4 GND 0.02346f
C4905 top_DAC_0/top_rseg_n_dcell_0.VL2.t6 GND 0.02766f
C4906 top_DAC_0/top_rseg_n_dcell_0.VL2.t1 GND 0.02638f
C4907 top_DAC_0/top_rseg_n_dcell_0.VL2.n0 GND 0.58962f
C4908 top_DAC_0/top_rseg_n_dcell_0.VL2.t8 GND 0.02638f
C4909 top_DAC_0/top_rseg_n_dcell_0.VL2.n1 GND 0.31558f
C4910 top_DAC_0/top_rseg_n_dcell_0.VL2.n2 GND 0.02488f
C4911 top_DAC_0/top_rseg_n_dcell_0.VL2.n3 GND 1.80854f
C4912 top_DAC_0/top_rseg_n_dcell_0.VL2.t5 GND 0.02427f
C4913 top_DAC_0/top_rseg_n_dcell_0.VL2.t7 GND 0.02314f
C4914 top_DAC_0/top_rseg_n_dcell_0.VL2.n4 GND 0.21836f
C4915 top_DAC_0/top_rseg_n_dcell_0.VL2.t3 GND 0.02314f
C4916 top_DAC_0/top_rseg_n_dcell_0.VL2.n5 GND 0.08405f
C4917 top_DAC_0/top_rseg_n_dcell_0.VL2.t2 GND 0.02314f
C4918 top_DAC_0/top_rseg_n_dcell_0.VL2.n6 GND 0.08405f
C4919 top_DAC_0/top_rseg_n_dcell_0.VL2.t0 GND 0.02314f
C4920 top_DAC_0/top_rseg_n_dcell_0.VL2.n7 GND 0.12636f
C4921 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t3 GND 0.24388f
C4922 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t2 GND 0.22393f
C4923 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n0 GND 3.24351f
C4924 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t0 GND 0.21007f
C4925 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n1 GND 1.67961f
C4926 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t1 GND 0.199f
C4927 top_DAC_0/top_rseg_n_dcell_0.VL3.t0 GND 0.01953f
C4928 top_DAC_0/top_rseg_n_dcell_0.VL3.t4 GND 0.02028f
C4929 top_DAC_0/top_rseg_n_dcell_0.VL3.n1 GND 1.11042f
C4930 top_DAC_0/top_rseg_n_dcell_0.VL3.t2 GND 0.01955f
C4931 top_DAC_0/top_rseg_n_dcell_0.VL3.t3 GND 0.01949f
C4932 top_DAC_0/top_rseg_n_dcell_0.VL3.n2 GND 0.10283f
C4933 top_DAC_0/top_rseg_n_dcell_0.VL3.t5 GND 0.01949f
C4934 top_DAC_0/top_rseg_n_dcell_0.VL3.n3 GND 0.07066f
C4935 top_DAC_0/top_rseg_n_dcell_0.VL3.t6 GND 0.01949f
C4936 top_DAC_0/top_rseg_n_dcell_0.VL3.n4 GND 0.06742f
C4937 top_DAC_0/top_rseg_n_dcell_0.VL3.t1 GND 0.01949f
C4938 top_DAC_0/top_rseg_n_dcell_0.VL3.n5 GND 0.13298f
C4939 top_DAC_0/top_rseg_n_dcell_0.SH[3].t0 GND 0.11227f
C4940 top_DAC_0/top_rseg_n_dcell_0.SH[3].n0 GND 0.04603f
C4941 top_DAC_0/top_rseg_n_dcell_0.SH[3].n1 GND 0.09909f
C4942 top_DAC_0/top_rseg_n_dcell_0.SH[3].n2 GND 0.06579f
C4943 top_DAC_0/top_rseg_n_dcell_0.SH[3].t1 GND 0.10756f
C4944 top_DAC_0/top_rseg_n_dcell_0.SH[3].n3 GND 0.01359f
C4945 top_DAC_0/top_rseg_n_dcell_0.SH[3].t3 GND 0.22037f
C4946 top_DAC_0/top_rseg_n_dcell_0.SH[3].t6 GND 0.2195f
C4947 top_DAC_0/top_rseg_n_dcell_0.SH[3].n4 GND 0.42193f
C4948 top_DAC_0/top_rseg_n_dcell_0.SH[3].t4 GND 0.2195f
C4949 top_DAC_0/top_rseg_n_dcell_0.SH[3].n5 GND 0.23437f
C4950 top_DAC_0/top_rseg_n_dcell_0.SH[3].t2 GND 0.2195f
C4951 top_DAC_0/top_rseg_n_dcell_0.SH[3].n6 GND 0.23437f
C4952 top_DAC_0/top_rseg_n_dcell_0.SH[3].t5 GND 0.2195f
C4953 top_DAC_0/top_rseg_n_dcell_0.SH[3].n7 GND 0.25474f
C4954 top_DAC_0/top_rseg_n_dcell_0.SH[3].n8 GND 0.07619f
C4955 a_31870_7686.t2 GND 0.05828f
C4956 a_31870_7686.t1 GND 0.04276f
C4957 a_31870_7686.n0 GND 2.03892f
C4958 a_31870_7686.t4 GND 0.04087f
C4959 a_31870_7686.n1 GND 1.29976f
C4960 a_31870_7686.t3 GND 0.07543f
C4961 a_31870_7686.n2 GND 3.00311f
C4962 a_31870_7686.t0 GND 0.04087f
C4963 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.t0 GND 0.03703f
C4964 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.t2 GND 0.12366f
C4965 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.t1 GND 0.36626f
C4966 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56.n0 GND 2.56502f
C4967 a_29780_7686.t1 GND 0.04115f
C4968 a_29780_7686.t2 GND 0.05703f
C4969 a_29780_7686.n0 GND 1.94212f
C4970 a_29780_7686.t3 GND 0.03868f
C4971 a_29780_7686.n1 GND 1.52384f
C4972 a_29780_7686.t4 GND 0.06894f
C4973 a_29780_7686.n2 GND 2.78956f
C4974 a_29780_7686.t0 GND 0.03868f
C4975 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t1 GND 0.08336f
C4976 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t0 GND 0.09794f
C4977 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n0 GND 0.50552f
C4978 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t9 GND 0.38933f
C4979 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t22 GND 0.38769f
C4980 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n1 GND 0.65162f
C4981 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t3 GND 0.38769f
C4982 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n2 GND 0.57279f
C4983 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n3 GND 0.8829f
C4984 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t6 GND 0.11878f
C4985 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t16 GND 0.11718f
C4986 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n4 GND 7.32954f
C4987 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t15 GND 0.11915f
C4988 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t11 GND 0.11855f
C4989 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n5 GND 0.38612f
C4990 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t21 GND 0.11855f
C4991 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n6 GND 0.19336f
C4992 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t14 GND 0.11855f
C4993 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n7 GND 0.19336f
C4994 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t24 GND 0.11855f
C4995 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n8 GND 0.19336f
C4996 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t20 GND 0.11855f
C4997 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n9 GND 0.19336f
C4998 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t23 GND 0.11855f
C4999 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n10 GND 0.19336f
C5000 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t2 GND 0.11718f
C5001 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t5 GND 0.11915f
C5002 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t17 GND 0.11954f
C5003 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t12 GND 0.11889f
C5004 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n11 GND 0.41817f
C5005 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t10 GND 0.11889f
C5006 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n12 GND 0.20941f
C5007 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t7 GND 0.11889f
C5008 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n13 GND 0.20941f
C5009 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t13 GND 0.11889f
C5010 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n14 GND 0.20941f
C5011 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t4 GND 0.11889f
C5012 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n15 GND 0.20941f
C5013 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n16 GND 0.32292f
C5014 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t8 GND 0.11718f
C5015 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n17 GND 0.40691f
C5016 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n18 GND 0.38834f
C5017 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n19 GND 0.09562f
C5018 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n20 GND 10.423f
C5019 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t18 GND 0.22031f
C5020 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].t19 GND 0.12221f
C5021 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n21 GND 0.19198f
C5022 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n22 GND 0.03351f
C5023 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3].n23 GND 0.26224f
C5024 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t1 GND 0.12074f
C5025 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t0 GND 0.12074f
C5026 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t2 GND 0.12074f
C5027 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n0 GND 0.65062f
C5028 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t4 GND 0.13368f
C5029 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t6 GND 0.13005f
C5030 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n1 GND 1.04458f
C5031 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t7 GND 0.13368f
C5032 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t5 GND 0.13005f
C5033 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n2 GND 0.85678f
C5034 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n3 GND 1.00824f
C5035 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n4 GND 0.9243f
C5036 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n5 GND 0.70506f
C5037 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t3 GND 0.12074f
C5038 top_DAC_0/top_final_switch_0.VOUT[4].n0 GND 0.02064f
C5039 top_DAC_0/top_final_switch_0.VOUT[4].n1 GND 0.02156f
C5040 top_DAC_0/top_final_switch_0.VOUT[4].n2 GND 1.24183f
C5041 top_DAC_0/top_final_switch_0.VOUT[4].t9 GND 0.84393f
C5042 top_DAC_0/top_final_switch_0.VOUT[4].t7 GND 0.83868f
C5043 top_DAC_0/top_final_switch_0.VOUT[4].n3 GND 1.39936f
C5044 top_DAC_0/top_final_switch_0.VOUT[4].t11 GND 0.83923f
C5045 top_DAC_0/top_final_switch_0.VOUT[4].t5 GND 0.8377f
C5046 top_DAC_0/top_final_switch_0.VOUT[4].n4 GND 1.08055f
C5047 top_DAC_0/top_final_switch_0.VOUT[4].n5 GND 0.70544f
C5048 top_DAC_0/top_final_switch_0.VOUT[4].t10 GND 0.3448f
C5049 top_DAC_0/top_final_switch_0.VOUT[4].t4 GND 0.34313f
C5050 top_DAC_0/top_final_switch_0.VOUT[4].n6 GND 0.91129f
C5051 top_DAC_0/top_final_switch_0.VOUT[4].t8 GND 0.35048f
C5052 top_DAC_0/top_final_switch_0.VOUT[4].t6 GND 0.34456f
C5053 top_DAC_0/top_final_switch_0.VOUT[4].n7 GND 1.01506f
C5054 top_DAC_0/top_final_switch_0.VOUT[4].n8 GND 0.53226f
C5055 top_DAC_0/top_final_switch_0.VOUT[4].n9 GND 0.18412f
C5056 top_DAC_0/top_final_switch_0.VOUT[4].n10 GND 0.53867f
C5057 top_DAC_0/top_final_switch_0.VOUT[4].n11 GND 0.2628f
C5058 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.t1 GND 0.02587f
C5059 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.t2 GND 0.07997f
C5060 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.t0 GND 0.07985f
C5061 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12.n0 GND 1.3573f
C5062 a_5050_12595.t7 GND 0.02366f
C5063 a_5050_12595.t9 GND 0.02366f
C5064 a_5050_12595.t1 GND 0.02366f
C5065 a_5050_12595.n0 GND 0.05487f
C5066 a_5050_12595.t0 GND 0.02366f
C5067 a_5050_12595.t8 GND 0.02366f
C5068 a_5050_12595.n1 GND 0.05487f
C5069 a_5050_12595.n2 GND 0.40357f
C5070 a_5050_12595.t4 GND 0.11399f
C5071 a_5050_12595.t5 GND 0.12455f
C5072 a_5050_12595.n3 GND 5.31895f
C5073 a_5050_12595.n4 GND 0.32667f
C5074 a_5050_12595.t6 GND 0.02366f
C5075 a_5050_12595.t2 GND 0.02366f
C5076 a_5050_12595.n5 GND 0.05487f
C5077 a_5050_12595.n6 GND 0.40357f
C5078 a_5050_12595.n7 GND 0.05487f
C5079 a_5050_12595.t3 GND 0.02366f
C5080 top_DAC_0/top_final_switch_0.VOUT[0].n0 GND 0.01656f
C5081 top_DAC_0/top_final_switch_0.VOUT[0].n1 GND 0.01729f
C5082 top_DAC_0/top_final_switch_0.VOUT[0].n2 GND 0.98633f
C5083 top_DAC_0/top_final_switch_0.VOUT[0].t7 GND 0.67691f
C5084 top_DAC_0/top_final_switch_0.VOUT[0].t5 GND 0.6727f
C5085 top_DAC_0/top_final_switch_0.VOUT[0].n3 GND 1.12242f
C5086 top_DAC_0/top_final_switch_0.VOUT[0].t11 GND 0.67314f
C5087 top_DAC_0/top_final_switch_0.VOUT[0].t10 GND 0.67191f
C5088 top_DAC_0/top_final_switch_0.VOUT[0].n4 GND 0.8667f
C5089 top_DAC_0/top_final_switch_0.VOUT[0].n5 GND 0.62892f
C5090 top_DAC_0/top_final_switch_0.VOUT[0].t9 GND 0.27656f
C5091 top_DAC_0/top_final_switch_0.VOUT[0].t8 GND 0.27523f
C5092 top_DAC_0/top_final_switch_0.VOUT[0].n6 GND 0.73094f
C5093 top_DAC_0/top_final_switch_0.VOUT[0].t6 GND 0.28112f
C5094 top_DAC_0/top_final_switch_0.VOUT[0].t4 GND 0.27637f
C5095 top_DAC_0/top_final_switch_0.VOUT[0].n7 GND 0.81417f
C5096 top_DAC_0/top_final_switch_0.VOUT[0].n8 GND 0.36383f
C5097 top_DAC_0/top_final_switch_0.VOUT[0].n9 GND 1.09627f
C5098 top_DAC_0/top_final_switch_0.VOUT[0].n10 GND 0.19303f
C5099 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.t2 GND 0.01519f
C5100 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.t1 GND 0.08976f
C5101 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.n0 GND 1.90489f
C5102 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23.t0 GND 0.09016f
C5103 a_24963_20174.t1 GND 0.15594f
C5104 a_24963_20174.t3 GND 0.06377f
C5105 a_24963_20174.n0 GND 5.11593f
C5106 a_24963_20174.t2 GND 0.06506f
C5107 a_24963_20174.n1 GND 3.89706f
C5108 a_24963_20174.t0 GND 0.10224f
C5109 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t2 GND 0.14561f
C5110 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n0 GND 0.18624f
C5111 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t13 GND 0.14561f
C5112 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n1 GND 0.23751f
C5113 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t7 GND 0.14561f
C5114 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n2 GND 0.23751f
C5115 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t19 GND 0.14561f
C5116 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n3 GND 0.23751f
C5117 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t12 GND 0.14561f
C5118 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n4 GND 0.23751f
C5119 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t21 GND 0.14561f
C5120 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n5 GND 0.23751f
C5121 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t17 GND 0.14561f
C5122 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n6 GND 0.23751f
C5123 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t8 GND 0.14561f
C5124 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n7 GND 0.22308f
C5125 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t15 GND 0.14635f
C5126 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t5 GND 0.14561f
C5127 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n8 GND 0.47428f
C5128 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t11 GND 0.14561f
C5129 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n9 GND 0.23751f
C5130 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t16 GND 0.14561f
C5131 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n10 GND 0.23751f
C5132 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t6 GND 0.14561f
C5133 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n11 GND 0.23751f
C5134 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t18 GND 0.14561f
C5135 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n12 GND 0.23751f
C5136 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t4 GND 0.14561f
C5137 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n13 GND 0.23751f
C5138 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t10 GND 0.14561f
C5139 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n14 GND 0.23751f
C5140 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t20 GND 0.14561f
C5141 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n15 GND 0.17196f
C5142 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n16 GND 16.048f
C5143 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t0 GND 0.1204f
C5144 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t1 GND 0.10238f
C5145 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n17 GND 0.82365f
C5146 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t3 GND 0.47802f
C5147 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t14 GND 0.47604f
C5148 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n18 GND 0.75563f
C5149 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n19 GND 0.48747f
C5150 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].t9 GND 0.50273f
C5151 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1].n20 GND 1.05121f
C5152 a_36888_19550.t2 GND 0.05539f
C5153 a_36888_19550.t3 GND 0.05331f
C5154 a_36888_19550.n0 GND 0.5884f
C5155 a_36888_19550.t1 GND 0.09815f
C5156 a_36888_19550.n1 GND 1.64869f
C5157 a_36888_19550.t0 GND 0.05605f
C5158 a_36888_19786.t5 GND 0.03016f
C5159 a_36888_19786.t4 GND 0.14825f
C5160 a_36888_19786.n0 GND 0.16973f
C5161 a_36888_19786.t7 GND 0.15058f
C5162 a_36888_19786.n1 GND 0.279f
C5163 a_36888_19786.t6 GND 0.15058f
C5164 a_36888_19786.t2 GND 0.14825f
C5165 a_36888_19786.t3 GND 0.03016f
C5166 a_36888_19786.n2 GND 0.16973f
C5167 a_36888_19786.n3 GND 0.29912f
C5168 a_36888_19786.t1 GND 0.03278f
C5169 a_36888_19786.n4 GND 0.83928f
C5170 a_36888_19786.t0 GND 0.05237f
C5171 a_31042_7686.t4 GND 0.10032f
C5172 a_31042_7686.t1 GND 0.08434f
C5173 a_31042_7686.n0 GND 3.60497f
C5174 a_31042_7686.t3 GND 0.07983f
C5175 a_31042_7686.n1 GND 2.75522f
C5176 a_31042_7686.t2 GND 0.14569f
C5177 a_31042_7686.n2 GND 5.84981f
C5178 a_31042_7686.t0 GND 0.07983f
C5179 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t0 GND 0.10226f
C5180 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t1 GND 0.08695f
C5181 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n0 GND 0.69951f
C5182 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t18 GND 0.40597f
C5183 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t23 GND 0.4043f
C5184 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n1 GND 0.64174f
C5185 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n2 GND 0.414f
C5186 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t24 GND 0.42696f
C5187 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n3 GND 0.89278f
C5188 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t4 GND 0.12394f
C5189 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t13 GND 0.12224f
C5190 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n4 GND 5.66133f
C5191 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t3 GND 0.12429f
C5192 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t5 GND 0.12366f
C5193 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n5 GND 0.4028f
C5194 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t22 GND 0.12366f
C5195 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n6 GND 0.20171f
C5196 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t2 GND 0.12366f
C5197 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n7 GND 0.20171f
C5198 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t15 GND 0.12366f
C5199 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n8 GND 0.20171f
C5200 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t7 GND 0.12366f
C5201 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n9 GND 0.20171f
C5202 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t10 GND 0.12366f
C5203 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n10 GND 0.20171f
C5204 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n11 GND 0.09544f
C5205 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t14 GND 0.12224f
C5206 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n12 GND 0.10215f
C5207 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t12 GND 0.12429f
C5208 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t20 GND 0.12471f
C5209 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t19 GND 0.12403f
C5210 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n13 GND 0.43623f
C5211 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t17 GND 0.12403f
C5212 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n14 GND 0.21846f
C5213 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t21 GND 0.12403f
C5214 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n15 GND 0.21846f
C5215 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t11 GND 0.12403f
C5216 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n16 GND 0.21846f
C5217 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t8 GND 0.12403f
C5218 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n17 GND 0.21846f
C5219 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n18 GND 0.33687f
C5220 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t16 GND 0.12224f
C5221 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n19 GND 0.42787f
C5222 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n20 GND 2.49587f
C5223 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n21 GND 11.4725f
C5224 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t6 GND 0.22982f
C5225 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].t9 GND 0.12749f
C5226 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n22 GND 0.20027f
C5227 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n23 GND 0.03496f
C5228 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1].n24 GND 0.27468f
C5229 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t0 GND 0.09672f
C5230 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n0 GND 0.03966f
C5231 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n1 GND 0.08537f
C5232 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n2 GND 0.05668f
C5233 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t1 GND 0.09266f
C5234 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n3 GND 0.0117f
C5235 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t2 GND 0.19122f
C5236 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n4 GND 0.24119f
C5237 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t4 GND 0.19213f
C5238 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n5 GND 0.49912f
C5239 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t6 GND 0.18909f
C5240 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n6 GND 14.5942f
C5241 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t3 GND 0.33825f
C5242 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].t5 GND 0.18764f
C5243 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n7 GND 0.29475f
C5244 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n8 GND 0.05864f
C5245 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4].n9 GND 0.08407f
C5246 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t23 GND 2.65181f
C5247 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t5 GND 0.10532f
C5248 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t4 GND 0.39669f
C5249 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n0 GND 0.35115f
C5250 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t2 GND 0.39669f
C5251 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n1 GND 0.16403f
C5252 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t3 GND 0.10454f
C5253 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n2 GND 0.19634f
C5254 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n3 GND 0.89301f
C5255 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t1 GND 0.03518f
C5256 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t0 GND 0.04509f
C5257 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n4 GND 0.51038f
C5258 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t11 GND 0.2035f
C5259 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t15 GND 0.20271f
C5260 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n5 GND 0.41896f
C5261 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t19 GND 0.20271f
C5262 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n6 GND 0.17856f
C5263 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t20 GND 0.20271f
C5264 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n7 GND 0.17856f
C5265 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t6 GND 0.20271f
C5266 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n8 GND 0.17856f
C5267 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t26 GND 0.20271f
C5268 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n9 GND 0.17856f
C5269 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t12 GND 0.20271f
C5270 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n10 GND 0.17856f
C5271 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t14 GND 0.20271f
C5272 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n11 GND 0.17856f
C5273 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t22 GND 0.20271f
C5274 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n12 GND 0.17856f
C5275 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t25 GND 0.20271f
C5276 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n13 GND 0.17856f
C5277 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t28 GND 0.20271f
C5278 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n14 GND 0.17856f
C5279 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t8 GND 0.20271f
C5280 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n15 GND 0.17856f
C5281 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t10 GND 0.20271f
C5282 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n16 GND 0.17856f
C5283 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t16 GND 0.20271f
C5284 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n17 GND 0.17856f
C5285 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t18 GND 0.20271f
C5286 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n18 GND 0.17856f
C5287 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t21 GND 0.20271f
C5288 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n19 GND 0.17856f
C5289 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t24 GND 0.20271f
C5290 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n20 GND 0.17856f
C5291 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t27 GND 0.20271f
C5292 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n21 GND 0.17856f
C5293 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t7 GND 0.20271f
C5294 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n22 GND 0.17856f
C5295 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t9 GND 0.20271f
C5296 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n23 GND 0.17856f
C5297 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t13 GND 0.20271f
C5298 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n24 GND 0.17856f
C5299 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t17 GND 0.20271f
C5300 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n25 GND 0.16737f
C5301 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n26 GND 1.68902f
C5302 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n27 GND 2.3067f
C5303 a_6923_9707.t4 GND 0.05554f
C5304 a_6923_9707.t1 GND 0.05553f
C5305 a_6923_9707.n0 GND 0.75856f
C5306 a_6923_9707.n1 GND 0.61998f
C5307 a_6923_9707.t5 GND 0.05546f
C5308 a_6923_9707.n2 GND 0.2593f
C5309 a_6923_9707.t15 GND 0.05546f
C5310 a_6923_9707.n3 GND 0.2593f
C5311 a_6923_9707.n4 GND 0.39892f
C5312 a_6923_9707.n5 GND 0.39892f
C5313 a_6923_9707.t12 GND 0.02477f
C5314 a_6923_9707.t23 GND 0.02477f
C5315 a_6923_9707.n6 GND 0.05745f
C5316 a_6923_9707.t20 GND 0.02477f
C5317 a_6923_9707.t13 GND 0.02477f
C5318 a_6923_9707.n7 GND 0.05745f
C5319 a_6923_9707.n8 GND 0.42255f
C5320 a_6923_9707.t22 GND 0.02477f
C5321 a_6923_9707.t11 GND 0.02477f
C5322 a_6923_9707.n9 GND 0.05745f
C5323 a_6923_9707.t14 GND 0.02477f
C5324 a_6923_9707.t21 GND 0.02477f
C5325 a_6923_9707.n10 GND 0.05745f
C5326 a_6923_9707.n11 GND 0.42255f
C5327 a_6923_9707.n12 GND 0.12609f
C5328 a_6923_9707.t3 GND 0.05546f
C5329 a_6923_9707.n13 GND 0.26103f
C5330 a_6923_9707.t16 GND 0.05553f
C5331 a_6923_9707.t2 GND 0.05554f
C5332 a_6923_9707.n14 GND 0.75856f
C5333 a_6923_9707.n15 GND 0.61998f
C5334 a_6923_9707.t6 GND 0.05546f
C5335 a_6923_9707.t10 GND 0.05546f
C5336 a_6923_9707.n16 GND 0.2593f
C5337 a_6923_9707.n17 GND 0.2593f
C5338 a_6923_9707.n18 GND 0.39892f
C5339 a_6923_9707.n19 GND 0.39892f
C5340 a_6923_9707.t17 GND 0.05546f
C5341 a_6923_9707.t9 GND 0.05546f
C5342 a_6923_9707.n20 GND 0.2593f
C5343 a_6923_9707.n21 GND 0.2593f
C5344 a_6923_9707.n22 GND 0.39892f
C5345 a_6923_9707.t19 GND 0.05546f
C5346 a_6923_9707.n23 GND 0.2593f
C5347 a_6923_9707.n24 GND 0.37714f
C5348 a_6923_9707.n25 GND 0.08229f
C5349 a_6923_9707.n26 GND 1.80716f
C5350 a_6923_9707.n27 GND 0.58376f
C5351 a_6923_9707.t18 GND 0.05546f
C5352 a_6923_9707.n28 GND 0.2593f
C5353 a_6923_9707.t8 GND 0.05546f
C5354 a_6923_9707.n29 GND 0.2593f
C5355 a_6923_9707.n30 GND 0.39892f
C5356 a_6923_9707.n31 GND 0.39892f
C5357 a_6923_9707.t7 GND 0.05546f
C5358 a_6923_9707.n32 GND 0.2593f
C5359 a_6923_9707.n33 GND 0.2593f
C5360 a_6923_9707.t0 GND 0.05546f
C5361 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t3 GND 0.52048f
C5362 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t1 GND 0.44012f
C5363 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t0 GND 0.46157f
C5364 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n0 GND 2.31307f
C5365 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n1 GND 1.44843f
C5366 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t21 GND 0.02401f
C5367 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t20 GND 0.02401f
C5368 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n2 GND 0.05274f
C5369 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t23 GND 0.08557f
C5370 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t13 GND 0.02401f
C5371 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t12 GND 0.02401f
C5372 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n3 GND 0.05274f
C5373 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t15 GND 0.08557f
C5374 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t4 GND 0.02401f
C5375 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t7 GND 0.02401f
C5376 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n4 GND 0.05274f
C5377 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t5 GND 0.08557f
C5378 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t8 GND 0.02401f
C5379 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t10 GND 0.02401f
C5380 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n5 GND 0.05274f
C5381 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t11 GND 0.08557f
C5382 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t19 GND 0.02401f
C5383 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t16 GND 0.02401f
C5384 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n6 GND 0.05274f
C5385 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t18 GND 0.12216f
C5386 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n7 GND 0.84523f
C5387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t17 GND 0.0856f
C5388 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n8 GND 0.32109f
C5389 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n9 GND 0.33237f
C5390 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n10 GND 0.42678f
C5391 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n11 GND 0.54022f
C5392 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t9 GND 0.0856f
C5393 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n12 GND 0.32109f
C5394 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n13 GND 0.33237f
C5395 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n14 GND 0.42678f
C5396 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n15 GND 0.54022f
C5397 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t6 GND 0.0856f
C5398 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n16 GND 0.32109f
C5399 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n17 GND 0.33237f
C5400 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n18 GND 0.42678f
C5401 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n19 GND 0.54022f
C5402 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t14 GND 0.0856f
C5403 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n20 GND 0.32109f
C5404 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n21 GND 0.33237f
C5405 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n22 GND 0.42678f
C5406 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n23 GND 0.54022f
C5407 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t22 GND 0.0856f
C5408 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n24 GND 0.32109f
C5409 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n25 GND 2.14651f
C5410 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t2 GND 0.52116f
C5411 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n26 GND 3.06731f
C5412 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t0 GND 0.08748f
C5413 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t36 GND 0.0844f
C5414 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n0 GND 1.3512f
C5415 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t34 GND 0.0844f
C5416 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n1 GND 0.72881f
C5417 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t6 GND 0.08748f
C5418 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t7 GND 0.08248f
C5419 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t38 GND 0.07822f
C5420 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n2 GND 1.08605f
C5421 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t3 GND 0.07822f
C5422 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n3 GND 0.46201f
C5423 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n4 GND 1.08984f
C5424 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t39 GND 0.0844f
C5425 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n5 GND 0.82131f
C5426 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t11 GND 0.0844f
C5427 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n6 GND 0.82131f
C5428 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t10 GND 0.0844f
C5429 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n7 GND 0.68473f
C5430 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n8 GND 0.57528f
C5431 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t4 GND 0.08748f
C5432 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t35 GND 0.08248f
C5433 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t12 GND 0.07822f
C5434 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n9 GND 1.08605f
C5435 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t5 GND 0.07822f
C5436 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n10 GND 0.46201f
C5437 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n11 GND 1.08984f
C5438 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t33 GND 0.0844f
C5439 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n12 GND 0.82131f
C5440 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t2 GND 0.0844f
C5441 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n13 GND 0.68617f
C5442 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t37 GND 0.08748f
C5443 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t8 GND 0.0844f
C5444 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n14 GND 1.3512f
C5445 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t1 GND 0.0844f
C5446 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n15 GND 0.82131f
C5447 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t9 GND 0.0844f
C5448 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n16 GND 0.64209f
C5449 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n17 GND 0.31437f
C5450 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n18 GND 1.77552f
C5451 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t32 GND 0.07826f
C5452 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t20 GND 0.07832f
C5453 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t29 GND 0.07822f
C5454 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n19 GND 0.41842f
C5455 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t31 GND 0.07822f
C5456 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n20 GND 0.19934f
C5457 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n21 GND 0.57069f
C5458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t13 GND 0.07826f
C5459 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t22 GND 0.07826f
C5460 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n22 GND 0.47705f
C5461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n23 GND 1.18839f
C5462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t26 GND 0.07826f
C5463 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t18 GND 0.07826f
C5464 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n24 GND 0.70457f
C5465 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t25 GND 0.07826f
C5466 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t24 GND 0.07826f
C5467 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n25 GND 0.47705f
C5468 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n26 GND 1.14431f
C5469 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n27 GND 0.71001f
C5470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t30 GND 0.07826f
C5471 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t21 GND 0.07826f
C5472 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n28 GND 0.70457f
C5473 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t28 GND 0.07826f
C5474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t17 GND 0.07826f
C5475 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n29 GND 0.47705f
C5476 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n30 GND 0.91667f
C5477 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t27 GND 0.07832f
C5478 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t19 GND 0.07822f
C5479 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n31 GND 0.41842f
C5480 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t16 GND 0.07822f
C5481 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n32 GND 0.19934f
C5482 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t15 GND 0.07826f
C5483 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n33 GND 0.57069f
C5484 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t23 GND 0.07826f
C5485 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t14 GND 0.07826f
C5486 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n34 GND 0.47705f
C5487 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n35 GND 1.41604f
C5488 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n36 GND 0.54346f
C5489 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n37 GND 1.19678f
C5490 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.t2 GND 0.10196f
C5491 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.t1 GND 0.09876f
C5492 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.n0 GND 1.88582f
C5493 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36.t0 GND 0.01345f
C5494 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t14 GND 0.14295f
C5495 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t6 GND 0.14218f
C5496 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n0 GND 0.50006f
C5497 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t18 GND 0.14218f
C5498 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n1 GND 0.25042f
C5499 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t4 GND 0.14218f
C5500 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n2 GND 0.22448f
C5501 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t5 GND 0.14218f
C5502 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n3 GND 0.19854f
C5503 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t15 GND 0.14218f
C5504 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n4 GND 0.25042f
C5505 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t2 GND 0.14218f
C5506 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n5 GND 0.25042f
C5507 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t17 GND 0.14218f
C5508 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n6 GND 0.23356f
C5509 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t8 GND 0.14295f
C5510 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t12 GND 0.14218f
C5511 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n7 GND 0.50006f
C5512 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t19 GND 0.14218f
C5513 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n8 GND 0.25042f
C5514 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t9 GND 0.14218f
C5515 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n9 GND 0.25042f
C5516 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t20 GND 0.14218f
C5517 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n10 GND 0.25042f
C5518 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t3 GND 0.14218f
C5519 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n11 GND 0.25042f
C5520 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t11 GND 0.14218f
C5521 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n12 GND 0.25042f
C5522 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t21 GND 0.14218f
C5523 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n13 GND 0.25042f
C5524 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t13 GND 0.14218f
C5525 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n14 GND 0.1892f
C5526 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n15 GND 14.7419f
C5527 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t10 GND 0.4559f
C5528 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t1 GND 0.09968f
C5529 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t0 GND 0.11713f
C5530 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n16 GND 0.6449f
C5531 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n17 GND 0.51336f
C5532 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t16 GND 0.46557f
C5533 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].t7 GND 0.46361f
C5534 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n18 GND 1.03065f
C5535 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2].n19 GND 0.7664f
C5536 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t5 GND 0.16429f
C5537 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t9 GND 0.16346f
C5538 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n0 GND 0.47064f
C5539 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t8 GND 0.16429f
C5540 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t4 GND 0.16346f
C5541 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n1 GND 0.53242f
C5542 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n2 GND 0.15152f
C5543 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t6 GND 0.16158f
C5544 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n3 GND 15.2195f
C5545 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t1 GND 0.11495f
C5546 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t0 GND 0.13506f
C5547 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n4 GND 0.69706f
C5548 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t7 GND 0.53685f
C5549 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t3 GND 0.53459f
C5550 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n5 GND 0.89852f
C5551 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].t2 GND 0.53459f
C5552 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n6 GND 0.78982f
C5553 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3].n7 GND 1.21743f
C5554 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t6 GND 0.17266f
C5555 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t3 GND 0.17211f
C5556 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n0 GND 0.24239f
C5557 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t8 GND 0.17306f
C5558 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t5 GND 0.17211f
C5559 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n1 GND 0.60536f
C5560 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n2 GND 0.18843f
C5561 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t9 GND 0.16963f
C5562 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n3 GND 16.2245f
C5563 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t2 GND 0.5519f
C5564 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t1 GND 0.12067f
C5565 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t0 GND 0.14179f
C5566 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n4 GND 0.78071f
C5567 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n5 GND 0.62147f
C5568 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t7 GND 0.56361f
C5569 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].t4 GND 0.56124f
C5570 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n6 GND 1.24769f
C5571 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2].n7 GND 0.92779f
C5572 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.t1 GND -0.04304f
C5573 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.t0 GND -0.04297f
C5574 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20.n0 GND -0.74313f
C5575 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t5 GND 0.33461f
C5576 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t4 GND 0.44915f
C5577 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t3 GND 0.33244f
C5578 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n0 GND 1.43209f
C5579 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t0 GND 0.45383f
C5580 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n1 GND 1.80141f
C5581 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n2 GND 1.63754f
C5582 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t9 GND 0.70064f
C5583 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t6 GND 0.69977f
C5584 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n3 GND 0.57765f
C5585 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t7 GND 0.70064f
C5586 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t8 GND 0.69977f
C5587 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n4 GND 0.57802f
C5588 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n5 GND 0.37137f
C5589 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n6 GND 0.42971f
C5590 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t1 GND 0.10481f
C5591 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.t2 GND 0.15924f
C5592 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A.n7 GND 1.27737f
C5593 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t2 GND 0.03483f
C5594 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t0 GND 0.03483f
C5595 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n0 GND 0.07139f
C5596 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n1 GND 0.36157f
C5597 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t10 GND 0.49404f
C5598 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t68 GND 0.49225f
C5599 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n2 GND 0.65036f
C5600 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t44 GND 0.49225f
C5601 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n3 GND 0.32608f
C5602 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t8 GND 0.49225f
C5603 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n4 GND 0.32608f
C5604 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t64 GND 0.49225f
C5605 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n5 GND 0.32608f
C5606 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t65 GND 0.49225f
C5607 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n6 GND 0.32608f
C5608 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t16 GND 0.49225f
C5609 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n7 GND 0.32608f
C5610 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t66 GND 0.49225f
C5611 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n8 GND 0.32608f
C5612 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t30 GND 0.49225f
C5613 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n9 GND 0.32608f
C5614 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t34 GND 0.49225f
C5615 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n10 GND 0.32608f
C5616 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t6 GND 0.49225f
C5617 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n11 GND 0.32608f
C5618 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t47 GND 0.49225f
C5619 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n12 GND 0.25142f
C5620 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t26 GND 0.49404f
C5621 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t42 GND 0.49225f
C5622 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n13 GND 0.65036f
C5623 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t9 GND 0.49225f
C5624 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n14 GND 0.32608f
C5625 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t7 GND 0.49225f
C5626 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n15 GND 0.32608f
C5627 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t43 GND 0.49225f
C5628 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n16 GND 0.32608f
C5629 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t67 GND 0.49225f
C5630 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n17 GND 0.32608f
C5631 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t5 GND 0.49225f
C5632 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n18 GND 0.32608f
C5633 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t25 GND 0.49225f
C5634 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n19 GND 0.32548f
C5635 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n20 GND 0.12706f
C5636 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t77 GND 0.49404f
C5637 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t56 GND 0.49225f
C5638 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n21 GND 0.65036f
C5639 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t29 GND 0.49225f
C5640 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n22 GND 0.32608f
C5641 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t74 GND 0.49225f
C5642 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n23 GND 0.32608f
C5643 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t45 GND 0.49225f
C5644 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n24 GND 0.32608f
C5645 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t46 GND 0.49225f
C5646 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n25 GND 0.32608f
C5647 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t84 GND 0.49225f
C5648 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n26 GND 0.32608f
C5649 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t49 GND 0.49225f
C5650 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n27 GND 0.32608f
C5651 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t19 GND 0.49225f
C5652 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n28 GND 0.32608f
C5653 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t20 GND 0.49225f
C5654 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n29 GND 0.32608f
C5655 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t70 GND 0.49225f
C5656 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n30 GND 0.32608f
C5657 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t37 GND 0.49225f
C5658 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n31 GND 0.25142f
C5659 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t14 GND 0.49404f
C5660 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t27 GND 0.49225f
C5661 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n32 GND 0.65036f
C5662 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t76 GND 0.49225f
C5663 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n33 GND 0.32608f
C5664 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t71 GND 0.49225f
C5665 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n34 GND 0.32608f
C5666 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t28 GND 0.49225f
C5667 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n35 GND 0.32608f
C5668 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t53 GND 0.49225f
C5669 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n36 GND 0.32608f
C5670 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t69 GND 0.49225f
C5671 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n37 GND 0.32608f
C5672 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t11 GND 0.49225f
C5673 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n38 GND 0.32548f
C5674 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n39 GND 0.07526f
C5675 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n40 GND 0.58913f
C5676 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t83 GND 0.49404f
C5677 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t61 GND 0.49225f
C5678 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n41 GND 0.65036f
C5679 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t35 GND 0.49225f
C5680 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n42 GND 0.32608f
C5681 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t80 GND 0.49225f
C5682 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n43 GND 0.32608f
C5683 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t48 GND 0.49225f
C5684 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n44 GND 0.32608f
C5685 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t50 GND 0.49225f
C5686 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n45 GND 0.32608f
C5687 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t86 GND 0.49225f
C5688 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n46 GND 0.32608f
C5689 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t52 GND 0.49225f
C5690 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n47 GND 0.32608f
C5691 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t21 GND 0.49225f
C5692 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n48 GND 0.32608f
C5693 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t23 GND 0.49225f
C5694 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n49 GND 0.32608f
C5695 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t75 GND 0.49225f
C5696 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n50 GND 0.32608f
C5697 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t39 GND 0.49225f
C5698 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n51 GND 0.25142f
C5699 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t18 GND 0.49404f
C5700 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t31 GND 0.49225f
C5701 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n52 GND 0.65036f
C5702 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t81 GND 0.49225f
C5703 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n53 GND 0.32608f
C5704 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t78 GND 0.49225f
C5705 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n54 GND 0.32608f
C5706 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t32 GND 0.49225f
C5707 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n55 GND 0.32608f
C5708 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t57 GND 0.49225f
C5709 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n56 GND 0.32608f
C5710 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t73 GND 0.49225f
C5711 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n57 GND 0.32608f
C5712 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t13 GND 0.49225f
C5713 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n58 GND 0.32548f
C5714 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n59 GND 0.07526f
C5715 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n60 GND 0.37231f
C5716 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t60 GND 0.49404f
C5717 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t41 GND 0.49225f
C5718 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n61 GND 0.65036f
C5719 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t17 GND 0.49225f
C5720 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n62 GND 0.32608f
C5721 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t58 GND 0.49225f
C5722 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n63 GND 0.32608f
C5723 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t33 GND 0.49225f
C5724 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n64 GND 0.32608f
C5725 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t36 GND 0.49225f
C5726 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n65 GND 0.32608f
C5727 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t63 GND 0.49225f
C5728 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n66 GND 0.32608f
C5729 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t38 GND 0.49225f
C5730 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n67 GND 0.32608f
C5731 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t85 GND 0.49225f
C5732 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n68 GND 0.32608f
C5733 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t87 GND 0.49225f
C5734 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n69 GND 0.32608f
C5735 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t54 GND 0.49225f
C5736 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n70 GND 0.32608f
C5737 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t22 GND 0.49225f
C5738 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n71 GND 0.25142f
C5739 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t62 GND 1.13006f
C5740 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t4 GND 1.12853f
C5741 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n72 GND 0.96689f
C5742 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t82 GND 1.13006f
C5743 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t24 GND 1.12853f
C5744 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n73 GND 1.14066f
C5745 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n74 GND 0.56996f
C5746 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t79 GND 0.49225f
C5747 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n75 GND 0.6695f
C5748 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t12 GND 0.49225f
C5749 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n76 GND 0.32608f
C5750 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t59 GND 0.49225f
C5751 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n77 GND 0.32608f
C5752 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t55 GND 0.49225f
C5753 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n78 GND 0.32608f
C5754 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t15 GND 0.49225f
C5755 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n79 GND 0.32608f
C5756 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t40 GND 0.49225f
C5757 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n80 GND 0.32608f
C5758 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t51 GND 0.49225f
C5759 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n81 GND 0.32608f
C5760 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t72 GND 0.49225f
C5761 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n82 GND 0.32548f
C5762 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n83 GND 0.07526f
C5763 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n84 GND 1.44386f
C5764 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t1 GND 0.03483f
C5765 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.t3 GND 0.03483f
C5766 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n85 GND 0.07139f
C5767 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n86 GND 0.46009f
C5768 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2.n87 GND 0.53996f
C5769 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t2 GND 0.04329f
C5770 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t3 GND 0.04329f
C5771 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n0 GND 0.09506f
C5772 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n1 GND 0.04101f
C5773 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t4 GND 0.04474f
C5774 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t17 GND 0.07165f
C5775 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n2 GND 0.13662f
C5776 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n3 GND 0.1482f
C5777 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n4 GND 0.5264f
C5778 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t6 GND 0.07295f
C5779 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t10 GND 0.04581f
C5780 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n5 GND 0.09982f
C5781 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n6 GND 0.12298f
C5782 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t8 GND 0.07295f
C5783 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t14 GND 0.04581f
C5784 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n7 GND 0.11271f
C5785 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n8 GND 0.15523f
C5786 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n9 GND 0.50079f
C5787 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n10 GND 0.64061f
C5788 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t15 GND 0.04476f
C5789 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t13 GND 0.07168f
C5790 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n11 GND 0.13717f
C5791 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n12 GND 0.47666f
C5792 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n13 GND 1.2109f
C5793 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t5 GND 0.07156f
C5794 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t9 GND 0.04466f
C5795 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n14 GND 0.1408f
C5796 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n15 GND 0.1064f
C5797 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n16 GND 0.7135f
C5798 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t7 GND 0.04466f
C5799 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t11 GND 0.07156f
C5800 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n17 GND 0.14228f
C5801 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t12 GND 0.04474f
C5802 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t16 GND 0.07165f
C5803 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n18 GND 0.1364f
C5804 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n19 GND 0.01603f
C5805 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n20 GND 0.16255f
C5806 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n21 GND 12.0678f
C5807 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n22 GND 8.45355f
C5808 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t1 GND 0.02814f
C5809 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t0 GND 0.02814f
C5810 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n23 GND 0.06709f
C5811 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n24 GND 0.1318f
C5812 VOUT.t84 GND 0.39129f
C5813 VOUT.n0 GND 0.37934f
C5814 VOUT.t80 GND 0.39174f
C5815 VOUT.n1 GND 0.3107f
C5816 VOUT.t56 GND 0.39129f
C5817 VOUT.n2 GND 0.24966f
C5818 VOUT.t72 GND 0.39174f
C5819 VOUT.n3 GND 0.3107f
C5820 VOUT.t85 GND 0.39129f
C5821 VOUT.n4 GND 0.24966f
C5822 VOUT.t52 GND 0.39129f
C5823 VOUT.n5 GND 0.47225f
C5824 VOUT.t67 GND 0.39174f
C5825 VOUT.n6 GND 0.5248f
C5826 VOUT.t76 GND 0.39174f
C5827 VOUT.n7 GND 0.3107f
C5828 VOUT.t61 GND 0.39174f
C5829 VOUT.n8 GND 0.27188f
C5830 VOUT.n9 GND 0.28449f
C5831 VOUT.n10 GND 0.34339f
C5832 VOUT.t79 GND 0.39129f
C5833 VOUT.n11 GND 0.21084f
C5834 VOUT.t70 GND 0.39129f
C5835 VOUT.n12 GND 0.24966f
C5836 VOUT.t71 GND 0.39129f
C5837 VOUT.n13 GND 0.21084f
C5838 VOUT.n14 GND 0.34339f
C5839 VOUT.n15 GND 0.28449f
C5840 VOUT.t63 GND 0.39174f
C5841 VOUT.n16 GND 0.27188f
C5842 VOUT.t57 GND 0.39174f
C5843 VOUT.n17 GND 0.3107f
C5844 VOUT.t59 GND 0.39174f
C5845 VOUT.n18 GND 0.27188f
C5846 VOUT.n19 GND 0.28449f
C5847 VOUT.n20 GND 0.34339f
C5848 VOUT.t86 GND 0.39129f
C5849 VOUT.n21 GND 0.21084f
C5850 VOUT.t51 GND 0.39129f
C5851 VOUT.n22 GND 0.24966f
C5852 VOUT.t83 GND 0.39129f
C5853 VOUT.n23 GND 0.21084f
C5854 VOUT.n24 GND 0.34339f
C5855 VOUT.n25 GND 0.28449f
C5856 VOUT.t54 GND 0.39174f
C5857 VOUT.n26 GND 0.27188f
C5858 VOUT.t69 GND 0.39174f
C5859 VOUT.n27 GND 0.30048f
C5860 VOUT.t38 GND 0.03027f
C5861 VOUT.t41 GND 0.03027f
C5862 VOUT.n28 GND 0.06343f
C5863 VOUT.t40 GND 0.03027f
C5864 VOUT.t39 GND 0.03027f
C5865 VOUT.n29 GND 0.06344f
C5866 VOUT.n30 GND 0.42057f
C5867 VOUT.t45 GND 0.01009f
C5868 VOUT.t44 GND 0.01009f
C5869 VOUT.n31 GND 0.02218f
C5870 VOUT.t47 GND 0.01009f
C5871 VOUT.t46 GND 0.01009f
C5872 VOUT.n32 GND 0.02218f
C5873 VOUT.n33 GND 0.14451f
C5874 VOUT.t17 GND 1.332f
C5875 VOUT.t4 GND 1.25774f
C5876 VOUT.n34 GND 0.42547f
C5877 VOUT.t43 GND 1.25774f
C5878 VOUT.n35 GND 0.21179f
C5879 VOUT.t16 GND 1.29039f
C5880 VOUT.n36 GND 0.2788f
C5881 VOUT.t11 GND 1.332f
C5882 VOUT.t6 GND 1.25774f
C5883 VOUT.n37 GND 0.42547f
C5884 VOUT.t2 GND 1.25774f
C5885 VOUT.n38 GND 0.21179f
C5886 VOUT.t9 GND 1.29039f
C5887 VOUT.n39 GND 0.25529f
C5888 VOUT.n40 GND 0.49984f
C5889 VOUT.t3 GND 1.332f
C5890 VOUT.t10 GND 1.25774f
C5891 VOUT.n41 GND 0.42547f
C5892 VOUT.t5 GND 1.25774f
C5893 VOUT.n42 GND 0.21179f
C5894 VOUT.t1 GND 1.29039f
C5895 VOUT.n43 GND 0.25529f
C5896 VOUT.n44 GND 0.33799f
C5897 VOUT.t0 GND 1.332f
C5898 VOUT.t15 GND 1.25774f
C5899 VOUT.n45 GND 0.42547f
C5900 VOUT.t13 GND 1.25774f
C5901 VOUT.n46 GND 0.21179f
C5902 VOUT.t42 GND 1.29039f
C5903 VOUT.n47 GND 0.25529f
C5904 VOUT.n48 GND 0.33799f
C5905 VOUT.t8 GND 1.332f
C5906 VOUT.t14 GND 1.25774f
C5907 VOUT.n49 GND 0.42547f
C5908 VOUT.t12 GND 1.25774f
C5909 VOUT.n50 GND 0.21179f
C5910 VOUT.t7 GND 1.29039f
C5911 VOUT.n51 GND 0.25529f
C5912 VOUT.n52 GND 0.50699f
C5913 VOUT.t19 GND 1.332f
C5914 VOUT.t32 GND 1.25774f
C5915 VOUT.n53 GND 0.42547f
C5916 VOUT.t26 GND 1.25774f
C5917 VOUT.n54 GND 0.21179f
C5918 VOUT.t20 GND 1.29039f
C5919 VOUT.n55 GND 0.25529f
C5920 VOUT.n56 GND 0.50699f
C5921 VOUT.t22 GND 1.332f
C5922 VOUT.t35 GND 1.25774f
C5923 VOUT.n57 GND 0.42547f
C5924 VOUT.t28 GND 1.25774f
C5925 VOUT.n58 GND 0.21179f
C5926 VOUT.t23 GND 1.29039f
C5927 VOUT.n59 GND 0.25529f
C5928 VOUT.n60 GND 0.33799f
C5929 VOUT.t30 GND 1.332f
C5930 VOUT.t25 GND 1.25774f
C5931 VOUT.n61 GND 0.42547f
C5932 VOUT.t18 GND 1.25774f
C5933 VOUT.n62 GND 0.21179f
C5934 VOUT.t31 GND 1.29039f
C5935 VOUT.n63 GND 0.25529f
C5936 VOUT.n64 GND 0.33799f
C5937 VOUT.t33 GND 1.332f
C5938 VOUT.t27 GND 1.25774f
C5939 VOUT.n65 GND 0.42547f
C5940 VOUT.t21 GND 1.25774f
C5941 VOUT.n66 GND 0.21179f
C5942 VOUT.t34 GND 1.29039f
C5943 VOUT.n67 GND 0.25529f
C5944 VOUT.n68 GND 0.33799f
C5945 VOUT.t36 GND 1.332f
C5946 VOUT.t29 GND 1.25774f
C5947 VOUT.n69 GND 0.42547f
C5948 VOUT.t24 GND 1.25774f
C5949 VOUT.n70 GND 0.21179f
C5950 VOUT.t37 GND 1.29039f
C5951 VOUT.n71 GND 0.25529f
C5952 VOUT.n72 GND 2.66762f
C5953 VOUT.n73 GND 1.16766f
C5954 VOUT.n74 GND 0.21357f
C5955 VOUT.n75 GND 0.70548f
C5956 VOUT.n76 GND 0.36499f
C5957 VOUT.n77 GND 0.34615f
C5958 VOUT.t64 GND 0.16094f
C5959 VOUT.n78 GND 0.3246f
C5960 VOUT.t87 GND 0.16028f
C5961 VOUT.n79 GND 0.19562f
C5962 VOUT.t53 GND 0.16094f
C5963 VOUT.n80 GND 0.25741f
C5964 VOUT.t65 GND 0.16028f
C5965 VOUT.n81 GND 0.19562f
C5966 VOUT.t73 GND 0.16094f
C5967 VOUT.n82 GND 0.25741f
C5968 VOUT.t62 GND 0.16094f
C5969 VOUT.n83 GND 0.38517f
C5970 VOUT.t48 GND 0.16028f
C5971 VOUT.n84 GND 0.3342f
C5972 VOUT.t81 GND 0.16028f
C5973 VOUT.n85 GND 0.19562f
C5974 VOUT.t74 GND 0.16028f
C5975 VOUT.n86 GND 0.15679f
C5976 VOUT.n87 GND 0.25717f
C5977 VOUT.n88 GND 0.20039f
C5978 VOUT.t58 GND 0.16094f
C5979 VOUT.n89 GND 0.21858f
C5980 VOUT.t68 GND 0.16094f
C5981 VOUT.n90 GND 0.25741f
C5982 VOUT.t60 GND 0.16094f
C5983 VOUT.n91 GND 0.21858f
C5984 VOUT.n92 GND 0.20039f
C5985 VOUT.n93 GND 0.25717f
C5986 VOUT.t66 GND 0.16028f
C5987 VOUT.n94 GND 0.15679f
C5988 VOUT.t50 GND 0.16028f
C5989 VOUT.n95 GND 0.19562f
C5990 VOUT.t82 GND 0.16028f
C5991 VOUT.n96 GND 0.15679f
C5992 VOUT.n97 GND 0.25717f
C5993 VOUT.n98 GND 0.20039f
C5994 VOUT.t55 GND 0.16094f
C5995 VOUT.n99 GND 0.21858f
C5996 VOUT.t75 GND 0.16094f
C5997 VOUT.n100 GND 0.25741f
C5998 VOUT.t49 GND 0.16094f
C5999 VOUT.n101 GND 0.21858f
C6000 VOUT.n102 GND 0.20039f
C6001 VOUT.n103 GND 0.25717f
C6002 VOUT.t77 GND 0.16028f
C6003 VOUT.n104 GND 0.15679f
C6004 VOUT.t78 GND 0.16028f
C6005 VOUT.n105 GND 0.25303f
C6006 VOUT.n106 GND 0.23589f
C6007 a_14948_18696.t1 GND 0.06282f
C6008 a_14948_18696.t2 GND 0.0622f
C6009 a_14948_18696.n0 GND 4.49915f
C6010 a_14948_18696.t0 GND 0.07583f
C6011 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t0 GND 0.09531f
C6012 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n0 GND 0.03908f
C6013 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n1 GND 0.08412f
C6014 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n2 GND 0.05585f
C6015 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t1 GND 0.09131f
C6016 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n3 GND 0.01153f
C6017 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t3 GND 0.18843f
C6018 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n4 GND 0.22732f
C6019 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t5 GND 0.18933f
C6020 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t2 GND 0.18843f
C6021 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n5 GND 0.59073f
C6022 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t4 GND 0.18843f
C6023 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n6 GND 0.29581f
C6024 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n7 GND 0.19692f
C6025 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t7 GND 0.18633f
C6026 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n8 GND 13.978f
C6027 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t6 GND 0.33331f
C6028 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].t8 GND 0.1849f
C6029 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n9 GND 0.29045f
C6030 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n10 GND 0.05778f
C6031 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5].n11 GND 0.08285f
C6032 a_23307_20174.t2 GND 0.12979f
C6033 a_23307_20174.t1 GND 0.07321f
C6034 a_23307_20174.n0 GND 4.33997f
C6035 a_23307_20174.t3 GND 0.1514f
C6036 a_23307_20174.t4 GND 0.06185f
C6037 a_23307_20174.n1 GND 4.46413f
C6038 a_23307_20174.n2 GND 1.20642f
C6039 a_23307_20174.t0 GND 0.07321f
C6040 a_22193_18133.t1 GND 0.04073f
C6041 a_22193_18133.t4 GND 0.04729f
C6042 a_22193_18133.t2 GND 0.0337f
C6043 a_22193_18133.n0 GND 1.6865f
C6044 a_22193_18133.t3 GND 0.0337f
C6045 a_22193_18133.n1 GND 0.82505f
C6046 a_22193_18133.n2 GND 1.39933f
C6047 a_22193_18133.t0 GND 0.0337f
C6048 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t6 GND 0.17284f
C6049 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t3 GND 0.17234f
C6050 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n0 GND 0.21906f
C6051 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t2 GND 0.17321f
C6052 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t4 GND 0.17234f
C6053 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n1 GND 0.56133f
C6054 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n2 GND 0.18922f
C6055 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t7 GND 0.17035f
C6056 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n3 GND 16.4341f
C6057 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t0 GND 0.1425f
C6058 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t1 GND 0.12117f
C6059 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n4 GND 0.97482f
C6060 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t8 GND 0.56576f
C6061 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t9 GND 0.56342f
C6062 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n5 GND 0.89432f
C6063 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n6 GND 0.57694f
C6064 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].t5 GND 0.595f
C6065 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1].n7 GND 1.24415f
C6066 a_19946_8950.t2 GND 0.07897f
C6067 a_19946_8950.t1 GND 0.06395f
C6068 a_19946_8950.n0 GND 5.77629f
C6069 a_19946_8950.t0 GND 0.08079f
C6070 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t0 GND 0.08787f
C6071 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n0 GND 0.03603f
C6072 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n1 GND 0.07755f
C6073 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n2 GND 0.05149f
C6074 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t1 GND 0.08418f
C6075 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n3 GND 0.01063f
C6076 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t3 GND 0.16833f
C6077 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t13 GND 0.17389f
C6078 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n4 GND 0.67814f
C6079 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t10 GND 0.17455f
C6080 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t6 GND 0.17372f
C6081 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n5 GND 0.54462f
C6082 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t8 GND 0.17372f
C6083 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n6 GND 0.22043f
C6084 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n7 GND 0.18155f
C6085 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t2 GND 0.17179f
C6086 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n8 GND 1.83198f
C6087 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n9 GND 8.61447f
C6088 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t12 GND 0.16619f
C6089 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t7 GND 0.16535f
C6090 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n10 GND 0.50865f
C6091 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t11 GND 0.16619f
C6092 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n11 GND 0.38958f
C6093 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t5 GND 0.16345f
C6094 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n12 GND 1.84501f
C6095 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n13 GND 9.22158f
C6096 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t9 GND 0.3073f
C6097 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.t4 GND 0.17047f
C6098 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n14 GND 0.26778f
C6099 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n15 GND 0.05327f
C6100 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2.n16 GND 0.07638f
C6101 top_DAC_0/top_rseg_n_dcell_0.VH2.t7 GND 0.02406f
C6102 top_DAC_0/top_rseg_n_dcell_0.VH2.t3 GND 0.02383f
C6103 top_DAC_0/top_rseg_n_dcell_0.VH2.t4 GND 0.03364f
C6104 top_DAC_0/top_rseg_n_dcell_0.VH2.n0 GND 0.53585f
C6105 top_DAC_0/top_rseg_n_dcell_0.VH2.t6 GND 0.02756f
C6106 top_DAC_0/top_rseg_n_dcell_0.VH2.n1 GND 0.4485f
C6107 top_DAC_0/top_rseg_n_dcell_0.VH2.n2 GND 0.01342f
C6108 top_DAC_0/top_rseg_n_dcell_0.VH2.n3 GND 1.85868f
C6109 top_DAC_0/top_rseg_n_dcell_0.VH2.t2 GND 0.02378f
C6110 top_DAC_0/top_rseg_n_dcell_0.VH2.t5 GND 0.0236f
C6111 top_DAC_0/top_rseg_n_dcell_0.VH2.n4 GND 0.15084f
C6112 top_DAC_0/top_rseg_n_dcell_0.VH2.t0 GND 0.0236f
C6113 top_DAC_0/top_rseg_n_dcell_0.VH2.n5 GND 0.08573f
C6114 top_DAC_0/top_rseg_n_dcell_0.VH2.t1 GND 0.0236f
C6115 top_DAC_0/top_rseg_n_dcell_0.VH2.n6 GND 0.12889f
C6116 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y GND 0.63154f
C6117 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t0 GND 0.1039f
C6118 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n0 GND 0.0426f
C6119 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n1 GND 0.09171f
C6120 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n2 GND 0.06089f
C6121 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t1 GND 0.09954f
C6122 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n3 GND 0.01257f
C6123 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t2 GND 0.204f
C6124 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t5 GND 0.20641f
C6125 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n4 GND 0.98607f
C6126 top_DAC_0/top_final_switch_0.b[0] GND 1.14816f
C6127 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t4 GND 0.29113f
C6128 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n5 GND 10.7165f
C6129 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.b[0] GND 0.20833f
C6130 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.t3 GND 0.19328f
C6131 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n6 GND 2.03795f
C6132 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n7 GND 12.8056f
C6133 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.b[0] GND 3.73787f
C6134 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUT GND 0.35647f
C6135 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0.n8 GND 0.06555f
C6136 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t3 GND 0.04249f
C6137 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t2 GND 0.04249f
C6138 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 GND 0.09332f
C6139 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y GND 0.21353f
C6140 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 GND 0.04026f
C6141 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t4 GND 0.72401f
C6142 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 GND 15.9934f
C6143 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t1 GND 0.02762f
C6144 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t0 GND 0.02762f
C6145 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 GND 0.06586f
C6146 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 GND 0.12938f
C6147 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t1 GND 0.02634f
C6148 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t2 GND 0.02634f
C6149 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 GND 0.06281f
C6150 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y GND 0.20365f
C6151 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 GND 0.1234f
C6152 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t5 GND 0.06304f
C6153 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t7 GND 0.03715f
C6154 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t4 GND 0.06304f
C6155 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t6 GND 0.03715f
C6156 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 GND 0.10577f
C6157 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 GND 0.15692f
C6158 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.A GND 0.01051f
C6159 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 GND 0.04732f
C6160 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t8 GND 0.51546f
C6161 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 GND 15.6837f
C6162 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 GND 0.02899f
C6163 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 GND 0.03839f
C6164 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t3 GND 0.04053f
C6165 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t0 GND 0.04053f
C6166 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 GND 0.089f
C6167 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t2 GND 0.01247f
C6168 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t1 GND 0.08855f
C6169 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t0 GND 0.09059f
C6170 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.n0 GND 1.58122f
C6171 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t2 GND 0.04184f
C6172 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t3 GND 0.04184f
C6173 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 GND 0.09189f
C6174 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y GND 0.21025f
C6175 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 GND 0.03964f
C6176 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t20 GND 0.06508f
C6177 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t9 GND 0.03835f
C6178 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t12 GND 0.06508f
C6179 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t4 GND 0.03835f
C6180 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 GND 0.1092f
C6181 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 GND 0.162f
C6182 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.A GND 0.01085f
C6183 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 GND 0.04886f
C6184 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t13 GND 0.06917f
C6185 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t6 GND 0.04317f
C6186 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 GND 0.13623f
C6187 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.B GND 0.01674f
C6188 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 GND 0.06232f
C6189 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t16 GND 0.06917f
C6190 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t8 GND 0.04317f
C6191 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 GND 0.13618f
C6192 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.B GND 0.01715f
C6193 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 GND 0.046f
C6194 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 GND 0.71314f
C6195 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[0] GND 1.82836f
C6196 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t15 GND 0.25867f
C6197 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 GND 5.84879f
C6198 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x1.B GND 0.01799f
C6199 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t5 GND 0.04317f
C6200 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t19 GND 0.06917f
C6201 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 GND 0.13609f
C6202 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 GND 0.12915f
C6203 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[6] GND 0.18f
C6204 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 GND 0.89598f
C6205 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t11 GND 0.07051f
C6206 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t17 GND 0.04428f
C6207 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 GND 0.09547f
C6208 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x2.C GND -0.02483f
C6209 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 GND 0.41728f
C6210 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 GND 1.14727f
C6211 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.A GND 0.01994f
C6212 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t18 GND 0.04344f
C6213 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t14 GND 0.06949f
C6214 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 GND 0.12217f
C6215 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 GND 0.19259f
C6216 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 GND 1.11131f
C6217 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t7 GND 0.04344f
C6218 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t10 GND 0.06949f
C6219 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 GND 0.12266f
C6220 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.A GND 0.01585f
C6221 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 GND 0.13712f
C6222 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 GND 5.41443f
C6223 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 GND 8.07493f
C6224 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 GND 1.01356f
C6225 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 GND 0.02993f
C6226 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t0 GND 0.0272f
C6227 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t1 GND 0.0272f
C6228 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 GND 0.06485f
C6229 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 GND 0.1274f
C6230 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t0 GND 0.22296f
C6231 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t18 GND 0.22296f
C6232 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t6 GND 0.22296f
C6233 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n0 GND 1.07167f
C6234 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t8 GND 0.22296f
C6235 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t7 GND 0.22296f
C6236 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n1 GND 0.84762f
C6237 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n2 GND 1.36355f
C6238 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t14 GND 0.22296f
C6239 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t13 GND 0.22296f
C6240 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n3 GND 0.84762f
C6241 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n4 GND 0.58565f
C6242 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t35 GND 0.2513f
C6243 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t23 GND 0.24374f
C6244 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n5 GND 1.86562f
C6245 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t24 GND 0.24374f
C6246 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n6 GND 1.07339f
C6247 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t20 GND 0.24374f
C6248 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n7 GND 0.98889f
C6249 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t36 GND 0.2513f
C6250 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t33 GND 0.24374f
C6251 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n8 GND 1.86562f
C6252 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t34 GND 0.24374f
C6253 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n9 GND 1.07339f
C6254 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t21 GND 0.24374f
C6255 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n10 GND 1.07339f
C6256 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t28 GND 0.24374f
C6257 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n11 GND 1.07339f
C6258 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t22 GND 0.24374f
C6259 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n12 GND 0.85936f
C6260 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n13 GND 0.79614f
C6261 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t31 GND 0.2513f
C6262 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t32 GND 0.24374f
C6263 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n14 GND 1.86562f
C6264 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t26 GND 0.24374f
C6265 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n15 GND 1.07339f
C6266 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t27 GND 0.24374f
C6267 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n16 GND 1.07339f
C6268 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t38 GND 0.24374f
C6269 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n17 GND 1.02698f
C6270 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t30 GND 0.2513f
C6271 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t37 GND 0.24374f
C6272 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n18 GND 1.86562f
C6273 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t29 GND 0.24374f
C6274 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n19 GND 1.07339f
C6275 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t25 GND 0.24374f
C6276 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n20 GND 1.07339f
C6277 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t39 GND 0.24374f
C6278 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n21 GND 0.89746f
C6279 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n22 GND 0.22235f
C6280 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n23 GND 2.09603f
C6281 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t3 GND 0.22296f
C6282 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t11 GND 0.22296f
C6283 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n24 GND 1.07167f
C6284 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t10 GND 0.22296f
C6285 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t17 GND 0.22296f
C6286 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n25 GND 0.84762f
C6287 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n26 GND 1.16787f
C6288 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t5 GND 0.22296f
C6289 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t9 GND 0.22296f
C6290 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n27 GND 1.07167f
C6291 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t16 GND 0.22296f
C6292 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t4 GND 0.22296f
C6293 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n28 GND 0.84762f
C6294 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n29 GND 1.36355f
C6295 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t12 GND 0.22296f
C6296 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t2 GND 0.22296f
C6297 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n30 GND 0.84762f
C6298 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n31 GND 0.71657f
C6299 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n32 GND 0.52089f
C6300 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n33 GND 1.30443f
C6301 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n34 GND 0.70528f
C6302 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t15 GND 0.22296f
C6303 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t1 GND 0.22296f
C6304 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n35 GND 0.84762f
C6305 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n36 GND 1.29878f
C6306 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n37 GND 1.07167f
C6307 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t19 GND 0.22296f
C6308 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t2 GND 0.04693f
C6309 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t3 GND 0.04693f
C6310 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n0 GND 0.10307f
C6311 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n1 GND 0.04446f
C6312 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t11 GND 0.073f
C6313 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t16 GND 0.04302f
C6314 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t8 GND 0.073f
C6315 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t14 GND 0.04302f
C6316 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n2 GND 0.12249f
C6317 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n3 GND 0.18172f
C6318 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n4 GND 0.0548f
C6319 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t15 GND 0.07759f
C6320 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t7 GND 0.04842f
C6321 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n5 GND 0.15426f
C6322 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t9 GND 0.07769f
C6323 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t19 GND 0.04851f
C6324 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n6 GND 0.14788f
C6325 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n7 GND 0.04318f
C6326 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t4 GND 0.04851f
C6327 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t18 GND 0.07769f
C6328 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n8 GND 0.14809f
C6329 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n9 GND 0.25203f
C6330 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n10 GND 0.72876f
C6331 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t5 GND 0.07749f
C6332 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t12 GND 0.04834f
C6333 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n11 GND 0.1591f
C6334 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n12 GND 1.10696f
C6335 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t17 GND 0.04966f
C6336 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t13 GND 0.07909f
C6337 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n13 GND 0.10732f
C6338 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n14 GND 1.43878f
C6339 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t6 GND 0.04966f
C6340 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t10 GND 0.07909f
C6341 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n15 GND 0.10732f
C6342 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n16 GND 5.7562f
C6343 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n17 GND 11.8589f
C6344 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n18 GND 1.22867f
C6345 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n19 GND 0.03358f
C6346 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t0 GND 0.0305f
C6347 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t1 GND 0.0305f
C6348 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n20 GND 0.07274f
C6349 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n21 GND 0.1429f
C6350 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t4 GND 0.18931f
C6351 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t1 GND 0.18936f
C6352 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t3 GND 0.18936f
C6353 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n0 GND 0.86568f
C6354 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t2 GND 0.18936f
C6355 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t5 GND 0.18936f
C6356 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n1 GND 0.95127f
C6357 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t6 GND 0.18931f
C6358 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t0 GND 0.18931f
C6359 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n2 GND 0.73533f
C6360 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n3 GND 1.158f
C6361 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t11 GND 0.21344f
C6362 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t12 GND 0.20701f
C6363 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n4 GND 1.77158f
C6364 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t8 GND 0.21344f
C6365 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t10 GND 0.20701f
C6366 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n5 GND 1.36507f
C6367 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n6 GND 0.47809f
C6368 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t13 GND 0.21344f
C6369 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t15 GND 0.20701f
C6370 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n7 GND 1.55038f
C6371 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t14 GND 0.21344f
C6372 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t9 GND 0.20701f
C6373 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n8 GND 1.58627f
C6374 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n9 GND 0.47475f
C6375 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n10 GND 0.91364f
C6376 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n11 GND 1.20528f
C6377 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n12 GND 1.09031f
C6378 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n13 GND 0.85788f
C6379 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t7 GND 0.18931f
C6380 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t2 GND 0.05236f
C6381 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t7 GND 0.04377f
C6382 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t4 GND 0.02732f
C6383 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n0 GND 0.08703f
C6384 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t5 GND 0.04383f
C6385 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t9 GND 0.02737f
C6386 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n1 GND 0.08343f
C6387 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n2 GND 0.01642f
C6388 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n3 GND 0.0358f
C6389 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n4 GND 5.85791f
C6390 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t6 GND 0.04386f
C6391 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t8 GND 0.02739f
C6392 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n5 GND 0.0822f
C6393 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n6 GND 0.02224f
C6394 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n7 GND 0.2998f
C6395 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n8 GND 0.13919f
C6396 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t1 GND 0.02648f
C6397 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t3 GND 0.02648f
C6398 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n9 GND 0.05886f
C6399 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t0 GND 0.12167f
C6400 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n10 GND 0.29364f
C6401 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t3 GND 0.04411f
C6402 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t2 GND 0.04411f
C6403 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 GND 0.09687f
C6404 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y GND 0.22166f
C6405 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 GND 0.04179f
C6406 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t4 GND 0.73789f
C6407 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 GND 16.6536f
C6408 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t1 GND 0.02867f
C6409 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t0 GND 0.02867f
C6410 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 GND 0.06836f
C6411 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 GND 0.1343f
C6412 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t2 GND 0.02769f
C6413 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t3 GND 0.02769f
C6414 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 GND 0.06602f
C6415 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y GND 0.21405f
C6416 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 GND 0.1297f
C6417 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t7 GND 0.06626f
C6418 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t5 GND 0.03905f
C6419 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t6 GND 0.06626f
C6420 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t4 GND 0.03905f
C6421 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 GND 0.11117f
C6422 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 GND 0.16493f
C6423 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.A GND 0.01104f
C6424 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 GND 0.04974f
C6425 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t8 GND 0.51398f
C6426 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 GND 16.3238f
C6427 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 GND 0.03047f
C6428 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 GND 0.04035f
C6429 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t0 GND 0.04259f
C6430 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t1 GND 0.04259f
C6431 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 GND 0.09355f
C6432 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t7 GND 0.23722f
C6433 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t9 GND 0.23722f
C6434 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t14 GND 0.23722f
C6435 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n0 GND 1.14024f
C6436 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t1 GND 0.23722f
C6437 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t8 GND 0.23722f
C6438 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n1 GND 0.90185f
C6439 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n2 GND 1.45079f
C6440 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t0 GND 0.23722f
C6441 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t6 GND 0.23722f
C6442 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n3 GND 0.90185f
C6443 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n4 GND 0.80884f
C6444 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t25 GND 0.26404f
C6445 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t21 GND 0.25657f
C6446 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n5 GND 1.86139f
C6447 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t32 GND 0.25657f
C6448 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n6 GND 1.07998f
C6449 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t20 GND 0.25657f
C6450 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n7 GND 1.07998f
C6451 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t34 GND 0.25657f
C6452 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n8 GND 0.98418f
C6453 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t24 GND 0.26404f
C6454 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t23 GND 0.25657f
C6455 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n9 GND 1.86139f
C6456 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t22 GND 0.25657f
C6457 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n10 GND 1.07998f
C6458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t39 GND 0.25657f
C6459 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n11 GND 1.07998f
C6460 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t29 GND 0.25657f
C6461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n12 GND 0.93922f
C6462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n13 GND 0.71895f
C6463 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t28 GND 0.26404f
C6464 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t37 GND 0.25657f
C6465 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n14 GND 1.86139f
C6466 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t31 GND 0.25657f
C6467 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n15 GND 1.07998f
C6468 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t30 GND 0.25657f
C6469 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n16 GND 0.94364f
C6470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t35 GND 0.26404f
C6471 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t26 GND 0.25657f
C6472 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n17 GND 1.86139f
C6473 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t27 GND 0.25657f
C6474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n18 GND 1.07998f
C6475 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t33 GND 0.25657f
C6476 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n19 GND 1.07998f
C6477 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t38 GND 0.25657f
C6478 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n20 GND 1.07998f
C6479 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t36 GND 0.25657f
C6480 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n21 GND 0.89869f
C6481 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n22 GND 0.31764f
C6482 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n23 GND 2.2018f
C6483 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t10 GND 0.23722f
C6484 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t15 GND 0.23722f
C6485 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n24 GND 1.14024f
C6486 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t17 GND 0.23722f
C6487 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t16 GND 0.23722f
C6488 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n25 GND 0.90185f
C6489 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n26 GND 1.45079f
C6490 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t4 GND 0.23722f
C6491 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t3 GND 0.23722f
C6492 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n27 GND 0.90185f
C6493 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n28 GND 0.57669f
C6494 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t12 GND 0.23722f
C6495 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t11 GND 0.23722f
C6496 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n29 GND 1.14024f
C6497 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t5 GND 0.23722f
C6498 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t13 GND 0.23722f
C6499 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n30 GND 0.90185f
C6500 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n31 GND 1.42831f
C6501 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n32 GND 0.55421f
C6502 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n33 GND 1.34907f
C6503 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n34 GND 0.71788f
C6504 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t18 GND 0.23722f
C6505 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t2 GND 0.23722f
C6506 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n35 GND 0.90185f
C6507 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n36 GND 1.19616f
C6508 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n37 GND 1.14024f
C6509 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t19 GND 0.23722f
C6510 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t17 GND 0.1404f
C6511 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t21 GND 0.3674f
C6512 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n0 GND 4.05473f
C6513 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t15 GND 0.13993f
C6514 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t3 GND 0.13993f
C6515 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n1 GND 0.57903f
C6516 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n2 GND 1.11378f
C6517 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t18 GND 0.13993f
C6518 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t10 GND 0.13993f
C6519 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n3 GND 0.71886f
C6520 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t5 GND 0.13993f
C6521 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t9 GND 0.13993f
C6522 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n4 GND 0.57903f
C6523 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n5 GND 0.86298f
C6524 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t19 GND 0.13993f
C6525 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t20 GND 0.13993f
C6526 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n6 GND 0.57903f
C6527 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n7 GND 0.37161f
C6528 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t25 GND 0.53665f
C6529 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t89 GND 0.5347f
C6530 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n8 GND 0.70644f
C6531 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t66 GND 0.5347f
C6532 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n9 GND 0.35419f
C6533 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t22 GND 0.5347f
C6534 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n10 GND 0.35419f
C6535 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t80 GND 0.5347f
C6536 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n11 GND 0.35419f
C6537 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t81 GND 0.5347f
C6538 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n12 GND 0.35419f
C6539 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t30 GND 0.5347f
C6540 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n13 GND 0.35419f
C6541 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t82 GND 0.5347f
C6542 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n14 GND 0.35354f
C6543 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t43 GND 0.53665f
C6544 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t64 GND 0.5347f
C6545 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n15 GND 0.70644f
C6546 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t24 GND 0.5347f
C6547 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n16 GND 0.35419f
C6548 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t101 GND 0.5347f
C6549 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n17 GND 0.35419f
C6550 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t65 GND 0.5347f
C6551 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n18 GND 0.35419f
C6552 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t87 GND 0.5347f
C6553 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n19 GND 0.35419f
C6554 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t98 GND 0.5347f
C6555 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n20 GND 0.35419f
C6556 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t42 GND 0.5347f
C6557 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n21 GND 0.35419f
C6558 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t70 GND 0.5347f
C6559 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n22 GND 0.35419f
C6560 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t99 GND 0.5347f
C6561 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n23 GND 0.35419f
C6562 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t50 GND 0.5347f
C6563 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n24 GND 0.35419f
C6564 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t46 GND 0.5347f
C6565 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n25 GND 0.2731f
C6566 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n26 GND 0.12073f
C6567 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t36 GND 0.53665f
C6568 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t96 GND 0.5347f
C6569 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n27 GND 0.70644f
C6570 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t71 GND 0.5347f
C6571 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n28 GND 0.35419f
C6572 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t33 GND 0.5347f
C6573 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n29 GND 0.35419f
C6574 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t85 GND 0.5347f
C6575 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n30 GND 0.35419f
C6576 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t88 GND 0.5347f
C6577 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n31 GND 0.35419f
C6578 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t39 GND 0.5347f
C6579 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n32 GND 0.35419f
C6580 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t90 GND 0.5347f
C6581 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n33 GND 0.35354f
C6582 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t49 GND 0.53665f
C6583 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t67 GND 0.5347f
C6584 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n34 GND 0.70644f
C6585 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t34 GND 0.5347f
C6586 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n35 GND 0.35419f
C6587 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t29 GND 0.5347f
C6588 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n36 GND 0.35419f
C6589 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t69 GND 0.5347f
C6590 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n37 GND 0.35419f
C6591 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t94 GND 0.5347f
C6592 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n38 GND 0.35419f
C6593 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t26 GND 0.5347f
C6594 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n39 GND 0.35419f
C6595 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t44 GND 0.5347f
C6596 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n40 GND 0.35419f
C6597 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t75 GND 0.5347f
C6598 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n41 GND 0.35419f
C6599 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t28 GND 0.5347f
C6600 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n42 GND 0.35419f
C6601 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t59 GND 0.5347f
C6602 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n43 GND 0.35419f
C6603 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t54 GND 0.5347f
C6604 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n44 GND 0.2731f
C6605 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n45 GND 0.08175f
C6606 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n46 GND 0.46995f
C6607 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t53 GND 0.53665f
C6608 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t37 GND 0.5347f
C6609 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n47 GND 0.70644f
C6610 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t86 GND 0.5347f
C6611 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n48 GND 0.35419f
C6612 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t51 GND 0.5347f
C6613 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n49 GND 0.35419f
C6614 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t100 GND 0.5347f
C6615 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n50 GND 0.35419f
C6616 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t23 GND 0.5347f
C6617 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n51 GND 0.35419f
C6618 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t57 GND 0.5347f
C6619 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n52 GND 0.35419f
C6620 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t27 GND 0.5347f
C6621 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n53 GND 0.35354f
C6622 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t72 GND 0.53665f
C6623 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t83 GND 0.5347f
C6624 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n54 GND 0.70644f
C6625 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t52 GND 0.5347f
C6626 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n55 GND 0.35419f
C6627 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t48 GND 0.5347f
C6628 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n56 GND 0.35419f
C6629 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t84 GND 0.5347f
C6630 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n57 GND 0.35419f
C6631 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t32 GND 0.5347f
C6632 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n58 GND 0.35419f
C6633 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t45 GND 0.5347f
C6634 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n59 GND 0.35419f
C6635 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t68 GND 0.5347f
C6636 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n60 GND 0.35419f
C6637 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t93 GND 0.5347f
C6638 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n61 GND 0.35419f
C6639 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t47 GND 0.5347f
C6640 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n62 GND 0.35419f
C6641 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t76 GND 0.5347f
C6642 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n63 GND 0.35419f
C6643 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t74 GND 0.5347f
C6644 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n64 GND 0.2731f
C6645 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n65 GND 0.08175f
C6646 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n66 GND 0.26882f
C6647 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t62 GND 0.53665f
C6648 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t41 GND 0.5347f
C6649 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n67 GND 0.70644f
C6650 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t95 GND 0.5347f
C6651 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n68 GND 0.35419f
C6652 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t60 GND 0.5347f
C6653 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n69 GND 0.35419f
C6654 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t31 GND 0.5347f
C6655 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n70 GND 0.35419f
C6656 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t35 GND 0.5347f
C6657 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n71 GND 0.35419f
C6658 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t63 GND 0.5347f
C6659 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n72 GND 0.35419f
C6660 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t38 GND 0.5347f
C6661 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n73 GND 0.35354f
C6662 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t77 GND 0.53665f
C6663 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t91 GND 0.5347f
C6664 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n74 GND 0.70644f
C6665 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t61 GND 0.5347f
C6666 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n75 GND 0.35419f
C6667 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t58 GND 0.5347f
C6668 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n76 GND 0.35419f
C6669 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t92 GND 0.5347f
C6670 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n77 GND 0.35419f
C6671 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t40 GND 0.5347f
C6672 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n78 GND 0.35419f
C6673 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t55 GND 0.5347f
C6674 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n79 GND 0.35419f
C6675 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t73 GND 0.5347f
C6676 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n80 GND 0.35419f
C6677 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t97 GND 0.5347f
C6678 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n81 GND 0.35419f
C6679 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t56 GND 0.5347f
C6680 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n82 GND 0.35419f
C6681 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t79 GND 0.5347f
C6682 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n83 GND 0.35419f
C6683 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t78 GND 0.5347f
C6684 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n84 GND 0.2731f
C6685 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n85 GND 0.08175f
C6686 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n86 GND 0.33195f
C6687 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t4 GND 0.13993f
C6688 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t0 GND 0.13993f
C6689 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n87 GND 0.57903f
C6690 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n88 GND 0.45206f
C6691 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t13 GND 0.13993f
C6692 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t16 GND 0.13993f
C6693 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n89 GND 0.71769f
C6694 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t1 GND 0.13993f
C6695 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t14 GND 0.13993f
C6696 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n90 GND 0.57903f
C6697 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n91 GND 0.86297f
C6698 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t2 GND 0.13993f
C6699 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t8 GND 0.13993f
C6700 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n92 GND 0.57903f
C6701 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n93 GND 0.53511f
C6702 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n94 GND 0.55982f
C6703 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n95 GND 1.16531f
C6704 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n96 GND 0.327f
C6705 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t6 GND 0.13993f
C6706 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t7 GND 0.13993f
C6707 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n97 GND 0.57903f
C6708 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n98 GND 0.61556f
C6709 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t11 GND 0.13993f
C6710 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t12 GND 0.13993f
C6711 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n99 GND 0.57787f
C6712 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n100 GND 0.72563f
C6713 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n101 GND 2.68137f
C6714 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n102 GND 0.36894f
C6715 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t3 GND 0.02431f
C6716 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t1 GND 0.02431f
C6717 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 GND 0.05796f
C6718 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y GND 0.18793f
C6719 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 GND 0.11387f
C6720 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.A GND 0.01066f
C6721 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t17 GND 0.0619f
C6722 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t11 GND 0.03865f
C6723 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 GND 0.11784f
C6724 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 GND 0.07161f
C6725 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.A GND 0.01066f
C6726 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t9 GND 0.0619f
C6727 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t16 GND 0.03865f
C6728 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 GND 0.11784f
C6729 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 GND 0.03158f
C6730 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 GND 0.64907f
C6731 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[0] GND 1.66982f
C6732 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t4 GND 0.23188f
C6733 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 GND 5.28977f
C6734 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[6] GND 0.11568f
C6735 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t13 GND 0.03865f
C6736 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t12 GND 0.0619f
C6737 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 GND 0.118f
C6738 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x2.A GND 0.0167f
C6739 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 GND 0.21334f
C6740 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 GND 0.62504f
C6741 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t15 GND 0.06302f
C6742 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t5 GND 0.03957f
C6743 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 GND 0.09737f
C6744 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x1.B GND 0.03102f
C6745 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 GND 0.34887f
C6746 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 GND 0.85432f
C6747 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t6 GND 0.03865f
C6748 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t18 GND 0.0619f
C6749 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 GND 0.11826f
C6750 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x3.A GND 0.01299f
C6751 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 GND 0.25368f
C6752 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 GND 0.89808f
C6753 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x2.A GND 0.01066f
C6754 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t8 GND 0.0619f
C6755 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t14 GND 0.03865f
C6756 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 GND 0.11784f
C6757 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 GND 0.1843f
C6758 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 GND 0.83617f
C6759 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t7 GND 0.03865f
C6760 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t10 GND 0.0619f
C6761 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 GND 0.11809f
C6762 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.A GND 0.0153f
C6763 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 GND 0.21398f
C6764 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 GND 4.36182f
C6765 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 GND 8.09385f
C6766 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 GND 0.43725f
C6767 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 GND 0.03543f
C6768 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t2 GND 0.0374f
C6769 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t0 GND 0.0374f
C6770 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n26 GND 0.08213f
C6771 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t3 GND 0.08659f
C6772 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t31 GND 0.08376f
C6773 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n0 GND 1.26472f
C6774 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t29 GND 0.08376f
C6775 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n1 GND 0.77891f
C6776 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t25 GND 0.08376f
C6777 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n2 GND 0.77891f
C6778 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t6 GND 0.08376f
C6779 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n3 GND 0.68725f
C6780 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t2 GND 0.08659f
C6781 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t28 GND 0.08376f
C6782 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n4 GND 1.26472f
C6783 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t26 GND 0.08376f
C6784 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n5 GND 0.63996f
C6785 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n6 GND 0.54086f
C6786 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t30 GND 0.08659f
C6787 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t24 GND 0.08376f
C6788 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n7 GND 1.26472f
C6789 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t7 GND 0.08376f
C6790 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n8 GND 0.77891f
C6791 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t0 GND 0.08376f
C6792 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n9 GND 0.64432f
C6793 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t4 GND 0.08659f
C6794 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t1 GND 0.08376f
C6795 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n10 GND 1.26472f
C6796 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t5 GND 0.08376f
C6797 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n11 GND 0.77891f
C6798 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t27 GND 0.08376f
C6799 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n12 GND 0.59704f
C6800 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n13 GND 0.31646f
C6801 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n14 GND 1.724f
C6802 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t20 GND 0.07878f
C6803 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t16 GND 0.07878f
C6804 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n15 GND 0.5907f
C6805 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t19 GND 0.07878f
C6806 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t13 GND 0.07878f
C6807 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n16 GND 0.35538f
C6808 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n17 GND 1.18222f
C6809 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t12 GND 0.07878f
C6810 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t11 GND 0.07878f
C6811 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n18 GND 0.5907f
C6812 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t17 GND 0.07878f
C6813 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t8 GND 0.07878f
C6814 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n19 GND 0.35538f
C6815 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n20 GND 1.13493f
C6816 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n21 GND 0.65639f
C6817 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t15 GND 0.07878f
C6818 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t14 GND 0.07878f
C6819 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n22 GND 0.5907f
C6820 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t18 GND 0.07878f
C6821 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t22 GND 0.07878f
C6822 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n23 GND 0.35538f
C6823 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n24 GND 1.43212f
C6824 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t9 GND 0.07878f
C6825 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t23 GND 0.07878f
C6826 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n25 GND 0.35538f
C6827 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n26 GND 0.57073f
C6828 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t10 GND 0.07878f
C6829 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t21 GND 0.07878f
C6830 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n27 GND 0.57514f
C6831 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n28 GND 0.87695f
C6832 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n29 GND 1.05186f
C6833 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t0 GND 0.03763f
C6834 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t18 GND 0.03763f
C6835 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n0 GND 0.55219f
C6836 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t20 GND 0.03762f
C6837 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t7 GND 0.03758f
C6838 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n1 GND 0.26539f
C6839 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t3 GND 0.03758f
C6840 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n2 GND 0.29049f
C6841 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t6 GND 0.03763f
C6842 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n3 GND 0.35844f
C6843 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n4 GND 0.43211f
C6844 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t13 GND 0.03758f
C6845 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t21 GND 0.03758f
C6846 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n5 GND 0.19468f
C6847 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n6 GND 0.19468f
C6848 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n7 GND 0.27467f
C6849 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n8 GND 0.27467f
C6850 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t16 GND 0.03758f
C6851 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t12 GND 0.03758f
C6852 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n9 GND 0.19468f
C6853 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n10 GND 0.19468f
C6854 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n11 GND 0.03513f
C6855 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n12 GND 0.60467f
C6856 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t5 GND 0.03758f
C6857 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t14 GND 0.03762f
C6858 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t17 GND 0.03758f
C6859 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n13 GND 0.26539f
C6860 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n14 GND 0.29049f
C6861 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t4 GND 0.03763f
C6862 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n15 GND 0.35844f
C6863 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n16 GND 0.43211f
C6864 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t15 GND 0.03758f
C6865 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n17 GND 0.19468f
C6866 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t2 GND 0.03758f
C6867 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n18 GND 0.19468f
C6868 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n19 GND 0.1431f
C6869 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t19 GND 0.03763f
C6870 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t8 GND 0.03763f
C6871 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n20 GND 0.55306f
C6872 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n21 GND 0.43211f
C6873 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t1 GND 0.03758f
C6874 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n22 GND 0.19468f
C6875 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t9 GND 0.03758f
C6876 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n23 GND 0.19468f
C6877 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n24 GND 0.16566f
C6878 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n25 GND 0.24058f
C6879 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n26 GND 0.91514f
C6880 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n27 GND 0.18865f
C6881 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t10 GND 0.03764f
C6882 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t11 GND 0.14374f
C6883 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n28 GND 3.02823f
C6884 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n29 GND 0.32533f
C6885 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t28 GND 0.19022f
C6886 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t63 GND 0.18766f
C6887 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n30 GND 0.5957f
C6888 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t43 GND 0.18766f
C6889 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n31 GND 0.23386f
C6890 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t30 GND 0.18766f
C6891 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n32 GND 0.23386f
C6892 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t68 GND 0.18766f
C6893 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n33 GND 0.23386f
C6894 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t46 GND 0.18766f
C6895 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n34 GND 0.23386f
C6896 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t45 GND 0.18766f
C6897 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n35 GND 0.23386f
C6898 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t25 GND 0.18766f
C6899 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n36 GND 0.21251f
C6900 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t23 GND 0.18766f
C6901 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n37 GND 0.35069f
C6902 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t24 GND 0.18766f
C6903 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n38 GND 0.23386f
C6904 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t44 GND 0.18766f
C6905 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n39 GND 0.23386f
C6906 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t64 GND 0.18766f
C6907 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n40 GND 0.23386f
C6908 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t66 GND 0.18766f
C6909 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n41 GND 0.23386f
C6910 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t42 GND 0.18766f
C6911 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n42 GND 0.23386f
C6912 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t48 GND 0.18766f
C6913 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n43 GND 0.18995f
C6914 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t77 GND 0.1893f
C6915 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t76 GND 0.18766f
C6916 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n44 GND 0.46608f
C6917 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t56 GND 0.18766f
C6918 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n45 GND 0.23386f
C6919 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t35 GND 0.18766f
C6920 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n46 GND 0.23386f
C6921 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t81 GND 0.18766f
C6922 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n47 GND 0.23386f
C6923 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t59 GND 0.18766f
C6924 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n48 GND 0.23386f
C6925 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t37 GND 0.18766f
C6926 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n49 GND 0.23386f
C6927 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t36 GND 0.18766f
C6928 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n50 GND 0.23386f
C6929 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t74 GND 0.18766f
C6930 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n51 GND 0.21251f
C6931 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n52 GND 0.0734f
C6932 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n53 GND 0.27713f
C6933 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n54 GND 0.06527f
C6934 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t55 GND 0.18766f
C6935 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n55 GND 0.18995f
C6936 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t50 GND 0.18766f
C6937 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n56 GND 0.23386f
C6938 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t73 GND 0.18766f
C6939 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n57 GND 0.23386f
C6940 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t71 GND 0.18766f
C6941 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n58 GND 0.23386f
C6942 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t52 GND 0.18766f
C6943 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n59 GND 0.23386f
C6944 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t31 GND 0.18766f
C6945 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n60 GND 0.44501f
C6946 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n61 GND 0.25344f
C6947 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t53 GND 0.19022f
C6948 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t33 GND 0.18766f
C6949 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n62 GND 0.5957f
C6950 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t69 GND 0.18766f
C6951 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n63 GND 0.23386f
C6952 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t54 GND 0.18766f
C6953 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n64 GND 0.23386f
C6954 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t34 GND 0.18766f
C6955 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n65 GND 0.23386f
C6956 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t72 GND 0.18766f
C6957 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n66 GND 0.23386f
C6958 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t70 GND 0.18766f
C6959 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n67 GND 0.23386f
C6960 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t51 GND 0.18766f
C6961 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n68 GND 0.21251f
C6962 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n69 GND 0.06527f
C6963 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t26 GND 0.18766f
C6964 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n70 GND 0.18995f
C6965 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t75 GND 0.18766f
C6966 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n71 GND 0.23386f
C6967 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t40 GND 0.18766f
C6968 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n72 GND 0.23386f
C6969 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t39 GND 0.18766f
C6970 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n73 GND 0.23386f
C6971 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t79 GND 0.18766f
C6972 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n74 GND 0.23386f
C6973 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t57 GND 0.18766f
C6974 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n75 GND 0.44501f
C6975 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n76 GND 0.3724f
C6976 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t65 GND 0.18766f
C6977 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n77 GND 0.35885f
C6978 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t67 GND 0.18766f
C6979 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n78 GND 0.23386f
C6980 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t29 GND 0.18766f
C6981 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n79 GND 0.23386f
C6982 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t47 GND 0.18766f
C6983 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n80 GND 0.23386f
C6984 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t49 GND 0.18766f
C6985 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n81 GND 0.23386f
C6986 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t27 GND 0.18766f
C6987 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n82 GND 0.23386f
C6988 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t32 GND 0.18766f
C6989 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n83 GND 0.18995f
C6990 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t61 GND 0.1893f
C6991 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t60 GND 0.18766f
C6992 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n84 GND 0.46608f
C6993 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t38 GND 0.18766f
C6994 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n85 GND 0.23386f
C6995 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t78 GND 0.18766f
C6996 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n86 GND 0.23386f
C6997 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t62 GND 0.18766f
C6998 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n87 GND 0.23386f
C6999 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t41 GND 0.18766f
C7000 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n88 GND 0.23386f
C7001 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t22 GND 0.18766f
C7002 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n89 GND 0.23386f
C7003 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t80 GND 0.18766f
C7004 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n90 GND 0.23386f
C7005 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t58 GND 0.18766f
C7006 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n91 GND 0.21251f
C7007 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n92 GND 0.06527f
C7008 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n93 GND 0.1306f
C7009 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t12 GND 0.07099f
C7010 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t18 GND 0.0702f
C7011 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n0 GND 0.14656f
C7012 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t17 GND 0.0702f
C7013 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n1 GND 0.06927f
C7014 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t24 GND 0.0702f
C7015 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n2 GND 0.06927f
C7016 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t23 GND 0.0702f
C7017 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n3 GND 0.06927f
C7018 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t13 GND 0.0702f
C7019 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n4 GND 0.06927f
C7020 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t6 GND 0.0702f
C7021 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n5 GND 0.06927f
C7022 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t8 GND 0.0702f
C7023 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n6 GND 0.06927f
C7024 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t25 GND 0.0702f
C7025 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n7 GND 0.06927f
C7026 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t15 GND 0.0702f
C7027 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n8 GND 0.06927f
C7028 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t7 GND 0.0702f
C7029 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n9 GND 0.06927f
C7030 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t20 GND 0.0702f
C7031 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n10 GND 0.06927f
C7032 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t14 GND 0.0702f
C7033 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n11 GND 0.06927f
C7034 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t27 GND 0.0702f
C7035 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n12 GND 0.06927f
C7036 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t19 GND 0.0702f
C7037 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n13 GND 0.06927f
C7038 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t10 GND 0.0702f
C7039 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n14 GND 0.06927f
C7040 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t26 GND 0.0702f
C7041 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n15 GND 0.06927f
C7042 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t16 GND 0.0702f
C7043 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n16 GND 0.06927f
C7044 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t9 GND 0.0702f
C7045 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n17 GND 0.06927f
C7046 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t22 GND 0.0702f
C7047 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n18 GND 0.06927f
C7048 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t21 GND 0.0702f
C7049 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n19 GND 0.06927f
C7050 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t28 GND 0.0702f
C7051 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n20 GND 0.06641f
C7052 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t11 GND 0.27283f
C7053 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n21 GND 0.09448f
C7054 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n22 GND 0.55544f
C7055 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t4 GND 0.04839f
C7056 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n23 GND 0.0364f
C7057 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n24 GND 0.04636f
C7058 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t2 GND 0.04832f
C7059 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n25 GND 0.02822f
C7060 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n26 GND 0.18252f
C7061 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t1 GND 0.0317f
C7062 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n27 GND 0.18304f
C7063 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t0 GND 0.03062f
C7064 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n28 GND 0.1181f
C7065 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.t1 GND 0.115f
C7066 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.t2 GND 0.10649f
C7067 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.n0 GND 1.95995f
C7068 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1.t0 GND 0.01856f
C7069 a_21927_20174.t3 GND 0.14562f
C7070 a_21927_20174.t1 GND 0.05846f
C7071 a_21927_20174.n0 GND 4.28874f
C7072 a_21927_20174.t2 GND 0.0771f
C7073 a_21927_20174.n1 GND 5.74363f
C7074 a_21927_20174.t0 GND 0.18645f
C7075 a_23629_18133.t5 GND 0.07067f
C7076 a_23629_18133.t3 GND 0.05945f
C7077 a_23629_18133.n0 GND 2.30243f
C7078 a_23629_18133.t2 GND 0.05945f
C7079 a_23629_18133.n1 GND 1.38823f
C7080 a_23629_18133.t1 GND 0.06045f
C7081 a_23629_18133.t4 GND 0.05907f
C7082 a_23629_18133.n2 GND 1.47888f
C7083 a_23629_18133.n3 GND 1.3619f
C7084 a_23629_18133.t0 GND 0.05945f
C7085 VDDH.n0 GND 10.6957f
C7086 VDDH.n2 GND 0.06535f
C7087 VDDH.t438 GND 0.08077f
C7088 VDDH.n5 GND 0.05513f
C7089 VDDH.n7 GND 0.06535f
C7090 VDDH.t504 GND 0.12385f
C7091 VDDH.n8 GND 0.04286f
C7092 VDDH.t516 GND 0.12385f
C7093 VDDH.n9 GND 0.04286f
C7094 VDDH.t573 GND 0.12385f
C7095 VDDH.n10 GND 0.04286f
C7096 VDDH.t436 GND 0.08077f
C7097 VDDH.n11 GND 0.05513f
C7098 VDDH.n13 GND 0.05722f
C7099 VDDH.n21 GND 0.05722f
C7100 VDDH.n22 GND 0.31817f
C7101 VDDH.t80 GND 0.01129f
C7102 VDDH.n24 GND 0.01665f
C7103 VDDH.n27 GND 0.04287f
C7104 VDDH.t81 GND 0.13243f
C7105 VDDH.t536 GND 0.01129f
C7106 VDDH.n32 GND 0.01665f
C7107 VDDH.n35 GND 0.04287f
C7108 VDDH.t537 GND 0.13243f
C7109 VDDH.n41 GND 0.05513f
C7110 VDDH.n43 GND 0.0554f
C7111 VDDH.n44 GND 0.04868f
C7112 VDDH.t428 GND 0.04153f
C7113 VDDH.n49 GND 0.04421f
C7114 VDDH.t354 GND 0.04287f
C7115 VDDH.n56 GND 0.0196f
C7116 VDDH.n59 GND 0.22505f
C7117 VDDH.t380 GND 0.42845f
C7118 VDDH.n67 GND 0.01157f
C7119 VDDH.n69 GND 0.0196f
C7120 VDDH.n70 GND 0.01157f
C7121 VDDH.n71 GND 0.0196f
C7122 VDDH.n73 GND 0.01157f
C7123 VDDH.n74 GND 0.0196f
C7124 VDDH.n77 GND 0.01157f
C7125 VDDH.n79 GND 0.01543f
C7126 VDDH.t452 GND 0.01129f
C7127 VDDH.n80 GND 0.03783f
C7128 VDDH.n81 GND 0.0164f
C7129 VDDH.n82 GND 0.02042f
C7130 VDDH.n87 GND 0.01543f
C7131 VDDH.t381 GND 0.01129f
C7132 VDDH.n88 GND 0.03783f
C7133 VDDH.n90 GND 0.04373f
C7134 VDDH.t365 GND 0.61416f
C7135 VDDH.n91 GND 0.1312f
C7136 VDDH.n92 GND 0.09959f
C7137 VDDH.n93 GND 0.09715f
C7138 VDDH.n94 GND 0.08537f
C7139 VDDH.n95 GND 0.02362f
C7140 VDDH.n96 GND 0.01687f
C7141 VDDH.n97 GND 0.02085f
C7142 VDDH.n98 GND 0.0146f
C7143 VDDH.n99 GND 0.03841f
C7144 VDDH.n100 GND 0.0679f
C7145 VDDH.n101 GND 0.05925f
C7146 VDDH.n102 GND 0.05437f
C7147 VDDH.n103 GND 0.05955f
C7148 VDDH.t236 GND 0.01754f
C7149 VDDH.t237 GND 0.01754f
C7150 VDDH.n104 GND 0.05822f
C7151 VDDH.t235 GND 0.06625f
C7152 VDDH.n105 GND 0.07705f
C7153 VDDH.t212 GND 0.01754f
C7154 VDDH.t213 GND 0.01754f
C7155 VDDH.n106 GND 0.05822f
C7156 VDDH.t211 GND 0.06625f
C7157 VDDH.n107 GND 0.07705f
C7158 VDDH.n108 GND 0.15954f
C7159 VDDH.n109 GND 0.10721f
C7160 VDDH.n110 GND 0.04469f
C7161 VDDH.n111 GND 0.39649f
C7162 VDDH.n112 GND 0.03771f
C7163 VDDH.t210 GND 0.01754f
C7164 VDDH.t116 GND 0.01754f
C7165 VDDH.t115 GND 0.01754f
C7166 VDDH.n113 GND 0.05822f
C7167 VDDH.t113 GND 0.06625f
C7168 VDDH.n114 GND 0.07705f
C7169 VDDH.t580 GND 0.01744f
C7170 VDDH.t209 GND 0.01744f
C7171 VDDH.n115 GND 0.06225f
C7172 VDDH.t57 GND 0.01744f
C7173 VDDH.t582 GND 0.01744f
C7174 VDDH.n116 GND 0.07069f
C7175 VDDH.t583 GND 0.01744f
C7176 VDDH.t347 GND 0.01744f
C7177 VDDH.n117 GND 0.07036f
C7178 VDDH.n118 GND 0.06285f
C7179 VDDH.n119 GND 0.03229f
C7180 VDDH.n120 GND 0.05663f
C7181 VDDH.n121 GND 0.07958f
C7182 VDDH.t56 GND 0.6f
C7183 VDDH.n122 GND 0.1047f
C7184 VDDH.n123 GND 0.02997f
C7185 VDDH.t581 GND 0.01744f
C7186 VDDH.t271 GND 0.01744f
C7187 VDDH.n124 GND 0.07069f
C7188 VDDH.n125 GND 0.0567f
C7189 VDDH.t272 GND 0.01744f
C7190 VDDH.t584 GND 0.01744f
C7191 VDDH.n126 GND 0.07069f
C7192 VDDH.t167 GND 0.01754f
C7193 VDDH.t185 GND 0.01754f
C7194 VDDH.t186 GND 0.01744f
C7195 VDDH.t346 GND 0.01744f
C7196 VDDH.n127 GND 0.06795f
C7197 VDDH.n128 GND 0.0612f
C7198 VDDH.t184 GND 0.06625f
C7199 VDDH.n129 GND 0.03408f
C7200 VDDH.n130 GND 0.04346f
C7201 VDDH.n131 GND 0.21942f
C7202 VDDH.n132 GND 0.15007f
C7203 VDDH.t230 GND 0.01754f
C7204 VDDH.t231 GND 0.01754f
C7205 VDDH.n133 GND 0.05822f
C7206 VDDH.t229 GND 0.06625f
C7207 VDDH.n134 GND 0.03339f
C7208 VDDH.t132 GND 0.01754f
C7209 VDDH.t131 GND 0.01754f
C7210 VDDH.n135 GND 0.05822f
C7211 VDDH.t129 GND 0.06625f
C7212 VDDH.n136 GND 0.08254f
C7213 VDDH.n137 GND 0.08786f
C7214 VDDH.n138 GND 0.1368f
C7215 VDDH.n139 GND 0.05275f
C7216 VDDH.n140 GND 0.09672f
C7217 VDDH.n141 GND 0.17039f
C7218 VDDH.n142 GND 0.02942f
C7219 VDDH.n143 GND 0.17173f
C7220 VDDH.n144 GND 0.49789f
C7221 VDDH.t417 GND 0.25392f
C7222 VDDH.t368 GND 0.32806f
C7223 VDDH.t418 GND 0.25392f
C7224 VDDH.t425 GND 0.74129f
C7225 VDDH.t382 GND 1.25867f
C7226 VDDH.t66 GND 0.42448f
C7227 VDDH.n145 GND 0.31426f
C7228 VDDH.t256 GND 0.41701f
C7229 VDDH.t538 GND 0.68764f
C7230 VDDH.t252 GND 0.5515f
C7231 VDDH.n147 GND 0.30827f
C7232 VDDH.t257 GND 0.34151f
C7233 VDDH.t392 GND 1.00146f
C7234 VDDH.n148 GND 0.72687f
C7235 VDDH.t338 GND 0.16284f
C7236 VDDH.t16 GND 3.09288f
C7237 VDDH.n149 GND 0.42567f
C7238 VDDH.n151 GND 0.15302f
C7239 VDDH.n152 GND 0.10138f
C7240 VDDH.n153 GND 0.09125f
C7241 VDDH.n154 GND 0.04141f
C7242 VDDH.n155 GND 0.03617f
C7243 VDDH.n156 GND 0.06762f
C7244 VDDH.n157 GND 0.01731f
C7245 VDDH.n159 GND 0.03764f
C7246 VDDH.n160 GND 0.81531f
C7247 VDDH.t466 GND 0.75794f
C7248 VDDH.t467 GND 0.75794f
C7249 VDDH.t251 GND 0.57415f
C7250 VDDH.n161 GND 0.53569f
C7251 VDDH.t30 GND 1.0329f
C7252 VDDH.t130 GND 0.88046f
C7253 VDDH.n163 GND 0.06711f
C7254 VDDH.n164 GND 0.56418f
C7255 VDDH.n165 GND 0.60977f
C7256 VDDH.n166 GND 0.08939f
C7257 VDDH.n167 GND 0.05077f
C7258 VDDH.n168 GND 0.05938f
C7259 VDDH.n169 GND 0.10165f
C7260 VDDH.n170 GND 0.18179f
C7261 VDDH.n171 GND 0.11596f
C7262 VDDH.n172 GND 1.95847f
C7263 VDDH.n173 GND 2.67348f
C7264 VDDH.t179 GND 0.01755f
C7265 VDDH.n174 GND 0.04261f
C7266 VDDH.n175 GND 0.27467f
C7267 VDDH.n176 GND 0.16036f
C7268 VDDH.n177 GND 0.08962f
C7269 VDDH.n178 GND 0.28316f
C7270 VDDH.n179 GND 0.15815f
C7271 VDDH.n180 GND 0.15866f
C7272 VDDH.n181 GND 2.74454f
C7273 VDDH.n182 GND 0.462f
C7274 VDDH.n183 GND 0.24856f
C7275 VDDH.n184 GND 0.24856f
C7276 VDDH.t540 GND 0.66812f
C7277 VDDH.n185 GND 0.29505f
C7278 VDDH.n186 GND 0.24856f
C7279 VDDH.n187 GND 0.15266f
C7280 VDDH.n188 GND 0.15266f
C7281 VDDH.n189 GND 0.07971f
C7282 VDDH.n190 GND 0.07946f
C7283 VDDH.t569 GND 0.01744f
C7284 VDDH.t296 GND 0.01744f
C7285 VDDH.n191 GND 0.06773f
C7286 VDDH.t385 GND 0.01744f
C7287 VDDH.t565 GND 0.01744f
C7288 VDDH.n192 GND 0.06773f
C7289 VDDH.n193 GND 0.14681f
C7290 VDDH.t362 GND 0.01744f
C7291 VDDH.t267 GND 0.01744f
C7292 VDDH.n194 GND 0.06773f
C7293 VDDH.n195 GND 0.14473f
C7294 VDDH.n196 GND 0.28316f
C7295 VDDH.n198 GND 0.04219f
C7296 VDDH.n199 GND 0.11165f
C7297 VDDH.n200 GND 0.03677f
C7298 VDDH.t135 GND 0.01754f
C7299 VDDH.t164 GND 0.01757f
C7300 VDDH.t162 GND 0.06625f
C7301 VDDH.t165 GND 0.01757f
C7302 VDDH.t269 GND 0.01744f
C7303 VDDH.t96 GND 0.01744f
C7304 VDDH.n201 GND 0.06225f
C7305 VDDH.t507 GND 0.01744f
C7306 VDDH.t282 GND 0.01744f
C7307 VDDH.n202 GND 0.06773f
C7308 VDDH.t283 GND 0.01744f
C7309 VDDH.t239 GND 0.01744f
C7310 VDDH.n203 GND 0.06773f
C7311 VDDH.t295 GND 0.01744f
C7312 VDDH.t43 GND 0.01744f
C7313 VDDH.n204 GND 0.06773f
C7314 VDDH.n205 GND 0.14681f
C7315 VDDH.n206 GND 0.14681f
C7316 VDDH.n207 GND 0.14524f
C7317 VDDH.n208 GND 0.10781f
C7318 VDDH.t95 GND 0.06625f
C7319 VDDH.n209 GND 0.06155f
C7320 VDDH.t97 GND 0.01744f
C7321 VDDH.t94 GND 0.01744f
C7322 VDDH.t207 GND 0.01744f
C7323 VDDH.t90 GND 0.01744f
C7324 VDDH.n210 GND 0.07543f
C7325 VDDH.t205 GND 0.06625f
C7326 VDDH.t92 GND 0.06625f
C7327 VDDH.n211 GND 0.06812f
C7328 VDDH.t88 GND 0.06625f
C7329 VDDH.t128 GND 0.01754f
C7330 VDDH.t91 GND 0.01754f
C7331 VDDH.n212 GND 0.05415f
C7332 VDDH.n214 GND 0.14084f
C7333 VDDH.n215 GND 0.01273f
C7334 VDDH.n216 GND 0.05382f
C7335 VDDH.t216 GND 0.01762f
C7336 VDDH.t214 GND 0.06625f
C7337 VDDH.n217 GND 0.05371f
C7338 VDDH.t176 GND 0.01762f
C7339 VDDH.t175 GND 0.06625f
C7340 VDDH.n218 GND 0.05371f
C7341 VDDH.t177 GND 0.01744f
C7342 VDDH.t215 GND 0.01744f
C7343 VDDH.n219 GND 0.06395f
C7344 VDDH.n220 GND 0.04225f
C7345 VDDH.t222 GND 0.01762f
C7346 VDDH.t220 GND 0.06625f
C7347 VDDH.n221 GND 0.05371f
C7348 VDDH.t182 GND 0.01762f
C7349 VDDH.t181 GND 0.06625f
C7350 VDDH.n222 GND 0.05371f
C7351 VDDH.t183 GND 0.01744f
C7352 VDDH.t221 GND 0.01744f
C7353 VDDH.n223 GND 0.06395f
C7354 VDDH.n224 GND 0.04225f
C7355 VDDH.n225 GND 0.19792f
C7356 VDDH.n226 GND 0.09499f
C7357 VDDH.n227 GND 0.02111f
C7358 VDDH.n228 GND 0.16791f
C7359 VDDH.t85 GND 1.69518f
C7360 VDDH.n229 GND 0.07302f
C7361 VDDH.n230 GND 0.07302f
C7362 VDDH.n231 GND 0.09549f
C7363 VDDH.n232 GND 0.02914f
C7364 VDDH.n233 GND 0.0411f
C7365 VDDH.n234 GND 0.07218f
C7366 VDDH.n235 GND 0.07218f
C7367 VDDH.t327 GND 0.51886f
C7368 VDDH.t337 GND 0.81738f
C7369 VDDH.n236 GND 0.07218f
C7370 VDDH.t42 GND 0.91689f
C7371 VDDH.t335 GND 1.33624f
C7372 VDDH.t52 GND 1.69518f
C7373 VDDH.t558 GND 1.33624f
C7374 VDDH.t268 GND 0.91689f
C7375 VDDH.t286 GND 1.33624f
C7376 VDDH.t50 GND 0.45844f
C7377 VDDH.n237 GND 0.47977f
C7378 VDDH.t325 GND 1.31492f
C7379 VDDH.t277 GND 0.91689f
C7380 VDDH.t559 GND 1.33624f
C7381 VDDH.t238 GND 1.69518f
C7382 VDDH.n238 GND 1.33624f
C7383 VDDH.n239 GND 0.05072f
C7384 VDDH.n240 GND 0.07218f
C7385 VDDH.t288 GND 1.57435f
C7386 VDDH.t54 GND 1.45707f
C7387 VDDH.t287 GND 0.91689f
C7388 VDDH.t336 GND 1.33624f
C7389 VDDH.t266 GND 1.69518f
C7390 VDDH.n241 GND 1.33624f
C7391 VDDH.n242 GND 0.05072f
C7392 VDDH.n243 GND 0.02914f
C7393 VDDH.n244 GND 0.07552f
C7394 VDDH.n245 GND 0.37714f
C7395 VDDH.n246 GND 0.01235f
C7396 VDDH.n247 GND 0.08734f
C7397 VDDH.n248 GND 0.09204f
C7398 VDDH.n249 GND 0.01235f
C7399 VDDH.t100 GND 0.01754f
C7400 VDDH.n250 GND 0.04171f
C7401 VDDH.n251 GND 0.24572f
C7402 VDDH.n252 GND 0.15304f
C7403 VDDH.n253 GND 0.16184f
C7404 VDDH.n254 GND 0.16707f
C7405 VDDH.t99 GND 1.69518f
C7406 VDDH.n255 GND 0.07302f
C7407 VDDH.n256 GND 0.07302f
C7408 VDDH.n257 GND 0.02653f
C7409 VDDH.n258 GND 0.11435f
C7410 VDDH.n259 GND 0.07345f
C7411 VDDH.n260 GND 0.07218f
C7412 VDDH.n261 GND 0.07218f
C7413 VDDH.t543 GND 1.33624f
C7414 VDDH.t103 GND 0.91689f
C7415 VDDH.t542 GND 0.80317f
C7416 VDDH.n262 GND 0.91689f
C7417 VDDH.t326 GND 0.53308f
C7418 VDDH.t279 GND 0.91689f
C7419 VDDH.t544 GND 1.33624f
C7420 VDDH.t46 GND 1.69518f
C7421 VDDH.n263 GND 0.04682f
C7422 VDDH.t453 GND 1.07326f
C7423 VDDH.n264 GND 0.04682f
C7424 VDDH.n265 GND 0.07218f
C7425 VDDH.n266 GND 0.0411f
C7426 VDDH.n267 GND 0.02653f
C7427 VDDH.n268 GND 0.04682f
C7428 VDDH.n269 GND 0.07218f
C7429 VDDH.t44 GND 0.91689f
C7430 VDDH.t454 GND 1.33624f
C7431 VDDH.t262 GND 1.69518f
C7432 VDDH.t320 GND 1.05904f
C7433 VDDH.t301 GND 0.91689f
C7434 VDDH.t541 GND 1.33624f
C7435 VDDH.t48 GND 1.69518f
C7436 VDDH.n270 GND 1.33624f
C7437 VDDH.n271 GND 0.05072f
C7438 VDDH.n272 GND 0.02914f
C7439 VDDH.n273 GND 0.07345f
C7440 VDDH.n274 GND 0.11435f
C7441 VDDH.n275 GND 0.04682f
C7442 VDDH.n276 GND 0.72143f
C7443 VDDH.t297 GND 0.45844f
C7444 VDDH.t455 GND 1.11235f
C7445 VDDH.t245 GND 1.14078f
C7446 VDDH.t275 GND 1.56013f
C7447 VDDH.t291 GND 1.47129f
C7448 VDDH.n277 GND 1.33624f
C7449 VDDH.n278 GND 0.05072f
C7450 VDDH.n279 GND 0.02914f
C7451 VDDH.n280 GND 0.0411f
C7452 VDDH.n281 GND 0.04137f
C7453 VDDH.n282 GND 0.04265f
C7454 VDDH.n283 GND 0.0991f
C7455 VDDH.n284 GND 0.93466f
C7456 VDDH.n285 GND 0.16791f
C7457 VDDH.n286 GND 0.04274f
C7458 VDDH.n287 GND 0.67878f
C7459 VDDH.n288 GND 0.02787f
C7460 VDDH.n291 GND 0.08728f
C7461 VDDH.t302 GND 0.01744f
C7462 VDDH.t274 GND 0.01744f
C7463 VDDH.n292 GND 0.0818f
C7464 VDDH.t552 GND 0.01744f
C7465 VDDH.t554 GND 0.01744f
C7466 VDDH.n293 GND 0.0818f
C7467 VDDH.t263 GND 0.01744f
C7468 VDDH.t49 GND 0.01744f
C7469 VDDH.n294 GND 0.0818f
C7470 VDDH.t305 GND 0.01744f
C7471 VDDH.t510 GND 0.01744f
C7472 VDDH.n295 GND 0.0818f
C7473 VDDH.t388 GND 0.01744f
C7474 VDDH.t45 GND 0.01744f
C7475 VDDH.n296 GND 0.0818f
C7476 VDDH.t298 GND 0.01744f
C7477 VDDH.t572 GND 0.01744f
C7478 VDDH.n297 GND 0.0818f
C7479 VDDH.t363 GND 0.01744f
C7480 VDDH.t315 GND 0.01744f
C7481 VDDH.n298 GND 0.0818f
C7482 VDDH.t389 GND 0.01744f
C7483 VDDH.t570 GND 0.01744f
C7484 VDDH.n299 GND 0.0818f
C7485 VDDH.t318 GND 0.01744f
C7486 VDDH.t293 GND 0.01744f
C7487 VDDH.n300 GND 0.0818f
C7488 VDDH.t300 GND 0.01744f
C7489 VDDH.t319 GND 0.01744f
C7490 VDDH.n301 GND 0.0818f
C7491 VDDH.t198 GND 0.01754f
C7492 VDDH.t174 GND 0.01754f
C7493 VDDH.t112 GND 0.01744f
C7494 VDDH.t101 GND 0.01744f
C7495 VDDH.t98 GND 0.06625f
C7496 VDDH.n302 GND 0.03408f
C7497 VDDH.t105 GND 0.01762f
C7498 VDDH.t102 GND 0.06625f
C7499 VDDH.n303 GND 0.05371f
C7500 VDDH.t203 GND 0.01762f
C7501 VDDH.t202 GND 0.06625f
C7502 VDDH.n304 GND 0.05371f
C7503 VDDH.t204 GND 0.01744f
C7504 VDDH.t104 GND 0.01744f
C7505 VDDH.n305 GND 0.06395f
C7506 VDDH.n306 GND 0.04499f
C7507 VDDH.t158 GND 0.01744f
C7508 VDDH.t280 GND 0.01744f
C7509 VDDH.n307 GND 0.06795f
C7510 VDDH.t265 GND 0.01744f
C7511 VDDH.t292 GND 0.01744f
C7512 VDDH.n308 GND 0.07069f
C7513 VDDH.t276 GND 0.01744f
C7514 VDDH.t313 GND 0.01744f
C7515 VDDH.n309 GND 0.07069f
C7516 VDDH.t317 GND 0.01744f
C7517 VDDH.t281 GND 0.01744f
C7518 VDDH.n310 GND 0.07069f
C7519 VDDH.t261 GND 0.01744f
C7520 VDDH.t556 GND 0.01744f
C7521 VDDH.n311 GND 0.07069f
C7522 VDDH.t234 GND 0.01754f
C7523 VDDH.n312 GND 0.04317f
C7524 VDDH.t232 GND 0.06625f
C7525 VDDH.n313 GND 0.03408f
C7526 VDDH.t195 GND 0.01744f
C7527 VDDH.t233 GND 0.01744f
C7528 VDDH.n314 GND 0.08113f
C7529 VDDH.t189 GND 0.01762f
C7530 VDDH.t187 GND 0.06625f
C7531 VDDH.n315 GND 0.05371f
C7532 VDDH.t154 GND 0.01762f
C7533 VDDH.t153 GND 0.06625f
C7534 VDDH.n316 GND 0.05371f
C7535 VDDH.t155 GND 0.01744f
C7536 VDDH.t188 GND 0.01744f
C7537 VDDH.n317 GND 0.06395f
C7538 VDDH.n318 GND 0.04499f
C7539 VDDH.n319 GND 0.05933f
C7540 VDDH.t193 GND 0.06625f
C7541 VDDH.n320 GND 0.03249f
C7542 VDDH.t555 GND 0.01744f
C7543 VDDH.t194 GND 0.01744f
C7544 VDDH.n321 GND 0.06795f
C7545 VDDH.n322 GND 0.0612f
C7546 VDDH.t278 GND 0.01744f
C7547 VDDH.t51 GND 0.01744f
C7548 VDDH.n323 GND 0.07069f
C7549 VDDH.n324 GND 0.07411f
C7550 VDDH.t53 GND 0.01744f
C7551 VDDH.t306 GND 0.01744f
C7552 VDDH.n325 GND 0.07069f
C7553 VDDH.n326 GND 0.07322f
C7554 VDDH.t303 GND 0.01744f
C7555 VDDH.t264 GND 0.01744f
C7556 VDDH.n327 GND 0.07069f
C7557 VDDH.n328 GND 0.07322f
C7558 VDDH.t294 GND 0.01744f
C7559 VDDH.t551 GND 0.01744f
C7560 VDDH.n329 GND 0.07069f
C7561 VDDH.n330 GND 0.07322f
C7562 VDDH.t557 GND 0.01744f
C7563 VDDH.t304 GND 0.01744f
C7564 VDDH.n331 GND 0.07069f
C7565 VDDH.n332 GND 0.07322f
C7566 VDDH.n333 GND 0.07322f
C7567 VDDH.n334 GND 0.07322f
C7568 VDDH.n335 GND 0.07322f
C7569 VDDH.n336 GND 0.07411f
C7570 VDDH.n337 GND 0.0612f
C7571 VDDH.t156 GND 0.06625f
C7572 VDDH.n338 GND 0.03249f
C7573 VDDH.n339 GND 0.05933f
C7574 VDDH.t157 GND 0.01744f
C7575 VDDH.n340 GND 0.08113f
C7576 VDDH.t173 GND 0.01744f
C7577 VDDH.n341 GND 0.07543f
C7578 VDDH.t151 GND 0.01754f
C7579 VDDH.t111 GND 0.01754f
C7580 VDDH.n342 GND 0.07518f
C7581 VDDH.t110 GND 0.06625f
C7582 VDDH.t150 GND 0.06625f
C7583 VDDH.n343 GND 0.06812f
C7584 VDDH.t218 GND 0.01757f
C7585 VDDH.t217 GND 0.06625f
C7586 VDDH.t219 GND 0.01757f
C7587 VDDH.t170 GND 0.01754f
C7588 VDDH.n346 GND 0.28031f
C7589 VDDH.n347 GND 0.25384f
C7590 VDDH.n348 GND 0.28765f
C7591 VDDH.n349 GND 0.0523f
C7592 VDDH.t169 GND 0.06625f
C7593 VDDH.n350 GND 0.03778f
C7594 VDDH.n351 GND 0.1144f
C7595 VDDH.t201 GND 0.01744f
C7596 VDDH.t508 GND 0.01744f
C7597 VDDH.n352 GND 0.06225f
C7598 VDDH.t47 GND 0.01744f
C7599 VDDH.t358 GND 0.01744f
C7600 VDDH.n353 GND 0.06773f
C7601 VDDH.t571 GND 0.01744f
C7602 VDDH.t383 GND 0.01744f
C7603 VDDH.n354 GND 0.06773f
C7604 VDDH.t384 GND 0.01744f
C7605 VDDH.t513 GND 0.01744f
C7606 VDDH.n355 GND 0.06773f
C7607 VDDH.n356 GND 0.14681f
C7608 VDDH.n357 GND 0.14681f
C7609 VDDH.n358 GND 0.14524f
C7610 VDDH.n359 GND 0.10781f
C7611 VDDH.t199 GND 0.06625f
C7612 VDDH.n360 GND 0.06155f
C7613 VDDH.n361 GND 0.05516f
C7614 VDDH.t171 GND 0.01744f
C7615 VDDH.t200 GND 0.01744f
C7616 VDDH.n362 GND 0.07543f
C7617 VDDH.t152 GND 0.01744f
C7618 VDDH.t197 GND 0.01744f
C7619 VDDH.n363 GND 0.07543f
C7620 VDDH.n364 GND 0.07145f
C7621 VDDH.t172 GND 0.06625f
C7622 VDDH.t196 GND 0.06625f
C7623 VDDH.n365 GND 0.06812f
C7624 VDDH.n366 GND 0.08466f
C7625 VDDH.n367 GND 0.08312f
C7626 VDDH.n368 GND 0.0921f
C7627 VDDH.n369 GND 0.0921f
C7628 VDDH.n370 GND 0.0921f
C7629 VDDH.n371 GND 0.08148f
C7630 VDDH.t93 GND 0.01754f
C7631 VDDH.t206 GND 0.01754f
C7632 VDDH.n372 GND 0.08466f
C7633 VDDH.t359 GND 0.01744f
C7634 VDDH.t568 GND 0.01744f
C7635 VDDH.n373 GND 0.0818f
C7636 VDDH.t386 GND 0.01744f
C7637 VDDH.t364 GND 0.01744f
C7638 VDDH.n374 GND 0.0818f
C7639 VDDH.n375 GND 0.08312f
C7640 VDDH.t512 GND 0.01744f
C7641 VDDH.t316 GND 0.01744f
C7642 VDDH.n376 GND 0.0818f
C7643 VDDH.t567 GND 0.01744f
C7644 VDDH.t299 GND 0.01744f
C7645 VDDH.n377 GND 0.0818f
C7646 VDDH.n378 GND 0.0921f
C7647 VDDH.t290 GND 0.01744f
C7648 VDDH.t361 GND 0.01744f
C7649 VDDH.n379 GND 0.0818f
C7650 VDDH.t314 GND 0.01744f
C7651 VDDH.t387 GND 0.01744f
C7652 VDDH.n380 GND 0.0818f
C7653 VDDH.n381 GND 0.0921f
C7654 VDDH.t270 GND 0.01744f
C7655 VDDH.t509 GND 0.01744f
C7656 VDDH.n382 GND 0.0818f
C7657 VDDH.t360 GND 0.01744f
C7658 VDDH.t564 GND 0.01744f
C7659 VDDH.n383 GND 0.0818f
C7660 VDDH.n384 GND 0.0921f
C7661 VDDH.t511 GND 0.01744f
C7662 VDDH.t553 GND 0.01744f
C7663 VDDH.n385 GND 0.0818f
C7664 VDDH.t566 GND 0.01744f
C7665 VDDH.t55 GND 0.01744f
C7666 VDDH.n386 GND 0.0818f
C7667 VDDH.n387 GND 0.08148f
C7668 VDDH.n388 GND 0.02124f
C7669 VDDH.n389 GND 0.14084f
C7670 VDDH.n391 GND 0.08653f
C7671 VDDH.n394 GND 0.24262f
C7672 VDDH.n395 GND 0.30711f
C7673 VDDH.n396 GND 0.36522f
C7674 VDDH.n397 GND 0.01331f
C7675 VDDH.n399 GND 0.01331f
C7676 VDDH.n400 GND 0.51342f
C7677 VDDH.t192 GND 0.01762f
C7678 VDDH.t190 GND 0.06625f
C7679 VDDH.n401 GND 0.05371f
C7680 VDDH.t145 GND 0.01762f
C7681 VDDH.t144 GND 0.06625f
C7682 VDDH.n402 GND 0.05371f
C7683 VDDH.t146 GND 0.01744f
C7684 VDDH.t191 GND 0.01744f
C7685 VDDH.n403 GND 0.06395f
C7686 VDDH.n404 GND 0.04225f
C7687 VDDH.n405 GND 0.24766f
C7688 VDDH.t125 GND 0.01762f
C7689 VDDH.t123 GND 0.06625f
C7690 VDDH.n406 GND 0.05371f
C7691 VDDH.t86 GND 0.01762f
C7692 VDDH.t84 GND 0.06625f
C7693 VDDH.n407 GND 0.05371f
C7694 VDDH.t87 GND 0.01744f
C7695 VDDH.t124 GND 0.01744f
C7696 VDDH.n408 GND 0.06395f
C7697 VDDH.n409 GND 0.04225f
C7698 VDDH.n410 GND 0.02475f
C7699 VDDH.t32 GND 0.04838f
C7700 VDDH.n411 GND 0.13558f
C7701 VDDH.n412 GND 0.04959f
C7702 VDDH.n413 GND 0.62619f
C7703 VDDH.n414 GND 0.04911f
C7704 VDDH.n415 GND 0.62619f
C7705 VDDH.t33 GND 0.52131f
C7706 VDDH.t31 GND 0.52131f
C7707 VDDH.n416 GND 0.08782f
C7708 VDDH.n417 GND 0.29662f
C7709 VDDH.n418 GND 0.08782f
C7710 VDDH.t34 GND 0.04838f
C7711 VDDH.n419 GND 0.13558f
C7712 VDDH.n420 GND 0.10507f
C7713 VDDH.n421 GND 0.06803f
C7714 VDDH.n422 GND 0.04959f
C7715 VDDH.n423 GND 0.04911f
C7716 VDDH.n424 GND 0.08886f
C7717 VDDH.n425 GND 0.47554f
C7718 VDDH.n426 GND 0.49034f
C7719 VDDH.n427 GND 0.18488f
C7720 VDDH.n428 GND 0.29291f
C7721 VDDH.n429 GND 0.05661f
C7722 VDDH.n430 GND 0.07345f
C7723 VDDH.n431 GND 0.11549f
C7724 VDDH.n432 GND 0.07345f
C7725 VDDH.n433 GND 0.11435f
C7726 VDDH.n434 GND 0.04682f
C7727 VDDH.n435 GND 0.91689f
C7728 VDDH.n436 GND 0.04682f
C7729 VDDH.n437 GND 0.02653f
C7730 VDDH.n438 GND 0.0411f
C7731 VDDH.n439 GND 0.04137f
C7732 VDDH.n440 GND 0.04265f
C7733 VDDH.n441 GND 0.0991f
C7734 VDDH.n442 GND 0.71788f
C7735 VDDH.t456 GND 2.40236f
C7736 VDDH.t82 GND 2.48287f
C7737 VDDH.n443 GND 3.48648f
C7738 VDDH.t89 GND 0.6827f
C7739 VDDH.t163 GND 0.02288f
C7740 VDDH.t107 GND 0.984f
C7741 VDDH.n444 GND 0.15304f
C7742 VDDH.n445 GND 0.02787f
C7743 VDDH.n446 GND 0.15863f
C7744 VDDH.n447 GND 0.15812f
C7745 VDDH.t108 GND 0.01757f
C7746 VDDH.t106 GND 0.06625f
C7747 VDDH.t109 GND 0.01757f
C7748 VDDH.t180 GND 0.01755f
C7749 VDDH.t178 GND 0.06625f
C7750 VDDH.n448 GND 0.02559f
C7751 VDDH.n449 GND 0.14641f
C7752 VDDH.n450 GND 0.41417f
C7753 VDDH.n451 GND 0.20697f
C7754 VDDH.n452 GND 0.18917f
C7755 VDDH.n453 GND 0.05168f
C7756 VDDH.t403 GND 0.04622f
C7757 VDDH.t527 GND 0.04622f
C7758 VDDH.n454 GND 0.18659f
C7759 VDDH.n455 GND 0.04866f
C7760 VDDH.n456 GND 0.06136f
C7761 VDDH.n457 GND 0.08675f
C7762 VDDH.n458 GND 0.04262f
C7763 VDDH.t404 GND 0.04622f
C7764 VDDH.t402 GND 0.04622f
C7765 VDDH.n459 GND 0.18659f
C7766 VDDH.n460 GND 0.08841f
C7767 VDDH.n461 GND 0.05219f
C7768 VDDH.n462 GND 0.09209f
C7769 VDDH.n463 GND 0.09209f
C7770 VDDH.t345 GND 2.80794f
C7771 VDDH.n464 GND 0.1172f
C7772 VDDH.t401 GND 1.1959f
C7773 VDDH.n465 GND 0.04059f
C7774 VDDH.n466 GND 0.04941f
C7775 VDDH.n467 GND 2.3033f
C7776 VDDH.n468 GND 0.07451f
C7777 VDDH.n469 GND 0.09643f
C7778 VDDH.n470 GND 0.04262f
C7779 VDDH.n471 GND 0.05464f
C7780 VDDH.n472 GND 0.01265f
C7781 VDDH.n473 GND 0.01265f
C7782 VDDH.t547 GND 0.35198f
C7783 VDDH.n474 GND 0.43037f
C7784 VDDH.n475 GND 0.03798f
C7785 VDDH.n476 GND 2.6592f
C7786 VDDH.n477 GND 1.20776f
C7787 VDDH.n478 GND 0.01104f
C7788 VDDH.n479 GND 0.27625f
C7789 VDDH.n480 GND 0.47173f
C7790 VDDH.n481 GND 0.43242f
C7791 VDDH.t548 GND 0.02964f
C7792 VDDH.t549 GND 0.02964f
C7793 VDDH.t546 GND 0.02964f
C7794 VDDH.t550 GND 0.02964f
C7795 VDDH.n482 GND 0.06425f
C7796 VDDH.n483 GND 0.01864f
C7797 VDDH.n484 GND 0.06461f
C7798 VDDH.n485 GND 0.023f
C7799 VDDH.n486 GND 0.05464f
C7800 VDDH.n487 GND 0.09643f
C7801 VDDH.n488 GND 0.07451f
C7802 VDDH.n489 GND 2.82293f
C7803 VDDH.n490 GND 0.09538f
C7804 VDDH.n491 GND 0.05232f
C7805 VDDH.n492 GND 0.03497f
C7806 VDDH.n493 GND 0.02046f
C7807 VDDH.n494 GND 0.06722f
C7808 VDDH.n495 GND 0.06722f
C7809 VDDH.t545 GND 0.35198f
C7810 VDDH.n496 GND 0.43037f
C7811 VDDH.n497 GND 0.03115f
C7812 VDDH.n498 GND 0.06299f
C7813 VDDH.n499 GND 0.09558f
C7814 VDDH.n500 GND 0.01864f
C7815 VDDH.n501 GND 0.09558f
C7816 VDDH.n502 GND 0.0873f
C7817 VDDH.n503 GND 0.03115f
C7818 VDDH.n504 GND 0.02046f
C7819 VDDH.n505 GND 0.03462f
C7820 VDDH.n506 GND 0.04287f
C7821 VDDH.n507 GND 0.09538f
C7822 VDDH.n508 GND 2.33182f
C7823 VDDH.n509 GND 0.08675f
C7824 VDDH.n510 GND 0.10844f
C7825 VDDH.n511 GND 1.40959f
C7826 VDDH.n512 GND 0.04059f
C7827 VDDH.n513 GND 0.023f
C7828 VDDH.n514 GND 0.05219f
C7829 VDDH.n515 GND 0.04941f
C7830 VDDH.n516 GND 0.10201f
C7831 VDDH.n517 GND 0.13946f
C7832 VDDH.n518 GND 0.09672f
C7833 VDDH.n519 GND 0.01972f
C7834 VDDH.n520 GND 0.08077f
C7835 VDDH.t142 GND 0.01757f
C7836 VDDH.t140 GND 0.06625f
C7837 VDDH.t143 GND 0.01757f
C7838 VDDH.t138 GND 0.01757f
C7839 VDDH.t136 GND 0.06625f
C7840 VDDH.t139 GND 0.01757f
C7841 VDDH.n521 GND 0.09993f
C7842 VDDH.n522 GND 0.20917f
C7843 VDDH.t224 GND 0.01757f
C7844 VDDH.t223 GND 0.06625f
C7845 VDDH.t225 GND 0.01757f
C7846 VDDH.t227 GND 0.01757f
C7847 VDDH.t226 GND 0.06625f
C7848 VDDH.t228 GND 0.01757f
C7849 VDDH.n523 GND 0.10074f
C7850 VDDH.n524 GND 0.20914f
C7851 VDDH.n525 GND 0.23325f
C7852 VDDH.n526 GND 0.24973f
C7853 VDDH.n527 GND 0.14151f
C7854 VDDH.n528 GND 0.0896f
C7855 VDDH.n530 GND 0.15863f
C7856 VDDH.n531 GND -0.3593f
C7857 VDDH.n532 GND 0.16184f
C7858 VDDH.n533 GND 0.04274f
C7859 VDDH.n534 GND 1.15562f
C7860 VDDH.n535 GND 0.16707f
C7861 VDDH.n536 GND 0.01273f
C7862 VDDH.n537 GND 0.096f
C7863 VDDH.n538 GND 0.14084f
C7864 VDDH.n539 GND 0.29291f
C7865 VDDH.t149 GND 0.01762f
C7866 VDDH.t147 GND 0.06625f
C7867 VDDH.n540 GND 0.05371f
C7868 VDDH.t118 GND 0.01762f
C7869 VDDH.t117 GND 0.06625f
C7870 VDDH.n541 GND 0.05371f
C7871 VDDH.t119 GND 0.01744f
C7872 VDDH.t148 GND 0.01744f
C7873 VDDH.n542 GND 0.06395f
C7874 VDDH.n543 GND 0.04225f
C7875 VDDH.t161 GND 0.01762f
C7876 VDDH.t159 GND 0.06625f
C7877 VDDH.n544 GND 0.05371f
C7878 VDDH.t121 GND 0.01762f
C7879 VDDH.t120 GND 0.06625f
C7880 VDDH.n545 GND 0.05371f
C7881 VDDH.t122 GND 0.01744f
C7882 VDDH.t160 GND 0.01744f
C7883 VDDH.n546 GND 0.06395f
C7884 VDDH.n547 GND 0.04225f
C7885 VDDH.n548 GND 0.19933f
C7886 VDDH.n549 GND 0.07293f
C7887 VDDH.n550 GND 0.05678f
C7888 VDDH.n551 GND 0.01293f
C7889 VDDH.n552 GND 0.09204f
C7890 VDDH.n554 GND 0.03677f
C7891 VDDH.n555 GND 0.04403f
C7892 VDDH.n556 GND 0.07666f
C7893 VDDH.t126 GND 0.06625f
C7894 VDDH.n557 GND 0.06812f
C7895 VDDH.n558 GND 0.07145f
C7896 VDDH.t127 GND 0.01744f
C7897 VDDH.n559 GND 0.07543f
C7898 VDDH.t134 GND 0.01744f
C7899 VDDH.n560 GND 0.07543f
C7900 VDDH.n561 GND 0.06017f
C7901 VDDH.t133 GND 0.06625f
C7902 VDDH.n562 GND 0.04023f
C7903 VDDH.n563 GND 0.10753f
C7904 VDDH.n564 GND 0.05503f
C7905 VDDH.n565 GND 0.06404f
C7906 VDDH.n566 GND 0.06924f
C7907 VDDH.n567 GND 0.04824f
C7908 VDDH.n568 GND 0.08077f
C7909 VDDH.n569 GND 0.15068f
C7910 VDDH.n570 GND 0.06248f
C7911 VDDH.n571 GND 0.08641f
C7912 VDDH.n572 GND 0.15769f
C7913 VDDH.n573 GND 0.27924f
C7914 VDDH.n574 GND 0.91689f
C7915 VDDH.t539 GND 0.66812f
C7916 VDDH.t273 GND 0.45489f
C7917 VDDH.n575 GND 2.67956f
C7918 VDDH.t83 GND 2.06018f
C7919 VDDH.t457 GND 2.69481f
C7920 VDDH.t141 GND 2.69481f
C7921 VDDH.t137 GND 0.35994f
C7922 VDDH.n576 GND 0.58609f
C7923 VDDH.n577 GND 0.15866f
C7924 VDDH.n579 GND 0.08079f
C7925 VDDH.n580 GND 0.26728f
C7926 VDDH.n581 GND 0.32477f
C7927 VDDH.n582 GND 1.73136f
C7928 VDDH.n583 GND 0.03393f
C7929 VDDH.n584 GND 0.0398f
C7930 VDDH.n585 GND 0.01409f
C7931 VDDH.n586 GND 0.02404f
C7932 VDDH.t419 GND 0.14737f
C7933 VDDH.t69 GND 0.16682f
C7934 VDDH.n588 GND 0.2213f
C7935 VDDH.n589 GND 0.02056f
C7936 VDDH.n590 GND 0.01242f
C7937 VDDH.n591 GND 0.23832f
C7938 VDDH.n592 GND 0.06957f
C7939 VDDH.n593 GND 0.041f
C7940 VDDH.n594 GND 0.02706f
C7941 VDDH.n595 GND 0.0156f
C7942 VDDH.n596 GND 0.02663f
C7943 VDDH.n597 GND 0.0737f
C7944 VDDH.t246 GND 0.12408f
C7945 VDDH.n598 GND 0.20245f
C7946 VDDH.t562 GND 0.13807f
C7947 VDDH.t502 GND 0.15428f
C7948 VDDH.n599 GND 0.10838f
C7949 VDDH.t563 GND 0.07101f
C7950 VDDH.n600 GND 0.10309f
C7951 VDDH.n601 GND 0.01177f
C7952 VDDH.n602 GND 0.02798f
C7953 VDDH.n603 GND 0.29696f
C7954 VDDH.n604 GND 0.81988f
C7955 VDDH.n605 GND 0.04345f
C7956 VDDH.n606 GND 0.17823f
C7957 VDDH.n607 GND 0.02588f
C7958 VDDH.n608 GND 0.05441f
C7959 VDDH.n609 GND 0.0737f
C7960 VDDH.t78 GND 0.15155f
C7961 VDDH.t289 GND 0.14776f
C7962 VDDH.t397 GND 0.15155f
C7963 VDDH.t76 GND 0.15155f
C7964 VDDH.t399 GND 0.15155f
C7965 VDDH.n611 GND 0.17823f
C7966 VDDH.n613 GND 0.04339f
C7967 VDDH.n614 GND 0.04021f
C7968 VDDH.t73 GND 0.14776f
C7969 VDDH.t501 GND 0.15155f
C7970 VDDH.t74 GND 0.15155f
C7971 VDDH.t70 GND 0.15155f
C7972 VDDH.t400 GND 0.15155f
C7973 VDDH.t77 GND 0.15155f
C7974 VDDH.t398 GND 0.13426f
C7975 VDDH.n615 GND 0.11696f
C7976 VDDH.t71 GND 0.13426f
C7977 VDDH.t499 GND 0.15155f
C7978 VDDH.t498 GND 0.15155f
C7979 VDDH.t72 GND 0.15155f
C7980 VDDH.n616 GND 0.03523f
C7981 VDDH.n617 GND 0.0487f
C7982 VDDH.n618 GND 0.18773f
C7983 VDDH.n619 GND 0.06396f
C7984 VDDH.t449 GND 0.14776f
C7985 VDDH.t240 GND 0.15924f
C7986 VDDH.t379 GND 0.15924f
C7987 VDDH.t375 GND 0.15924f
C7988 VDDH.t405 GND 0.11751f
C7989 VDDH.t409 GND 0.11723f
C7990 VDDH.n620 GND 0.06393f
C7991 VDDH.n622 GND 0.02644f
C7992 VDDH.n623 GND 0.04479f
C7993 VDDH.t408 GND 0.15924f
C7994 VDDH.t396 GND 0.15924f
C7995 VDDH.t284 GND 0.15155f
C7996 VDDH.t395 GND 0.13426f
C7997 VDDH.n625 GND 0.11696f
C7998 VDDH.t440 GND 0.13426f
C7999 VDDH.t443 GND 0.15155f
C8000 VDDH.t444 GND 0.15155f
C8001 VDDH.n626 GND 0.04479f
C8002 VDDH.n628 GND 0.1491f
C8003 VDDH.t442 GND 0.13426f
C8004 VDDH.n630 GND 0.11696f
C8005 VDDH.t494 GND 0.13426f
C8006 VDDH.t525 GND 0.15155f
C8007 VDDH.t496 GND 0.14776f
C8008 VDDH.t493 GND 0.15155f
C8009 VDDH.n631 GND 0.02496f
C8010 VDDH.n632 GND 0.02654f
C8011 VDDH.n633 GND 0.04508f
C8012 VDDH.t495 GND 0.15155f
C8013 VDDH.n634 GND 0.04508f
C8014 VDDH.n635 GND 0.01695f
C8015 VDDH.n636 GND 0.02644f
C8016 VDDH.n637 GND 0.02349f
C8017 VDDH.n638 GND 0.04007f
C8018 VDDH.t441 GND 0.15155f
C8019 VDDH.n639 GND 0.04007f
C8020 VDDH.n640 GND 0.02349f
C8021 VDDH.n641 GND 0.03766f
C8022 VDDH.n642 GND 0.04897f
C8023 VDDH.n643 GND 0.08329f
C8024 VDDH.n644 GND 0.04173f
C8025 VDDH.n645 GND 0.03432f
C8026 VDDH.n646 GND 0.08329f
C8027 VDDH.n647 GND 0.04044f
C8028 VDDH.n648 GND 0.03714f
C8029 VDDH.n650 GND 0.03471f
C8030 VDDH.n651 GND 0.04044f
C8031 VDDH.n652 GND 0.07388f
C8032 VDDH.t500 GND 0.15155f
C8033 VDDH.n653 GND 0.07388f
C8034 VDDH.n654 GND 0.0737f
C8035 VDDH.n655 GND 0.07388f
C8036 VDDH.t75 GND 0.15155f
C8037 VDDH.n656 GND 0.07388f
C8038 VDDH.n657 GND 0.04044f
C8039 VDDH.n658 GND 0.03471f
C8040 VDDH.n659 GND 0.13323f
C8041 VDDH.n660 GND 6.28439f
C8042 VDDH.n661 GND 6.83032f
C8043 VDDH.t168 GND 0.01755f
C8044 VDDH.n662 GND 0.05587f
C8045 VDDH.n663 GND 0.11511f
C8046 VDDH.t166 GND 0.06625f
C8047 VDDH.n664 GND 0.02998f
C8048 VDDH.n665 GND 0.05115f
C8049 VDDH.n666 GND 0.06054f
C8050 VDDH.n667 GND 0.02124f
C8051 VDDH.n668 GND 0.0591f
C8052 VDDH.n669 GND 0.02997f
C8053 VDDH.n671 GND 0.06711f
C8054 VDDH.n672 GND 0.61041f
C8055 VDDH.t114 GND 0.88046f
C8056 VDDH.t28 GND 1.07137f
C8057 VDDH.t29 GND 1.00441f
C8058 VDDH.n673 GND 0.53569f
C8059 VDDH.n674 GND 0.07424f
C8060 VDDH.n675 GND 0.02222f
C8061 VDDH.n676 GND 0.02031f
C8062 VDDH.n677 GND 0.02124f
C8063 VDDH.n678 GND 0.05484f
C8064 VDDH.n679 GND 0.06027f
C8065 VDDH.t208 GND 0.06625f
C8066 VDDH.n680 GND 0.09593f
C8067 VDDH.n681 GND 0.04239f
C8068 VDDH.n682 GND 0.02824f
C8069 VDDH.n683 GND 0.03797f
C8070 VDDH.n684 GND 0.07878f
C8071 VDDH.n685 GND 0.03017f
C8072 VDDH.n686 GND 0.04371f
C8073 VDDH.n687 GND 0.0468f
C8074 VDDH.n688 GND 0.0815f
C8075 VDDH.n689 GND 0.09664f
C8076 VDDH.n690 GND 0.06291f
C8077 VDDH.n691 GND 0.02825f
C8078 VDDH.n693 GND 0.02382f
C8079 VDDH.n694 GND 0.05211f
C8080 VDDH.n695 GND 0.05708f
C8081 VDDH.n696 GND 0.04846f
C8082 VDDH.n697 GND 0.02559f
C8083 VDDH.n698 GND 0.16252f
C8084 VDDH.n699 GND 0.06081f
C8085 VDDH.n700 GND 0.05231f
C8086 VDDH.n701 GND 0.01543f
C8087 VDDH.t560 GND 0.01129f
C8088 VDDH.n702 GND 0.03783f
C8089 VDDH.n704 GND 0.05462f
C8090 VDDH.n705 GND 0.04683f
C8091 VDDH.n706 GND 0.03027f
C8092 VDDH.n707 GND 0.05231f
C8093 VDDH.n708 GND 0.04948f
C8094 VDDH.n709 GND 0.05462f
C8095 VDDH.n710 GND 0.04683f
C8096 VDDH.n711 GND 0.03027f
C8097 VDDH.n712 GND 0.08217f
C8098 VDDH.n713 GND 0.47893f
C8099 VDDH.n714 GND 0.07716f
C8100 VDDH.n715 GND 0.07716f
C8101 VDDH.n716 GND 0.04373f
C8102 VDDH.n717 GND 0.01527f
C8103 VDDH.n718 GND 0.02042f
C8104 VDDH.n723 GND 0.01543f
C8105 VDDH.t492 GND 0.01129f
C8106 VDDH.n724 GND 0.03783f
C8107 VDDH.n725 GND 0.01752f
C8108 VDDH.n726 GND 0.01929f
C8109 VDDH.n731 GND 0.21127f
C8110 VDDH.n734 GND 0.02042f
C8111 VDDH.n735 GND 0.12544f
C8112 VDDH.n736 GND 0.35303f
C8113 VDDH.n737 GND 0.01468f
C8114 VDDH.n742 GND 0.0111f
C8115 VDDH.n744 GND 0.05513f
C8116 VDDH.n745 GND 0.04421f
C8117 VDDH.t523 GND 0.04287f
C8118 VDDH.t1 GND 0.01129f
C8119 VDDH.n753 GND 0.01665f
C8120 VDDH.n756 GND 0.04287f
C8121 VDDH.t58 GND 0.16528f
C8122 VDDH.n762 GND 0.05513f
C8123 VDDH.n763 GND 0.0554f
C8124 VDDH.t475 GND 0.01129f
C8125 VDDH.n765 GND 0.03783f
C8126 VDDH.n766 GND 0.09491f
C8127 VDDH.n769 GND 0.08083f
C8128 VDDH.t474 GND 0.04287f
C8129 VDDH.n770 GND 0.01652f
C8130 VDDH.t4 GND 0.04287f
C8131 VDDH.n771 GND 0.04868f
C8132 VDDH.n774 GND 0.04868f
C8133 VDDH.t434 GND 0.04153f
C8134 VDDH.t0 GND 0.01608f
C8135 VDDH.n775 GND 0.04421f
C8136 VDDH.n776 GND 0.08083f
C8137 VDDH.t459 GND 0.13243f
C8138 VDDH.t503 GND 0.13282f
C8139 VDDH.n777 GND 0.08128f
C8140 VDDH.n781 GND 0.01468f
C8141 VDDH.n782 GND 0.0111f
C8142 VDDH.n783 GND 0.03783f
C8143 VDDH.n785 GND 0.04069f
C8144 VDDH.n788 GND 0.0554f
C8145 VDDH.t524 GND 0.01129f
C8146 VDDH.n790 GND 0.03783f
C8147 VDDH.n791 GND 0.0111f
C8148 VDDH.n792 GND 0.01468f
C8149 VDDH.n795 GND 0.01652f
C8150 VDDH.t426 GND 0.04287f
C8151 VDDH.n796 GND 0.04868f
C8152 VDDH.n797 GND 0.04287f
C8153 VDDH.t371 GND 0.01608f
C8154 VDDH.t470 GND 0.04153f
C8155 VDDH.n798 GND 0.04868f
C8156 VDDH.n801 GND 0.01665f
C8157 VDDH.n802 GND 0.01468f
C8158 VDDH.n803 GND 0.0111f
C8159 VDDH.t372 GND 0.01129f
C8160 VDDH.n804 GND 0.03783f
C8161 VDDH.n809 GND 0.08128f
C8162 VDDH.t373 GND 0.13282f
C8163 VDDH.t351 GND 0.13243f
C8164 VDDH.n810 GND 0.08083f
C8165 VDDH.t406 GND 0.04287f
C8166 VDDH.n811 GND 0.01652f
C8167 VDDH.t24 GND 0.04287f
C8168 VDDH.n812 GND 0.04868f
C8169 VDDH.t18 GND 0.04153f
C8170 VDDH.n815 GND 0.01665f
C8171 VDDH.t353 GND 0.01129f
C8172 VDDH.n818 GND 0.03783f
C8173 VDDH.n819 GND 0.0111f
C8174 VDDH.n820 GND 0.01468f
C8175 VDDH.t352 GND 0.01608f
C8176 VDDH.n822 GND 0.08083f
C8177 VDDH.t38 GND 0.13243f
C8178 VDDH.t561 GND 0.13282f
C8179 VDDH.n823 GND 0.08128f
C8180 VDDH.n824 GND 0.04421f
C8181 VDDH.n827 GND 0.04868f
C8182 VDDH.n828 GND 0.04287f
C8183 VDDH.n829 GND 0.05513f
C8184 VDDH.n830 GND 0.0554f
C8185 VDDH.t407 GND 0.01129f
C8186 VDDH.n831 GND 0.03783f
C8187 VDDH.n837 GND 0.04069f
C8188 VDDH.n838 GND 0.31817f
C8189 VDDH.n839 GND 0.31817f
C8190 VDDH.n840 GND 0.31817f
C8191 VDDH.n841 GND 0.31817f
C8192 VDDH.n842 GND 0.04069f
C8193 VDDH.n845 GND 0.0554f
C8194 VDDH.t355 GND 0.01129f
C8195 VDDH.n847 GND 0.03783f
C8196 VDDH.n848 GND 0.0111f
C8197 VDDH.n849 GND 0.01468f
C8198 VDDH.n852 GND 0.01652f
C8199 VDDH.t12 GND 0.04287f
C8200 VDDH.n853 GND 0.04868f
C8201 VDDH.n854 GND 0.04287f
C8202 VDDH.t348 GND 0.01608f
C8203 VDDH.t6 GND 0.04153f
C8204 VDDH.n855 GND 0.04868f
C8205 VDDH.n858 GND 0.01665f
C8206 VDDH.n859 GND 0.01468f
C8207 VDDH.n860 GND 0.0111f
C8208 VDDH.t349 GND 0.01129f
C8209 VDDH.n861 GND 0.03783f
C8210 VDDH.n866 GND 0.08128f
C8211 VDDH.t339 GND 0.13282f
C8212 VDDH.t451 GND 0.13243f
C8213 VDDH.t2 GND 0.04287f
C8214 VDDH.n867 GND 0.01652f
C8215 VDDH.t309 GND 0.04287f
C8216 VDDH.n868 GND 0.08083f
C8217 VDDH.n871 GND 0.04069f
C8218 VDDH.n872 GND 0.01468f
C8219 VDDH.n873 GND 0.0111f
C8220 VDDH.t310 GND 0.01129f
C8221 VDDH.n874 GND 0.03783f
C8222 VDDH.t328 GND 0.01608f
C8223 VDDH.n879 GND 0.04421f
C8224 VDDH.t374 GND 0.13282f
C8225 VDDH.n880 GND 0.08128f
C8226 VDDH.t329 GND 0.01129f
C8227 VDDH.n885 GND 0.03783f
C8228 VDDH.n886 GND 0.0111f
C8229 VDDH.n887 GND 0.01468f
C8230 VDDH.n888 GND 0.01665f
C8231 VDDH.n891 GND 0.04868f
C8232 VDDH.n892 GND 0.04287f
C8233 VDDH.n893 GND 0.05513f
C8234 VDDH.n894 GND 0.05513f
C8235 VDDH.n895 GND 0.0554f
C8236 VDDH.t68 GND 0.01129f
C8237 VDDH.n897 GND 0.03783f
C8238 VDDH.n898 GND 0.0111f
C8239 VDDH.n899 GND 0.01468f
C8240 VDDH.n900 GND 0.04069f
C8241 VDDH.n903 GND 0.08083f
C8242 VDDH.t67 GND 0.04287f
C8243 VDDH.n904 GND 0.01652f
C8244 VDDH.t472 GND 0.04287f
C8245 VDDH.n905 GND 0.04868f
C8246 VDDH.n908 GND 0.04868f
C8247 VDDH.t26 GND 0.04153f
C8248 VDDH.t535 GND 0.01608f
C8249 VDDH.n909 GND 0.04421f
C8250 VDDH.t244 GND 0.13282f
C8251 VDDH.n910 GND 0.08128f
C8252 VDDH.n914 GND 0.01468f
C8253 VDDH.n915 GND 0.0111f
C8254 VDDH.n916 GND 0.03783f
C8255 VDDH.n920 GND 0.0554f
C8256 VDDH.t529 GND 0.01129f
C8257 VDDH.n922 GND 0.03783f
C8258 VDDH.n923 GND 0.0111f
C8259 VDDH.n924 GND 0.01468f
C8260 VDDH.n925 GND 0.04069f
C8261 VDDH.n928 GND 0.08083f
C8262 VDDH.t528 GND 0.04287f
C8263 VDDH.n929 GND 0.01652f
C8264 VDDH.t20 GND 0.04287f
C8265 VDDH.n930 GND 0.04868f
C8266 VDDH.n933 GND 0.04868f
C8267 VDDH.t14 GND 0.04153f
C8268 VDDH.t79 GND 0.01608f
C8269 VDDH.n934 GND 0.04421f
C8270 VDDH.t575 GND 0.13292f
C8271 VDDH.t521 GND 0.1365f
C8272 VDDH.n935 GND 0.08128f
C8273 VDDH.n939 GND 0.01468f
C8274 VDDH.n940 GND 0.0111f
C8275 VDDH.n941 GND 0.03783f
C8276 VDDH.n943 GND 0.31817f
C8277 VDDH.t517 GND 0.01129f
C8278 VDDH.n952 GND 0.06535f
C8279 VDDH.n953 GND 0.0111f
C8280 VDDH.n954 GND 0.03783f
C8281 VDDH.n958 GND 0.0111f
C8282 VDDH.t505 GND 0.01129f
C8283 VDDH.n959 GND 0.03783f
C8284 VDDH.n966 GND 0.05722f
C8285 VDDH.n967 GND 0.31022f
C8286 VDDH.n968 GND 0.31817f
C8287 VDDH.t574 GND 0.01129f
C8288 VDDH.n970 GND 0.03783f
C8289 VDDH.n971 GND 0.0111f
C8290 VDDH.n972 GND 0.06535f
C8291 VDDH.n973 GND 0.05513f
C8292 VDDH.n974 GND 0.05479f
C8293 VDDH.t432 GND 0.08077f
C8294 VDDH.t497 GND 0.13684f
C8295 VDDH.t515 GND 0.13684f
C8296 VDDH.t22 GND 0.08077f
C8297 VDDH.n975 GND 0.05479f
C8298 VDDH.t468 GND 0.08077f
C8299 VDDH.t331 GND 0.13684f
C8300 VDDH.t506 GND 0.13684f
C8301 VDDH.t10 GND 0.08077f
C8302 VDDH.t334 GND 0.13684f
C8303 VDDH.t514 GND 0.13684f
C8304 VDDH.t8 GND 0.08077f
C8305 VDDH.n976 GND 0.05479f
C8306 VDDH.n977 GND 0.05513f
C8307 VDDH.n978 GND 0.05513f
C8308 VDDH.t526 GND 0.16945f
C8309 VDDH.t430 GND 0.08077f
C8310 VDDH.n979 GND 0.05479f
C8311 VDDH.t332 GND 0.12385f
C8312 VDDH.n980 GND 0.04286f
C8313 VDDH.n982 GND 0.0111f
C8314 VDDH.t333 GND 0.01129f
C8315 VDDH.n983 GND 0.03783f
C8316 VDDH.n989 GND 0.05722f
C8317 VDDH.n990 GND 0.71449f
C8318 VDDH.n991 GND 14.417f
C8319 VDDH.t285 GND 0.03754f
C8320 VDDH.n992 GND 0.78306f
C8321 VDDH.n993 GND 9.99452f
C8322 VDDH.n994 GND 0.02719f
C8323 VDDH.n995 GND 0.17097f
C8324 VDDH.n996 GND 0.03217f
C8325 VDDH.n997 GND 0.02711f
C8326 VDDH.n998 GND 0.02445f
C8327 VDDH.n999 GND 0.04666f
C8328 VDDH.n1000 GND 0.17097f
C8329 VDDH.n1001 GND 0.17097f
C8330 VDDH.t488 GND 0.14776f
C8331 VDDH.t486 GND 0.15155f
C8332 VDDH.t484 GND 0.15155f
C8333 VDDH.t489 GND 0.11367f
C8334 VDDH.t481 GND 0.14776f
C8335 VDDH.t482 GND 0.15155f
C8336 VDDH.t485 GND 0.15155f
C8337 VDDH.t487 GND 0.11367f
C8338 VDDH.n1003 GND 0.03514f
C8339 VDDH.n1004 GND 0.02257f
C8340 VDDH.n1005 GND 0.17097f
C8341 VDDH.n1006 GND 0.17097f
C8342 VDDH.t531 GND 0.14776f
C8343 VDDH.t322 GND 0.15155f
C8344 VDDH.t424 GND 0.15155f
C8345 VDDH.t534 GND 0.11367f
C8346 VDDH.n1008 GND 0.04773f
C8347 VDDH.n1009 GND 0.02664f
C8348 VDDH.n1010 GND 0.0321f
C8349 VDDH.n1011 GND 0.17097f
C8350 VDDH.n1012 GND 0.17097f
C8351 VDDH.t532 GND 0.14776f
C8352 VDDH.t421 GND 0.15155f
C8353 VDDH.t422 GND 0.15155f
C8354 VDDH.t423 GND 0.11367f
C8355 VDDH.n1015 GND 0.03491f
C8356 VDDH.n1016 GND 0.17097f
C8357 VDDH.n1017 GND 0.17097f
C8358 VDDH.t341 GND 0.14776f
C8359 VDDH.t35 GND 0.15155f
C8360 VDDH.t39 GND 0.15155f
C8361 VDDH.t255 GND 0.11367f
C8362 VDDH.t357 GND 0.14776f
C8363 VDDH.t254 GND 0.15155f
C8364 VDDH.t253 GND 0.15155f
C8365 VDDH.t518 GND 0.11367f
C8366 VDDH.n1018 GND 0.04773f
C8367 VDDH.n1021 GND 0.0501f
C8368 VDDH.n1023 GND 0.043f
C8369 VDDH.n1024 GND 0.17097f
C8370 VDDH.n1025 GND 0.17097f
C8371 VDDH.t63 GND 0.14776f
C8372 VDDH.t460 GND 0.15155f
C8373 VDDH.t461 GND 0.15155f
C8374 VDDH.t60 GND 0.11367f
C8375 VDDH.t61 GND 0.14776f
C8376 VDDH.t59 GND 0.15155f
C8377 VDDH.t579 GND 0.15155f
C8378 VDDH.t465 GND 0.11367f
C8379 VDDH.n1026 GND 0.03514f
C8380 VDDH.n1028 GND 0.07066f
C8381 VDDH.n1030 GND 0.17097f
C8382 VDDH.n1031 GND 0.17097f
C8383 VDDH.t342 GND 0.14776f
C8384 VDDH.t377 GND 0.15155f
C8385 VDDH.t344 GND 0.15155f
C8386 VDDH.t343 GND 0.11367f
C8387 VDDH.t414 GND 0.14776f
C8388 VDDH.t376 GND 0.15155f
C8389 VDDH.t416 GND 0.15155f
C8390 VDDH.t415 GND 0.11367f
C8391 VDDH.n1032 GND 0.05708f
C8392 VDDH.n1033 GND 0.03826f
C8393 VDDH.n1034 GND 0.03626f
C8394 VDDH.n1035 GND 0.07159f
C8395 VDDH.n1036 GND 0.0362f
C8396 VDDH.n1037 GND 0.07159f
C8397 VDDH.n1038 GND 0.02445f
C8398 VDDH.n1039 GND 0.17097f
C8399 VDDH.t243 GND 0.14776f
C8400 VDDH.t450 GND 0.15155f
C8401 VDDH.t448 GND 0.15155f
C8402 VDDH.t242 GND 0.11367f
C8403 VDDH.n1040 GND 0.07578f
C8404 VDDH.t259 GND 0.11367f
C8405 VDDH.t260 GND 0.15155f
C8406 VDDH.t241 GND 0.15155f
C8407 VDDH.t258 GND 0.14776f
C8408 VDDH.n1041 GND 0.17097f
C8409 VDDH.n1043 GND 0.04195f
C8410 VDDH.n1044 GND 0.02776f
C8411 VDDH.n1045 GND 0.04502f
C8412 VDDH.n1046 GND 0.21817f
C8413 VDDH.n1047 GND 0.21817f
C8414 VDDH.t311 GND 0.14776f
C8415 VDDH.t307 GND 0.15155f
C8416 VDDH.t378 GND 0.15155f
C8417 VDDH.t308 GND 0.15924f
C8418 VDDH.t250 GND 0.15924f
C8419 VDDH.t248 GND 0.15155f
C8420 VDDH.t247 GND 0.1252f
C8421 VDDH.t530 GND 0.15544f
C8422 VDDH.t312 GND 0.16693f
C8423 VDDH.t330 GND 0.15924f
C8424 VDDH.t350 GND 0.15924f
C8425 VDDH.t522 GND 0.15924f
C8426 VDDH.t458 GND 0.15924f
C8427 VDDH.t249 GND 0.10982f
C8428 VDDH.n1048 GND 0.03826f
C8429 VDDH.n1049 GND 0.06976f
C8430 VDDH.n1050 GND 0.11847f
C8431 VDDH.n1051 GND 0.07578f
C8432 VDDH.n1052 GND 0.11847f
C8433 VDDH.n1053 GND 0.06378f
C8434 VDDH.n1054 GND 0.04502f
C8435 VDDH.n1055 GND 0.01773f
C8436 VDDH.n1056 GND 0.03081f
C8437 VDDH.n1057 GND 0.02478f
C8438 VDDH.n1058 GND 0.07159f
C8439 VDDH.n1059 GND 0.07578f
C8440 VDDH.n1060 GND 0.07159f
C8441 VDDH.n1061 GND 0.0362f
C8442 VDDH.n1062 GND 0.07066f
C8443 VDDH.n1063 GND 0.02625f
C8444 VDDH.n1064 GND 0.03221f
C8445 VDDH.n1065 GND 0.17097f
C8446 VDDH.n1067 GND 0.17097f
C8447 VDDH.t37 GND 0.14776f
C8448 VDDH.t340 GND 0.15155f
C8449 VDDH.t519 GND 0.15155f
C8450 VDDH.t36 GND 0.11367f
C8451 VDDH.n1068 GND 0.0362f
C8452 VDDH.n1069 GND 0.07159f
C8453 VDDH.t40 GND 0.14776f
C8454 VDDH.t520 GND 0.15155f
C8455 VDDH.t356 GND 0.15155f
C8456 VDDH.t41 GND 0.11367f
C8457 VDDH.n1070 GND 0.07578f
C8458 VDDH.n1071 GND 0.07159f
C8459 VDDH.n1072 GND 0.02487f
C8460 VDDH.n1073 GND 0.03167f
C8461 VDDH.n1074 GND 0.02932f
C8462 VDDH.n1075 GND 0.02782f
C8463 VDDH.n1076 GND 0.03167f
C8464 VDDH.n1077 GND 0.0294f
C8465 VDDH.n1078 GND 0.07159f
C8466 VDDH.n1079 GND 0.07578f
C8467 VDDH.n1080 GND 0.07159f
C8468 VDDH.n1081 GND 0.03922f
C8469 VDDH.n1082 GND 0.0501f
C8470 VDDH.n1083 GND 0.03517f
C8471 VDDH.n1084 GND 0.17097f
C8472 VDDH.n1085 GND 0.17097f
C8473 VDDH.t464 GND 0.14776f
C8474 VDDH.t65 GND 0.15155f
C8475 VDDH.t62 GND 0.15155f
C8476 VDDH.t463 GND 0.11367f
C8477 VDDH.n1086 GND 0.03467f
C8478 VDDH.n1087 GND 0.03491f
C8479 VDDH.n1088 GND 0.03922f
C8480 VDDH.n1089 GND 0.07159f
C8481 VDDH.t576 GND 0.14776f
C8482 VDDH.t462 GND 0.15155f
C8483 VDDH.t578 GND 0.15155f
C8484 VDDH.t577 GND 0.11367f
C8485 VDDH.n1090 GND 0.07578f
C8486 VDDH.n1091 GND 0.07159f
C8487 VDDH.n1092 GND 0.01505f
C8488 VDDH.n1093 GND 0.0321f
C8489 VDDH.n1094 GND 0.02814f
C8490 VDDH.n1095 GND 0.02782f
C8491 VDDH.n1096 GND 0.0321f
C8492 VDDH.n1097 GND 0.02761f
C8493 VDDH.n1098 GND 0.0321f
C8494 VDDH.n1099 GND 0.01268f
C8495 VDDH.n1100 GND 0.07159f
C8496 VDDH.n1101 GND 0.07578f
C8497 VDDH.n1102 GND 0.07159f
C8498 VDDH.n1103 GND 0.0362f
C8499 VDDH.n1104 GND 0.03319f
C8500 VDDH.n1105 GND 0.03319f
C8501 VDDH.n1107 GND 0.03217f
C8502 VDDH.n1108 GND 0.0362f
C8503 VDDH.n1109 GND 0.07159f
C8504 VDDH.t533 GND 0.14776f
C8505 VDDH.t447 GND 0.15155f
C8506 VDDH.t445 GND 0.15155f
C8507 VDDH.t420 GND 0.11367f
C8508 VDDH.n1110 GND 0.07578f
C8509 VDDH.n1111 GND 0.07159f
C8510 VDDH.n1112 GND 0.01161f
C8511 VDDH.n1113 GND 0.0321f
C8512 VDDH.n1114 GND 0.04666f
C8513 VDDH.n1115 GND 0.0362f
C8514 VDDH.n1116 GND 0.07159f
C8515 VDDH.t323 GND 0.14776f
C8516 VDDH.t321 GND 0.15155f
C8517 VDDH.t446 GND 0.15155f
C8518 VDDH.t324 GND 0.11367f
C8519 VDDH.n1117 GND 0.07578f
C8520 VDDH.n1118 GND 0.07159f
C8521 VDDH.n1119 GND 0.03468f
C8522 VDDH.n1120 GND 0.03167f
C8523 VDDH.n1121 GND 0.01607f
C8524 VDDH.n1123 GND 0.03266f
C8525 VDDH.n1124 GND 0.03922f
C8526 VDDH.n1125 GND 0.07159f
C8527 VDDH.n1126 GND 0.07578f
C8528 VDDH.n1127 GND 0.07159f
C8529 VDDH.n1128 GND 0.0362f
C8530 VDDH.n1129 GND 0.02636f
C8531 VDDH.n1130 GND 0.02731f
C8532 VDDH.n1131 GND 0.0261f
C8533 VDDH.n1133 GND 0.17097f
C8534 VDDH.t483 GND 0.14776f
C8535 VDDH.t476 GND 0.15155f
C8536 VDDH.t480 GND 0.15155f
C8537 VDDH.t479 GND 0.11367f
C8538 VDDH.t478 GND 0.14776f
C8539 VDDH.t490 GND 0.15155f
C8540 VDDH.t491 GND 0.15155f
C8541 VDDH.t477 GND 0.11367f
C8542 VDDH.n1134 GND 0.07159f
C8543 VDDH.n1135 GND 0.07578f
C8544 VDDH.n1136 GND 0.07159f
C8545 VDDH.n1137 GND 0.03922f
C8546 VDDH.n1138 GND 0.14057f
C8547 VDDH.n1139 GND 6.48486f
C8548 a_14331_6250.t4 GND 0.0968f
C8549 a_14331_6250.t3 GND 0.09483f
C8550 a_14331_6250.t2 GND 0.07529f
C8551 a_14331_6250.n0 GND 4.30036f
C8552 a_14331_6250.t1 GND 0.1106f
C8553 a_14331_6250.n1 GND 4.73412f
C8554 a_14331_6250.n2 GND 5.41272f
C8555 a_14331_6250.t0 GND 0.07529f
C8556 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y GND 0.52167f
C8557 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t0 GND 0.08583f
C8558 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n0 GND 0.03519f
C8559 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n1 GND 0.07575f
C8560 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n2 GND 0.05029f
C8561 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t1 GND 0.08222f
C8562 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n3 GND 0.01039f
C8563 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t10 GND 0.1705f
C8564 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t17 GND 0.16969f
C8565 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n4 GND 0.53197f
C8566 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t13 GND 0.16969f
C8567 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n5 GND 0.26639f
C8568 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t14 GND 0.16969f
C8569 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n6 GND 0.22129f
C8570 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t15 GND 0.1705f
C8571 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t3 GND 0.16969f
C8572 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n7 GND 0.53197f
C8573 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t2 GND 0.16969f
C8574 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n8 GND 0.26639f
C8575 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t16 GND 0.16969f
C8576 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n9 GND 0.22129f
C8577 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n10 GND 0.65118f
C8578 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t12 GND 0.16969f
C8579 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n11 GND 1.05719f
C8580 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t11 GND 0.16969f
C8581 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n12 GND 0.26639f
C8582 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t8 GND 0.16969f
C8583 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n13 GND 0.26639f
C8584 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t6 GND 0.16969f
C8585 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n14 GND 0.26639f
C8586 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t4 GND 0.16969f
C8587 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n15 GND 0.26639f
C8588 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t9 GND 0.16969f
C8589 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n16 GND 0.26639f
C8590 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t7 GND 0.16969f
C8591 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n17 GND 0.26639f
C8592 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.t5 GND 0.16969f
C8593 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n18 GND 14.7741f
C8594 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec2b[0] GND 0.1379f
C8595 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n19 GND 12.494f
C8596 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0.n20 GND 0.07003f
C8597 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t6 GND 0.16908f
C8598 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t2 GND 0.16823f
C8599 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n0 GND 0.50612f
C8600 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t9 GND 0.16908f
C8601 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t3 GND 0.16823f
C8602 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n1 GND 0.54795f
C8603 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n2 GND 0.13418f
C8604 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t4 GND 0.16629f
C8605 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n3 GND 15.1749f
C8606 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t0 GND 0.13933f
C8607 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t1 GND 0.11828f
C8608 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n4 GND 1.15353f
C8609 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t5 GND 0.55227f
C8610 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t7 GND 0.54999f
C8611 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n5 GND 0.91171f
C8612 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].t8 GND 0.54999f
C8613 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n6 GND 0.47041f
C8614 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0].n7 GND 0.86048f
C8615 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t0 GND 0.05358f
C8616 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t12 GND 0.85572f
C8617 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n0 GND 0.12606f
C8618 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t1 GND 0.08482f
C8619 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n1 GND 0.05712f
C8620 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t3 GND 0.08482f
C8621 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t2 GND 0.01718f
C8622 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n2 GND 0.1007f
C8623 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t4 GND 0.01718f
C8624 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n3 GND 0.13843f
C8625 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n4 GND 0.05663f
C8626 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t18 GND 0.12218f
C8627 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n5 GND 0.07605f
C8628 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t9 GND 0.12218f
C8629 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n6 GND 0.0851f
C8630 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t17 GND 0.12218f
C8631 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n7 GND 0.0851f
C8632 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t8 GND 0.12218f
C8633 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n8 GND 0.05779f
C8634 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t14 GND 0.12218f
C8635 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n9 GND 0.06025f
C8636 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t7 GND 0.12218f
C8637 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n10 GND 0.0851f
C8638 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t13 GND 0.12218f
C8639 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n11 GND 0.0851f
C8640 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t10 GND 0.12218f
C8641 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n12 GND 0.08168f
C8642 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t6 GND 0.12218f
C8643 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n13 GND 0.06025f
C8644 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t16 GND 0.12218f
C8645 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n14 GND 0.0851f
C8646 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t15 GND 0.12218f
C8647 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n15 GND 0.0851f
C8648 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t11 GND 0.12218f
C8649 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n16 GND 0.08168f
C8650 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n17 GND 0.27847f
C8651 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n18 GND 0.75769f
C8652 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n19 GND 0.13016f
C8653 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n20 GND 0.39284f
C8654 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n21 GND 0.26288f
C8655 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t5 GND 0.05626f
C8656 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n22 GND 0.23923f
C8657 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.t1 GND 0.04754f
C8658 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.t0 GND 0.14298f
C8659 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.t2 GND 0.14263f
C8660 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9.n0 GND 2.55569f
C8661 a_30056_7686.t2 GND 0.0855f
C8662 a_30056_7686.t3 GND 0.14007f
C8663 a_30056_7686.t1 GND 0.07805f
C8664 a_30056_7686.n0 GND 5.65951f
C8665 a_30056_7686.t4 GND 0.07805f
C8666 a_30056_7686.n1 GND 2.99489f
C8667 a_30056_7686.n2 GND 3.75935f
C8668 a_30056_7686.t0 GND 0.10458f
C8669 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t0 GND 0.09748f
C8670 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t1 GND 0.08275f
C8671 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n0 GND 0.80704f
C8672 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t7 GND 0.38639f
C8673 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t19 GND 0.38479f
C8674 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n1 GND 0.63787f
C8675 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t11 GND 0.38479f
C8676 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n2 GND 0.32912f
C8677 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n3 GND 0.60202f
C8678 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t22 GND 0.11796f
C8679 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t6 GND 0.11634f
C8680 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n4 GND 3.73702f
C8681 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t5 GND 0.1183f
C8682 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t8 GND 0.1177f
C8683 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n5 GND 0.38336f
C8684 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t10 GND 0.1177f
C8685 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n6 GND 0.19198f
C8686 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t4 GND 0.1177f
C8687 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n7 GND 0.1585f
C8688 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t14 GND 0.1183f
C8689 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t12 GND 0.1177f
C8690 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n8 GND 0.38336f
C8691 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t9 GND 0.1177f
C8692 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n9 GND 0.19198f
C8693 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t15 GND 0.1177f
C8694 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n10 GND 0.1585f
C8695 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n11 GND 0.20637f
C8696 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t18 GND 0.1183f
C8697 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t21 GND 0.1177f
C8698 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n12 GND 0.38336f
C8699 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t16 GND 0.1177f
C8700 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n13 GND 0.19198f
C8701 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t17 GND 0.1177f
C8702 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n14 GND 0.19198f
C8703 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t20 GND 0.1177f
C8704 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n15 GND 0.19198f
C8705 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t3 GND 0.1177f
C8706 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n16 GND 0.19198f
C8707 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t2 GND 0.1177f
C8708 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n17 GND 0.19198f
C8709 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t23 GND 0.1177f
C8710 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n18 GND 0.15678f
C8711 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n19 GND 3.06972f
C8712 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n20 GND 10.845f
C8713 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t13 GND 0.21873f
C8714 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].t24 GND 0.12134f
C8715 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n21 GND 0.1906f
C8716 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n22 GND 0.03327f
C8717 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0].n23 GND 0.26302f
C8718 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t14 GND 0.04436f
C8719 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t1 GND 0.04436f
C8720 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t5 GND 0.04436f
C8721 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t3 GND 0.01245f
C8722 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t6 GND 0.01245f
C8723 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n0 GND 0.02734f
C8724 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t4 GND 0.04436f
C8725 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t20 GND 0.04436f
C8726 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t22 GND 0.01245f
C8727 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t23 GND 0.01245f
C8728 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n1 GND 0.02734f
C8729 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t21 GND 0.04436f
C8730 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t7 GND 0.27187f
C8731 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t8 GND 0.22818f
C8732 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t13 GND 0.30968f
C8733 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n2 GND 1.11186f
C8734 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t12 GND 0.27344f
C8735 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n3 GND 0.70969f
C8736 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n4 GND 1.26622f
C8737 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t42 GND 0.8241f
C8738 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t41 GND 0.93054f
C8739 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t35 GND 0.68684f
C8740 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n5 GND 0.8925f
C8741 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t29 GND 0.68684f
C8742 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n6 GND 0.53851f
C8743 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n7 GND 0.48945f
C8744 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t39 GND 0.8241f
C8745 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t38 GND 0.93054f
C8746 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t33 GND 0.68684f
C8747 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n8 GND 0.8925f
C8748 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t26 GND 0.68684f
C8749 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n9 GND 0.53851f
C8750 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n10 GND 0.46043f
C8751 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n11 GND 0.61675f
C8752 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t31 GND 0.8241f
C8753 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t30 GND 0.93054f
C8754 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t43 GND 0.68684f
C8755 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n12 GND 0.8925f
C8756 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t36 GND 0.68684f
C8757 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n13 GND 0.53851f
C8758 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n14 GND 0.46043f
C8759 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n15 GND 0.34287f
C8760 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t25 GND 0.8241f
C8761 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t24 GND 0.93054f
C8762 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t37 GND 0.68684f
C8763 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n16 GND 0.8925f
C8764 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t32 GND 0.68684f
C8765 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n17 GND 0.53851f
C8766 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n18 GND 0.48929f
C8767 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t28 GND 0.8241f
C8768 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t27 GND 0.93054f
C8769 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t40 GND 0.68684f
C8770 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n19 GND 0.8925f
C8771 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t34 GND 0.68684f
C8772 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n20 GND 0.53851f
C8773 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n21 GND 0.46043f
C8774 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n22 GND 0.48153f
C8775 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n23 GND 1.98328f
C8776 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n24 GND 1.84928f
C8777 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n25 GND 0.31773f
C8778 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n26 GND 0.19617f
C8779 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n27 GND 0.26296f
C8780 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n28 GND 0.20871f
C8781 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n29 GND 0.17232f
C8782 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n30 GND 0.19617f
C8783 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n31 GND 0.26296f
C8784 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n32 GND 0.20871f
C8785 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n33 GND 0.17232f
C8786 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n34 GND 0.19617f
C8787 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t15 GND 0.01245f
C8788 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t0 GND 0.01245f
C8789 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n35 GND 0.02734f
C8790 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n36 GND 0.26297f
C8791 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n37 GND 0.2087f
C8792 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t11 GND 0.01245f
C8793 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t9 GND 0.01245f
C8794 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n38 GND 0.02734f
C8795 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t2 GND 0.04436f
C8796 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t16 GND 0.01245f
C8797 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t19 GND 0.01245f
C8798 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n39 GND 0.02734f
C8799 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t17 GND 0.04624f
C8800 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n40 GND 0.42562f
C8801 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t18 GND 0.04436f
C8802 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n41 GND 0.19617f
C8803 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n42 GND 0.17232f
C8804 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n43 GND 0.2087f
C8805 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n44 GND 0.26297f
C8806 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t10 GND 0.04436f
C8807 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n45 GND 0.19617f
C8808 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n46 GND 0.17232f
C8809 a_6778_12595.t2 GND 0.01193f
C8810 a_6778_12595.t7 GND 0.01193f
C8811 a_6778_12595.t4 GND 0.01193f
C8812 a_6778_12595.n0 GND 0.02768f
C8813 a_6778_12595.t3 GND 0.01193f
C8814 a_6778_12595.t8 GND 0.01193f
C8815 a_6778_12595.n1 GND 0.02768f
C8816 a_6778_12595.n2 GND 0.2036f
C8817 a_6778_12595.t6 GND 0.05399f
C8818 a_6778_12595.t9 GND 0.04624f
C8819 a_6778_12595.n3 GND 2.06772f
C8820 a_6778_12595.n4 GND 0.11865f
C8821 a_6778_12595.t1 GND 0.01193f
C8822 a_6778_12595.t5 GND 0.01193f
C8823 a_6778_12595.n5 GND 0.02768f
C8824 a_6778_12595.n6 GND 0.2036f
C8825 a_6778_12595.n7 GND 0.02768f
C8826 a_6778_12595.t0 GND 0.01193f
C8827 top_DAC_0/top_final_switch_0.VOUT[1].t2 GND 0.01026f
C8828 top_DAC_0/top_final_switch_0.VOUT[1].t3 GND 0.01026f
C8829 top_DAC_0/top_final_switch_0.VOUT[1].n0 GND 0.02336f
C8830 top_DAC_0/top_final_switch_0.VOUT[1].t0 GND 0.01026f
C8831 top_DAC_0/top_final_switch_0.VOUT[1].t1 GND 0.01026f
C8832 top_DAC_0/top_final_switch_0.VOUT[1].n1 GND 0.02438f
C8833 top_DAC_0/top_final_switch_0.VOUT[1].n2 GND 1.39086f
C8834 top_DAC_0/top_final_switch_0.VOUT[1].t9 GND 0.95454f
C8835 top_DAC_0/top_final_switch_0.VOUT[1].t7 GND 0.9486f
C8836 top_DAC_0/top_final_switch_0.VOUT[1].n3 GND 1.58277f
C8837 top_DAC_0/top_final_switch_0.VOUT[1].t5 GND 0.94923f
C8838 top_DAC_0/top_final_switch_0.VOUT[1].t11 GND 0.94749f
C8839 top_DAC_0/top_final_switch_0.VOUT[1].n4 GND 1.22217f
C8840 top_DAC_0/top_final_switch_0.VOUT[1].n5 GND 0.86462f
C8841 top_DAC_0/top_final_switch_0.VOUT[1].t4 GND 0.38998f
C8842 top_DAC_0/top_final_switch_0.VOUT[1].t10 GND 0.38811f
C8843 top_DAC_0/top_final_switch_0.VOUT[1].n6 GND 1.03073f
C8844 top_DAC_0/top_final_switch_0.VOUT[1].t8 GND 0.39642f
C8845 top_DAC_0/top_final_switch_0.VOUT[1].t6 GND 0.38972f
C8846 top_DAC_0/top_final_switch_0.VOUT[1].n7 GND 1.1481f
C8847 top_DAC_0/top_final_switch_0.VOUT[1].n8 GND 0.5353f
C8848 top_DAC_0/top_final_switch_0.VOUT[1].n9 GND 1.75445f
C8849 top_DAC_0/top_final_switch_0.VOUT[1].n10 GND 0.25027f
C8850 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t2 GND 0.04535f
C8851 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t3 GND 0.04535f
C8852 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n0 GND 0.09959f
C8853 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n1 GND 0.04296f
C8854 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t7 GND 0.07054f
C8855 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t12 GND 0.04157f
C8856 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t13 GND 0.07054f
C8857 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t8 GND 0.04157f
C8858 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n2 GND 0.11836f
C8859 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n3 GND 0.17559f
C8860 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n4 GND 0.05295f
C8861 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t10 GND 0.04679f
C8862 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t6 GND 0.07497f
C8863 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n5 GND 0.14751f
C8864 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n6 GND 0.23906f
C8865 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n7 GND 1.13361f
C8866 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t11 GND 0.04687f
C8867 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t9 GND 0.07507f
C8868 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n8 GND 0.14345f
C8869 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n9 GND 0.63171f
C8870 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n10 GND 1.9824f
C8871 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t4 GND 0.04689f
C8872 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t5 GND 0.07509f
C8873 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n11 GND 0.14293f
C8874 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n12 GND 0.27598f
C8875 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n13 GND 12.0537f
C8876 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n14 GND 9.98745f
C8877 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n15 GND 0.03244f
C8878 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t0 GND 0.02948f
C8879 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t1 GND 0.02948f
C8880 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n16 GND 0.07028f
C8881 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n17 GND 0.13808f
C8882 VDD.n0 GND 1.73611f
C8883 VDD.n3 GND 0.06722f
C8884 VDD.t20 GND 0.02776f
C8885 VDD.n11 GND 0.0482f
C8886 VDD.t69 GND 0.02776f
C8887 VDD.n13 GND 0.06691f
C8888 VDD.n78 GND 0.10878f
C8889 VDD.t67 GND 0.01142f
C8890 VDD.n85 GND 0.01744f
C8891 VDD.n111 GND 0.01267f
C8892 VDD.n112 GND 0.01544f
C8893 VDD.n144 GND 0.01336f
C8894 VDD.n167 GND 0.02834f
C8895 VDD.n172 GND 0.01267f
C8896 VDD.n173 GND 0.01544f
C8897 VDD.n178 GND 0.02834f
C8898 VDD.n179 GND 3.71926f
C8899 VDD.n180 GND 6.87453f
C8900 VDD.n181 GND 0.19374f
C8901 VDD.n192 GND 0.01864f
C8902 VDD.n193 GND 0.01386f
C8903 VDD.t63 GND 0.01429f
C8904 VDD.n194 GND 0.01038f
C8905 VDD.n217 GND 0.01038f
C8906 VDD.n218 GND 0.01038f
C8907 VDD.n241 GND 0.01038f
C8908 VDD.n242 GND 0.01038f
C8909 VDD.n265 GND 0.01038f
C8910 VDD.n266 GND 0.01038f
C8911 VDD.n289 GND 0.01038f
C8912 VDD.n290 GND 0.01038f
C8913 VDD.n301 GND 0.20066f
C8914 VDD.n302 GND 0.14162f
C8915 VDD.n303 GND 0.01887f
C8916 VDD.t179 GND 0.01065f
C8917 VDD.t49 GND 0.01531f
C8918 VDD.t203 GND 0.01426f
C8919 VDD.n343 GND 0.01451f
C8920 VDD.n381 GND 0.01223f
C8921 VDD.t77 GND 0.01229f
C8922 VDD.n382 GND 0.01012f
C8923 VDD.n384 GND 0.02583f
C8924 VDD.n385 GND 0.03536f
C8925 VDD.n387 GND 0.01915f
C8926 VDD.n400 GND 0.0103f
C8927 VDD.t43 GND 0.01036f
C8928 VDD.n417 GND 0.0109f
C8929 VDD.t129 GND 0.02898f
C8930 VDD.n418 GND 0.02978f
C8931 VDD.n419 GND 0.01286f
C8932 VDD.n420 GND 0.06614f
C8933 VDD.n421 GND 0.02983f
C8934 VDD.n422 GND 0.01331f
C8935 VDD.n436 GND 0.03978f
C8936 VDD.n440 GND 0.09626f
C8937 VDD.n441 GND 0.08433f
C8938 VDD.n442 GND 4.46151f
C8939 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t2 GND 0.04341f
C8940 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t3 GND 0.04341f
C8941 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n0 GND 0.09533f
C8942 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n1 GND 0.04112f
C8943 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t4 GND 0.07176f
C8944 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t11 GND 0.04479f
C8945 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n2 GND 0.14268f
C8946 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t8 GND 0.07186f
C8947 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t16 GND 0.04486f
C8948 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n3 GND 0.13678f
C8949 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n4 GND 0.02691f
C8950 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n5 GND 0.06791f
C8951 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t9 GND 0.04479f
C8952 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t6 GND 0.07176f
C8953 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n6 GND 0.14129f
C8954 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n7 GND 0.19926f
C8955 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n8 GND 0.69128f
C8956 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t10 GND 0.07196f
C8957 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t14 GND 0.04495f
C8958 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n9 GND 0.13234f
C8959 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n10 GND 0.10406f
C8960 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n11 GND 0.77672f
C8961 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t15 GND 0.04479f
C8962 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t13 GND 0.07176f
C8963 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n12 GND 0.14129f
C8964 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n13 GND 0.19036f
C8965 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n14 GND 0.75233f
C8966 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t7 GND 0.07186f
C8967 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t12 GND 0.04486f
C8968 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n15 GND 0.13678f
C8969 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n16 GND 0.30498f
C8970 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n17 GND 1.04101f
C8971 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t17 GND 0.04479f
C8972 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t5 GND 0.07176f
C8973 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n18 GND 0.14124f
C8974 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n19 GND 0.13864f
C8975 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n20 GND 4.55762f
C8976 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n21 GND 12.0001f
C8977 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n22 GND 0.56248f
C8978 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t0 GND 0.02821f
C8979 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t1 GND 0.02821f
C8980 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n23 GND 0.06728f
C8981 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n24 GND 0.13217f
.ends

