magic
tech sky130A
magscale 1 2
timestamp 1750847318
<< pwell >>
rect -278 -1109 278 1109
<< mvnmos >>
rect -50 767 50 851
rect -50 527 50 611
rect -50 287 50 371
rect -50 47 50 131
rect -50 -193 50 -109
rect -50 -433 50 -349
rect -50 -673 50 -589
rect -50 -913 50 -829
<< mvndiff >>
rect -108 839 -50 851
rect -108 779 -96 839
rect -62 779 -50 839
rect -108 767 -50 779
rect 50 839 108 851
rect 50 779 62 839
rect 96 779 108 839
rect 50 767 108 779
rect -108 599 -50 611
rect -108 539 -96 599
rect -62 539 -50 599
rect -108 527 -50 539
rect 50 599 108 611
rect 50 539 62 599
rect 96 539 108 599
rect 50 527 108 539
rect -108 359 -50 371
rect -108 299 -96 359
rect -62 299 -50 359
rect -108 287 -50 299
rect 50 359 108 371
rect 50 299 62 359
rect 96 299 108 359
rect 50 287 108 299
rect -108 119 -50 131
rect -108 59 -96 119
rect -62 59 -50 119
rect -108 47 -50 59
rect 50 119 108 131
rect 50 59 62 119
rect 96 59 108 119
rect 50 47 108 59
rect -108 -121 -50 -109
rect -108 -181 -96 -121
rect -62 -181 -50 -121
rect -108 -193 -50 -181
rect 50 -121 108 -109
rect 50 -181 62 -121
rect 96 -181 108 -121
rect 50 -193 108 -181
rect -108 -361 -50 -349
rect -108 -421 -96 -361
rect -62 -421 -50 -361
rect -108 -433 -50 -421
rect 50 -361 108 -349
rect 50 -421 62 -361
rect 96 -421 108 -361
rect 50 -433 108 -421
rect -108 -601 -50 -589
rect -108 -661 -96 -601
rect -62 -661 -50 -601
rect -108 -673 -50 -661
rect 50 -601 108 -589
rect 50 -661 62 -601
rect 96 -661 108 -601
rect 50 -673 108 -661
rect -108 -841 -50 -829
rect -108 -901 -96 -841
rect -62 -901 -50 -841
rect -108 -913 -50 -901
rect 50 -841 108 -829
rect 50 -901 62 -841
rect 96 -901 108 -841
rect 50 -913 108 -901
<< mvndiffc >>
rect -96 779 -62 839
rect 62 779 96 839
rect -96 539 -62 599
rect 62 539 96 599
rect -96 299 -62 359
rect 62 299 96 359
rect -96 59 -62 119
rect 62 59 96 119
rect -96 -181 -62 -121
rect 62 -181 96 -121
rect -96 -421 -62 -361
rect 62 -421 96 -361
rect -96 -661 -62 -601
rect 62 -661 96 -601
rect -96 -901 -62 -841
rect 62 -901 96 -841
<< mvpsubdiff >>
rect -242 1061 242 1073
rect -242 1027 -134 1061
rect 134 1027 242 1061
rect -242 1015 242 1027
rect -242 965 -184 1015
rect -242 -965 -230 965
rect -196 -965 -184 965
rect 184 965 242 1015
rect -242 -1015 -184 -965
rect 184 -965 196 965
rect 230 -965 242 965
rect 184 -1015 242 -965
rect -242 -1027 242 -1015
rect -242 -1061 -134 -1027
rect 134 -1061 242 -1027
rect -242 -1073 242 -1061
<< mvpsubdiffcont >>
rect -134 1027 134 1061
rect -230 -965 -196 965
rect 196 -965 230 965
rect -134 -1061 134 -1027
<< poly >>
rect -50 923 50 939
rect -50 889 -34 923
rect 34 889 50 923
rect -50 851 50 889
rect -50 741 50 767
rect -50 683 50 699
rect -50 649 -34 683
rect 34 649 50 683
rect -50 611 50 649
rect -50 501 50 527
rect -50 443 50 459
rect -50 409 -34 443
rect 34 409 50 443
rect -50 371 50 409
rect -50 261 50 287
rect -50 203 50 219
rect -50 169 -34 203
rect 34 169 50 203
rect -50 131 50 169
rect -50 21 50 47
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -219 50 -193
rect -50 -277 50 -261
rect -50 -311 -34 -277
rect 34 -311 50 -277
rect -50 -349 50 -311
rect -50 -459 50 -433
rect -50 -517 50 -501
rect -50 -551 -34 -517
rect 34 -551 50 -517
rect -50 -589 50 -551
rect -50 -699 50 -673
rect -50 -757 50 -741
rect -50 -791 -34 -757
rect 34 -791 50 -757
rect -50 -829 50 -791
rect -50 -939 50 -913
<< polycont >>
rect -34 889 34 923
rect -34 649 34 683
rect -34 409 34 443
rect -34 169 34 203
rect -34 -71 34 -37
rect -34 -311 34 -277
rect -34 -551 34 -517
rect -34 -791 34 -757
<< locali >>
rect -230 1027 -134 1061
rect 134 1027 230 1061
rect -230 965 -196 1027
rect 196 965 230 1027
rect -50 889 -34 923
rect 34 889 50 923
rect -96 839 -62 855
rect -96 763 -62 779
rect 62 839 96 855
rect 62 763 96 779
rect -50 649 -34 683
rect 34 649 50 683
rect -96 599 -62 615
rect -96 523 -62 539
rect 62 599 96 615
rect 62 523 96 539
rect -50 409 -34 443
rect 34 409 50 443
rect -96 359 -62 375
rect -96 283 -62 299
rect 62 359 96 375
rect 62 283 96 299
rect -50 169 -34 203
rect 34 169 50 203
rect -96 119 -62 135
rect -96 43 -62 59
rect 62 119 96 135
rect 62 43 96 59
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -197 -62 -181
rect 62 -121 96 -105
rect 62 -197 96 -181
rect -50 -311 -34 -277
rect 34 -311 50 -277
rect -96 -361 -62 -345
rect -96 -437 -62 -421
rect 62 -361 96 -345
rect 62 -437 96 -421
rect -50 -551 -34 -517
rect 34 -551 50 -517
rect -96 -601 -62 -585
rect -96 -677 -62 -661
rect 62 -601 96 -585
rect 62 -677 96 -661
rect -50 -791 -34 -757
rect 34 -791 50 -757
rect -96 -841 -62 -825
rect -96 -917 -62 -901
rect 62 -841 96 -825
rect 62 -917 96 -901
rect -230 -1027 -196 -965
rect 196 -1027 230 -965
rect -230 -1061 -134 -1027
rect 134 -1061 230 -1027
<< viali >>
rect -26 889 26 923
rect -96 779 -62 839
rect 62 779 96 839
rect -26 649 26 683
rect -96 539 -62 599
rect 62 539 96 599
rect -26 409 26 443
rect -96 299 -62 359
rect 62 299 96 359
rect -26 169 26 203
rect -96 59 -62 119
rect 62 59 96 119
rect -26 -71 26 -37
rect -96 -181 -62 -121
rect 62 -181 96 -121
rect -26 -311 26 -277
rect -96 -421 -62 -361
rect 62 -421 96 -361
rect -26 -551 26 -517
rect -96 -661 -62 -601
rect 62 -661 96 -601
rect -26 -791 26 -757
rect -96 -901 -62 -841
rect 62 -901 96 -841
<< metal1 >>
rect -38 923 38 929
rect -38 889 -26 923
rect 26 889 38 923
rect -38 883 38 889
rect -102 839 -56 851
rect -102 779 -96 839
rect -62 779 -56 839
rect -102 767 -56 779
rect 56 839 102 851
rect 56 779 62 839
rect 96 779 102 839
rect 56 767 102 779
rect -38 683 38 689
rect -38 649 -26 683
rect 26 649 38 683
rect -38 643 38 649
rect -102 599 -56 611
rect -102 539 -96 599
rect -62 539 -56 599
rect -102 527 -56 539
rect 56 599 102 611
rect 56 539 62 599
rect 96 539 102 599
rect 56 527 102 539
rect -38 443 38 449
rect -38 409 -26 443
rect 26 409 38 443
rect -38 403 38 409
rect -102 359 -56 371
rect -102 299 -96 359
rect -62 299 -56 359
rect -102 287 -56 299
rect 56 359 102 371
rect 56 299 62 359
rect 96 299 102 359
rect 56 287 102 299
rect -38 203 38 209
rect -38 169 -26 203
rect 26 169 38 203
rect -38 163 38 169
rect -102 119 -56 131
rect -102 59 -96 119
rect -62 59 -56 119
rect -102 47 -56 59
rect 56 119 102 131
rect 56 59 62 119
rect 96 59 102 119
rect 56 47 102 59
rect -38 -37 38 -31
rect -38 -71 -26 -37
rect 26 -71 38 -37
rect -38 -77 38 -71
rect -102 -121 -56 -109
rect -102 -181 -96 -121
rect -62 -181 -56 -121
rect -102 -193 -56 -181
rect 56 -121 102 -109
rect 56 -181 62 -121
rect 96 -181 102 -121
rect 56 -193 102 -181
rect -38 -277 38 -271
rect -38 -311 -26 -277
rect 26 -311 38 -277
rect -38 -317 38 -311
rect -102 -361 -56 -349
rect -102 -421 -96 -361
rect -62 -421 -56 -361
rect -102 -433 -56 -421
rect 56 -361 102 -349
rect 56 -421 62 -361
rect 96 -421 102 -361
rect 56 -433 102 -421
rect -38 -517 38 -511
rect -38 -551 -26 -517
rect 26 -551 38 -517
rect -38 -557 38 -551
rect -102 -601 -56 -589
rect -102 -661 -96 -601
rect -62 -661 -56 -601
rect -102 -673 -56 -661
rect 56 -601 102 -589
rect 56 -661 62 -601
rect 96 -661 102 -601
rect 56 -673 102 -661
rect -38 -757 38 -751
rect -38 -791 -26 -757
rect 26 -791 38 -757
rect -38 -797 38 -791
rect -102 -841 -56 -829
rect -102 -901 -96 -841
rect -62 -901 -56 -841
rect -102 -913 -56 -901
rect 56 -841 102 -829
rect 56 -901 62 -841
rect 96 -901 102 -841
rect 56 -913 102 -901
<< properties >>
string FIXED_BBOX -213 -1044 213 1044
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.420 l 0.50 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
