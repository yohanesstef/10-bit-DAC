magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1104 307 1104
<< psubdiff >>
rect -271 1034 -175 1068
rect 175 1034 271 1068
rect -271 972 -237 1034
rect 237 972 271 1034
rect -271 -1034 -237 -972
rect 237 -1034 271 -972
rect -271 -1068 -175 -1034
rect 175 -1068 271 -1034
<< psubdiffcont >>
rect -175 1034 175 1068
rect -271 -972 -237 972
rect 237 -972 271 972
rect -175 -1068 175 -1034
<< xpolycontact >>
rect -141 506 141 938
rect -141 -938 141 -506
<< xpolyres >>
rect -141 -506 141 506
<< locali >>
rect -271 1034 -175 1068
rect 175 1034 271 1068
rect -271 972 -237 1034
rect 237 972 271 1034
rect -271 -1034 -237 -972
rect 237 -1034 271 -972
rect -271 -1068 -175 -1034
rect 175 -1068 271 -1034
<< viali >>
rect -125 523 125 920
rect -125 -920 125 -523
<< metal1 >>
rect -131 920 131 932
rect -131 523 -125 920
rect 125 523 131 920
rect -131 511 131 523
rect -131 -523 131 -511
rect -131 -920 -125 -523
rect 125 -920 131 -523
rect -131 -932 131 -920
<< properties >>
string FIXED_BBOX -254 -1051 254 1051
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 5.218 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 7.668k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
