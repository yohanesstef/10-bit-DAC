* NGSPICE file created from rseg_3_v3.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_SEMVNL a_n141_n733# a_n141_301# VSUBS
X0 a_n141_301# a_n141_n733# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.17
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_SEMXNL a_n141_n733# a_n141_301# VSUBS
X0 a_n141_301# a_n141_n733# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.17
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_GLTCMD a_n141_311# a_n141_n743# VSUBS
X0 a_n141_311# a_n141_n743# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.27
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_42QADH a_n141_n748# a_n141_316# VSUBS
X0 a_n141_316# a_n141_n748# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.32
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_AFTT8S a_n141_n769# a_n141_337# VSUBS
X0 a_n141_337# a_n141_n769# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.53
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_GVNVJY a_n141_n753# a_n141_321# VSUBS
X0 a_n141_321# a_n141_n753# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.37
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_DZKNT5 a_n141_367# a_n141_n799# VSUBS
X0 a_n141_367# a_n141_n799# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.83
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_J5YLPL a_n141_n774# a_n141_342# VSUBS
X0 a_n141_342# a_n141_n774# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.58
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_47PAZ6 a_n141_n784# a_n141_352# VSUBS
X0 a_n141_352# a_n141_n784# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.68
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_DZKLT5 a_n141_367# a_n141_n799# VSUBS
X0 a_n141_367# a_n141_n799# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.83
.ends

.subckt rseg_3_1 sky130_fd_pr__res_xhigh_po_1p41_DZKNT5_0/a_n141_367# XR1/a_n141_n733#
+ sky130_fd_pr__res_xhigh_po_1p41_SEMVNL_0/a_n141_301# sky130_fd_pr__res_xhigh_po_1p41_DZKNT5_0/a_n141_n799#
+ m1_6357_n4745# m1_4812_n3449# sky130_fd_pr__res_xhigh_po_1p41_SEMVNL_0/a_n141_n733#
+ m1_6332_n4421# m1_4786_n4097# m1_6301_n2801# m1_4827_n2539# m1_6311_n3773# VSUBS
+ m1_4745_n4745#
Xsky130_fd_pr__res_xhigh_po_1p41_SEMVNL_0 sky130_fd_pr__res_xhigh_po_1p41_SEMVNL_0/a_n141_n733#
+ sky130_fd_pr__res_xhigh_po_1p41_SEMVNL_0/a_n141_301# VSUBS sky130_fd_pr__res_xhigh_po_1p41_SEMVNL
XXR1 XR1/a_n141_n733# m1_4827_n2539# VSUBS sky130_fd_pr__res_xhigh_po_1p41_SEMXNL
XXR2 m1_4827_n2539# m1_6301_n2801# VSUBS sky130_fd_pr__res_xhigh_po_1p41_GLTCMD
XXR3 m1_6301_n2801# m1_4812_n3449# VSUBS sky130_fd_pr__res_xhigh_po_1p41_42QADH
XXR5 m1_6311_n3773# m1_4786_n4097# VSUBS sky130_fd_pr__res_xhigh_po_1p41_AFTT8S
XXR4 m1_6311_n3773# m1_4812_n3449# VSUBS sky130_fd_pr__res_xhigh_po_1p41_GVNVJY
Xsky130_fd_pr__res_xhigh_po_1p41_DZKNT5_0 sky130_fd_pr__res_xhigh_po_1p41_DZKNT5_0/a_n141_367#
+ sky130_fd_pr__res_xhigh_po_1p41_DZKNT5_0/a_n141_n799# VSUBS sky130_fd_pr__res_xhigh_po_1p41_DZKNT5
XXR6 m1_6332_n4421# m1_4786_n4097# VSUBS sky130_fd_pr__res_xhigh_po_1p41_J5YLPL
XXR7 m1_6332_n4421# m1_4745_n4745# VSUBS sky130_fd_pr__res_xhigh_po_1p41_47PAZ6
XXR8 m1_4745_n4745# m1_6357_n4745# VSUBS sky130_fd_pr__res_xhigh_po_1p41_DZKLT5
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_QX57C3 a_n141_n825# a_n141_393# VSUBS
X0 a_n141_393# a_n141_n825# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=4.09
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_H2U5BC a_n141_n835# a_n141_403# VSUBS
X0 a_n141_403# a_n141_n835# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=4.19
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_E2U9YT a_n141_n861# a_n141_429# VSUBS
X0 a_n141_429# a_n141_n861# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=4.45
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_YY58WS a_n141_378# a_n141_n810# VSUBS
X0 a_n141_378# a_n141_n810# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.94
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_KLD4QF a_n141_n902# a_n141_470# VSUBS
X0 a_n141_470# a_n141_n902# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=4.86
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_4F76E7 a_n141_n876# a_n141_444# VSUBS
X0 a_n141_444# a_n141_n876# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=4.6
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_HDPFLR a_n141_n928# a_n141_496# VSUBS
X0 a_n141_496# a_n141_n928# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=5.12
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_5X53DF a_n141_526# a_n141_n958# VSUBS
X0 a_n141_526# a_n141_n958# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=5.42
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_YY56WS a_n141_378# a_n141_n810# VSUBS
X0 a_n141_378# a_n141_n810# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.94
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF a_n141_526# a_n141_n958# VSUBS
X0 a_n141_526# a_n141_n958# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=5.42
.ends

.subckt rseg_3_2 XR9/a_n141_n810# m1_8330_n3320# sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF_0/a_n141_526#
+ XR16/a_n141_n958# sky130_fd_pr__res_xhigh_po_1p41_YY58WS_0/a_n141_n810# m1_8304_n3968#
+ sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF_0/a_n141_n958# m1_10152_n3644# m1_10116_n4292#
+ m1_8375_n2410# m1_10193_n2996# m1_8263_n4616# sky130_fd_pr__res_xhigh_po_1p41_YY58WS_0/a_n141_378#
+ VSUBS
XXR10 m1_10116_n4292# m1_8263_n4616# VSUBS sky130_fd_pr__res_xhigh_po_1p41_QX57C3
XXR11 m1_10116_n4292# m1_8304_n3968# VSUBS sky130_fd_pr__res_xhigh_po_1p41_H2U5BC
XXR12 m1_10152_n3644# m1_8304_n3968# VSUBS sky130_fd_pr__res_xhigh_po_1p41_E2U9YT
Xsky130_fd_pr__res_xhigh_po_1p41_YY58WS_0 sky130_fd_pr__res_xhigh_po_1p41_YY58WS_0/a_n141_378#
+ sky130_fd_pr__res_xhigh_po_1p41_YY58WS_0/a_n141_n810# VSUBS sky130_fd_pr__res_xhigh_po_1p41_YY58WS
XXR14 m1_10193_n2996# m1_8330_n3320# VSUBS sky130_fd_pr__res_xhigh_po_1p41_KLD4QF
XXR13 m1_10152_n3644# m1_8330_n3320# VSUBS sky130_fd_pr__res_xhigh_po_1p41_4F76E7
XXR15 m1_10193_n2996# m1_8375_n2410# VSUBS sky130_fd_pr__res_xhigh_po_1p41_HDPFLR
XXR16 m1_8375_n2410# XR16/a_n141_n958# VSUBS sky130_fd_pr__res_xhigh_po_1p41_5X53DF
XXR9 m1_8263_n4616# XR9/a_n141_n810# VSUBS sky130_fd_pr__res_xhigh_po_1p41_YY56WS
Xsky130_fd_pr__res_xhigh_po_1p41_5X5ZCF_0 sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF_0/a_n141_526#
+ sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF_0/a_n141_n958# VSUBS sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF
.ends

.subckt rseg_3_v3 v0 v1 v2 v3 v4 v5 v6 v7 v8 v9 v10 v11 v12 v13 v14 v15 v16 gnd
Xrseg_3_1_0 gnd v0 gnd gnd v8 v3 gnd v6 v5 v2 v1 v4 gnd v7 rseg_3_1
Xrseg_3_2_0 v8 v13 gnd v16 gnd v11 gnd v12 v10 v15 v14 v9 gnd gnd rseg_3_2
.ends

