magic
tech sky130A
magscale 1 2
timestamp 1749057406
<< pwell >>
rect -307 -965 307 965
<< psubdiff >>
rect -271 895 -175 929
rect 175 895 271 929
rect -271 833 -237 895
rect 237 833 271 895
rect -271 -895 -237 -833
rect 237 -895 271 -833
rect -271 -929 -175 -895
rect 175 -929 271 -895
<< psubdiffcont >>
rect -175 895 175 929
rect -271 -833 -237 833
rect 237 -833 271 833
rect -175 -929 175 -895
<< xpolycontact >>
rect -141 367 141 799
rect -141 -799 141 -367
<< xpolyres >>
rect -141 -367 141 367
<< locali >>
rect -271 895 -175 929
rect 175 895 271 929
rect -271 833 -237 895
rect 237 833 271 895
rect -271 -895 -237 -833
rect 237 -895 271 -833
rect -271 -929 -175 -895
rect 175 -929 271 -895
<< viali >>
rect -125 384 125 781
rect -125 -781 125 -384
<< metal1 >>
rect -131 781 131 793
rect -131 384 -125 781
rect 125 384 131 781
rect -131 372 131 384
rect -131 -384 131 -372
rect -131 -781 -125 -384
rect 125 -781 131 -384
rect -131 -793 131 -781
<< properties >>
string FIXED_BBOX -254 -912 254 912
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 3.834 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 5.705k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
