* PEX produced on Fri Jun 13 01:01:18 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from logic_shift_seg2.ext - technology: sky130A

.subckt logic_shift_seg2_posim b[6] b[7] b[8] b[9] bb[6] bb[7] bb[8] BS[8] BS[9] BSB[8]
+ BSB[9] VDD GND
X0 VDD.t32 b[6].t0 x5.C.t1 VDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 x5.C.t2 b[6].t1 a_5195_n3687.t1 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 x3.Y.t2 b[9].t0 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 BSB[9].t1 BS[9].t4 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4 x2.Y.t2 b[9].t1 VDD.t27 VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_6203_n3687.t1 bb[8].t0 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VDD.t37 x6.Y.t3 BS[8].t2 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7 x5.A.t3 bb[8].t1 VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 a_5643_n3687.t1 x6.Y.t4 a_5559_n3687.t1 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VDD.t7 b[7].t0 x3.Y.t0 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 BS[8].t0 x5.C.t3 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_5559_n3687.t0 x5.C.t4 GND.t12 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VDD.t31 b[6].t2 x2.Y.t1 VDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_6287_n3687.t1 bb[7].t0 a_6203_n3687.t0 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 x1.Y.t1 b[9].t2 a_4919_n2823.t1 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VDD.t5 bb[7].t1 x5.A.t2 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X16 a_5919_n2823.t0 x2.Y.t3 a_5835_n2823.t1 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_4919_n2823.t0 b[8].t0 GND.t18 GND.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X18 x5.A.t0 bb[6].t0 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X19 x6.Y.t0 b[8].t1 a_4919_n3687.t0 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 x5.A.t1 bb[6].t1 a_6287_n3687.t0 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X21 BS[9].t3 x1.Y.t3 a_5919_n2823.t1 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X22 VDD.t9 b[8].t2 x6.Y.t1 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 x6.Y.t2 b[7].t1 VDD.t35 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X24 a_4919_n3687.t1 b[7].t2 GND.t16 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X25 BS[8].t3 x5.A.t4 a_5643_n3687.t0 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X26 a_5835_n2823.t0 x3.Y.t3 GND.t6 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 BS[8].t1 x5.A.t5 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X28 a_5563_n2823.t1 b[9].t3 GND.t14 GND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X29 BSB[9].t0 BS[9].t5 GND.t22 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X30 a_5195_n2823.t1 b[9].t4 GND.t29 GND.t28 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VDD.t14 b[9].t5 x1.Y.t2 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X32 VDD.t13 x2.Y.t4 BS[9].t0 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X33 x1.Y.t0 b[8].t3 VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 a_5195_n3687.t0 b[8].t4 GND.t8 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X35 x5.C.t0 b[8].t5 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X36 x3.Y.t1 b[7].t3 a_5563_n2823.t0 GND.t26 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 BS[9].t1 x1.Y.t4 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X38 BS[9].t2 x3.Y.t4 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X39 x2.Y.t0 b[6].t3 a_5195_n2823.t0 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X40 BSB[8].t1 BS[8].t4 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X41 BSB[8].t0 BS[8].t5 GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 b[6].n0 b[6].t2 230.155
R1 b[6].n3 b[6].t0 230.155
R2 b[6].n0 b[6].t3 157.856
R3 b[6].n3 b[6].t1 157.856
R4 b[6].n1 b[6].n0 154.867
R5 b[6].n4 b[6].n3 152
R6 b[6].n4 b[6].n2 21.3533
R7 b[6].n2 b[6].n1 18.3823
R8 b[6] b[6].n4 2.10199
R9 b[6].n1 b[6] 1.52886
R10 b[6].n2 b[6] 0.484875
R11 x5.C x5.C.n0 237.577
R12 x5.C.n2 x5.C.t3 230.363
R13 x5.C.n2 x5.C.t4 158.064
R14 x5.C.n3 x5.C.n2 152.553
R15 x5.C.n1 x5.C.t2 140.53
R16 x5.C.n0 x5.C.t1 26.5955
R17 x5.C.n0 x5.C.t0 26.5955
R18 x5.C.n4 x5.C.n3 20.0033
R19 x5.C x5.C.n4 11.2946
R20 x5.C.n1 x5.C 9.03579
R21 x5.C.n4 x5.C.n1 5.27109
R22 x5.C.n1 x5.C 1.72748
R23 x5.C.n3 x5.C 1.54533
R24 VDD.n16 VDD.n13 318.305
R25 VDD.n22 VDD.n8 318.303
R26 VDD.n29 VDD.n4 313.575
R27 VDD.n6 VDD.t34 255.905
R28 VDD.n12 VDD.t29 255.904
R29 VDD.n26 VDD.t3 249.901
R30 VDD.n2 VDD.t11 249.52
R31 VDD.n20 VDD.t16 249.387
R32 VDD.n40 VDD.t9 249.363
R33 VDD.n1 VDD.t32 249.363
R34 VDD.n40 VDD.t14 249.362
R35 VDD.n1 VDD.t31 249.362
R36 VDD.n36 VDD.t35 247.394
R37 VDD.n41 VDD.t22 247.394
R38 VDD.n36 VDD.t24 247.394
R39 VDD.n41 VDD.t27 247.394
R40 VDD.n2 VDD.t26 247.394
R41 VDD.n27 VDD.t7 245.178
R42 VDD.t30 VDD.n47 234.982
R43 VDD.t0 VDD 216.519
R44 VDD.n20 VDD.n10 213.119
R45 VDD VDD.t19 208.127
R46 VDD.t8 VDD 204.77
R47 VDD.n48 VDD 197.325
R48 VDD.t17 VDD.t6 154.417
R49 VDD.t21 VDD.t30 140.989
R50 VDD.t23 VDD.t8 140.989
R51 VDD.t36 VDD.t25 134.276
R52 VDD.n47 VDD 124.206
R53 VDD VDD.t21 117.492
R54 VDD VDD.t23 117.492
R55 VDD.t2 VDD 107.421
R56 VDD.t10 VDD 107.421
R57 VDD.n47 VDD.n46 106.559
R58 VDD VDD.t4 95.6719
R59 VDD.t12 VDD 95.6719
R60 VDD.t4 VDD.t28 82.2443
R61 VDD.t33 VDD.t12 82.2443
R62 VDD.n10 VDD.t15 80.5659
R63 VDD.t28 VDD.t0 78.8874
R64 VDD.t19 VDD.t33 78.8874
R65 VDD VDD.t17 53.7107
R66 VDD.t15 VDD 45.3185
R67 VDD VDD.t2 45.3185
R68 VDD.n15 VDD.n14 42.2367
R69 VDD.n4 VDD.t18 38.4155
R70 VDD.n8 VDD.t20 38.4155
R71 VDD.n13 VDD.t1 38.4155
R72 VDD.n30 VDD.n29 33.1299
R73 VDD.n22 VDD.n21 27.4829
R74 VDD.n16 VDD.n15 27.4829
R75 VDD.n10 VDD 26.8556
R76 VDD.n4 VDD.t37 26.5955
R77 VDD.n8 VDD.t13 26.5955
R78 VDD.n13 VDD.t5 26.5955
R79 VDD.n40 VDD.n34 25.977
R80 VDD.n42 VDD.n1 25.977
R81 VDD.n26 VDD.n25 25.977
R82 VDD.n36 VDD.n34 24.4711
R83 VDD.n42 VDD.n41 24.4711
R84 VDD.n30 VDD.n2 24.4711
R85 VDD.n21 VDD.n20 23.7181
R86 VDD.n20 VDD.n9 23.7181
R87 VDD.n27 VDD.n26 22.9652
R88 VDD.n49 VDD.n48 18.084
R89 VDD.n36 VDD.n0 12.8005
R90 VDD.n41 VDD.n40 12.8005
R91 VDD.n46 VDD.n1 12.8005
R92 VDD.n46 VDD.n2 12.8005
R93 VDD.n15 VDD.n11 9.3005
R94 VDD.n17 VDD.n16 9.3005
R95 VDD.n18 VDD.n9 9.3005
R96 VDD.n20 VDD.n19 9.3005
R97 VDD.n21 VDD.n7 9.3005
R98 VDD.n23 VDD.n22 9.3005
R99 VDD.n25 VDD.n24 9.3005
R100 VDD.n26 VDD.n5 9.3005
R101 VDD.n28 VDD.n3 9.3005
R102 VDD.n31 VDD.n30 9.3005
R103 VDD.n32 VDD.n2 9.3005
R104 VDD.n46 VDD.n45 9.3005
R105 VDD.n44 VDD.n1 9.3005
R106 VDD.n43 VDD.n42 9.3005
R107 VDD.n41 VDD.n33 9.3005
R108 VDD.n40 VDD.n39 9.3005
R109 VDD.n38 VDD.n34 9.3005
R110 VDD.n37 VDD.n36 9.3005
R111 VDD.n35 VDD.n0 9.3005
R112 VDD.n25 VDD.n6 8.28285
R113 VDD.n12 VDD.n9 8.28285
R114 VDD.t6 VDD.t36 6.71428
R115 VDD.t25 VDD.t10 6.71428
R116 VDD.n48 VDD.n0 3.58719
R117 VDD.n29 VDD.n28 1.50638
R118 VDD.n28 VDD.n27 1.12991
R119 VDD.n22 VDD.n6 0.376971
R120 VDD.n16 VDD.n12 0.376971
R121 VDD.n14 VDD 0.324797
R122 VDD.n17 VDD.n11 0.120292
R123 VDD.n18 VDD.n17 0.120292
R124 VDD.n23 VDD.n7 0.120292
R125 VDD.n24 VDD.n23 0.120292
R126 VDD.n31 VDD.n3 0.120292
R127 VDD.n32 VDD.n31 0.120292
R128 VDD.n44 VDD.n43 0.120292
R129 VDD.n43 VDD.n33 0.120292
R130 VDD.n39 VDD.n38 0.120292
R131 VDD.n38 VDD.n37 0.120292
R132 VDD VDD.n11 0.104667
R133 VDD.n19 VDD 0.0603958
R134 VDD VDD.n7 0.0603958
R135 VDD VDD.n5 0.0603958
R136 VDD VDD.n3 0.0603958
R137 VDD.n45 VDD 0.0603958
R138 VDD VDD.n44 0.0603958
R139 VDD.n39 VDD 0.0603958
R140 VDD VDD.n35 0.0603958
R141 VDD.n49 VDD 0.0603958
R142 VDD.n14 VDD 0.0427777
R143 VDD.n45 VDD 0.03175
R144 VDD.n35 VDD 0.03175
R145 VDD VDD.n49 0.03175
R146 VDD VDD.n33 0.0239375
R147 VDD.n37 VDD 0.0239375
R148 VDD VDD.n18 0.0226354
R149 VDD.n24 VDD 0.0226354
R150 VDD.n19 VDD 0.0213333
R151 VDD.n5 VDD 0.0213333
R152 VDD VDD.n32 0.0213333
R153 a_5195_n3687.t0 a_5195_n3687.t1 49.8467
R154 GND.n77 GND.n76 8012.67
R155 GND GND.t4 5766.99
R156 GND.t21 GND 2506.15
R157 GND GND.t9 2434.95
R158 GND.n46 GND.t27 1993.53
R159 GND.n45 GND.t23 1993.53
R160 GND.n44 GND.t24 1993.53
R161 GND GND.t26 1765.7
R162 GND GND.t25 1751.46
R163 GND GND.t30 1737.22
R164 GND GND.t3 1737.22
R165 GND GND.t21 1509.39
R166 GND.t9 GND 1509.39
R167 GND.t27 GND.t19 1366.99
R168 GND.t4 GND.t2 1366.99
R169 GND.t25 GND.t20 1366.99
R170 GND.n76 GND.n2 1310.03
R171 GND.n77 GND.n1 1310.03
R172 GND.n1 GND.n0 1198.25
R173 GND.n44 GND.n43 1198.25
R174 GND.n76 GND.n75 1198.25
R175 GND.n74 GND.n2 1198.25
R176 GND.n45 GND.n8 1198.25
R177 GND.n47 GND.n46 1198.25
R178 GND.n78 GND.n77 1198.25
R179 GND.t19 GND.t5 1196.12
R180 GND.t26 GND.t13 1196.12
R181 GND.t23 GND.t28 1196.12
R182 GND.t30 GND.t17 1196.12
R183 GND.t2 GND.t0 1196.12
R184 GND.t20 GND.t11 1196.12
R185 GND.t24 GND.t7 1196.12
R186 GND.t3 GND.t15 1196.12
R187 GND GND.n44 1082.2
R188 GND.n46 GND 1067.96
R189 GND GND.n45 1053.72
R190 GND GND.n2 1053.72
R191 GND GND.n1 1053.72
R192 GND.t13 GND 996.764
R193 GND.t28 GND 996.764
R194 GND.t17 GND 996.764
R195 GND.t7 GND 996.764
R196 GND.t15 GND 996.764
R197 GND.t5 GND 911.327
R198 GND.t0 GND 911.327
R199 GND.t11 GND 911.327
R200 GND.n13 GND.t12 274.812
R201 GND.n18 GND.t1 274.812
R202 GND.n10 GND.t6 274.812
R203 GND.n20 GND.t10 158.361
R204 GND.n49 GND.t22 158.361
R205 GND.n33 GND.t16 150.922
R206 GND.n38 GND.t8 150.922
R207 GND.n73 GND.t18 150.922
R208 GND.n68 GND.t29 150.922
R209 GND.n62 GND.t14 150.922
R210 GND.n37 GND.n31 34.6358
R211 GND.n39 GND.n12 34.6358
R212 GND.n25 GND.n15 34.6358
R213 GND.n26 GND.n25 34.6358
R214 GND.n27 GND.n26 34.6358
R215 GND.n21 GND.n19 34.6358
R216 GND.n72 GND.n6 34.6358
R217 GND.n67 GND.n66 34.6358
R218 GND.n61 GND.n60 34.6358
R219 GND.n55 GND.n54 34.6358
R220 GND.n56 GND.n55 34.6358
R221 GND.n27 GND.n13 25.977
R222 GND.n56 GND.n10 25.977
R223 GND.n19 GND.n18 24.0946
R224 GND.n60 GND.n10 24.0946
R225 GND.n38 GND.n37 23.7181
R226 GND.n43 GND.n12 23.7181
R227 GND.n68 GND.n6 23.7181
R228 GND.n66 GND.n8 23.7181
R229 GND.n54 GND.n47 23.7181
R230 GND.n50 GND.n47 23.7181
R231 GND.n33 GND.n31 22.2123
R232 GND.n39 GND.n38 22.2123
R233 GND.n73 GND.n72 22.2123
R234 GND.n68 GND.n67 22.2123
R235 GND.n62 GND.n61 22.2123
R236 GND.n49 GND.n48 18.1437
R237 GND.n43 GND.n13 13.177
R238 GND.n33 GND.n0 12.8005
R239 GND.n78 GND.n0 12.8005
R240 GND.n75 GND.n74 12.8005
R241 GND.n74 GND.n73 12.8005
R242 GND.n62 GND.n8 12.8005
R243 GND.n21 GND.n20 10.5417
R244 GND.n51 GND.n50 9.3005
R245 GND.n54 GND.n53 9.3005
R246 GND.n55 GND.n11 9.3005
R247 GND.n57 GND.n56 9.3005
R248 GND.n58 GND.n10 9.3005
R249 GND.n60 GND.n59 9.3005
R250 GND.n61 GND.n9 9.3005
R251 GND.n63 GND.n62 9.3005
R252 GND.n64 GND.n8 9.3005
R253 GND.n66 GND.n65 9.3005
R254 GND.n67 GND.n7 9.3005
R255 GND.n69 GND.n68 9.3005
R256 GND.n70 GND.n6 9.3005
R257 GND.n72 GND.n71 9.3005
R258 GND.n73 GND.n5 9.3005
R259 GND.n74 GND.n4 9.3005
R260 GND.n75 GND.n3 9.3005
R261 GND.n52 GND.n47 9.3005
R262 GND.n79 GND.n78 9.3005
R263 GND.n19 GND.n16 9.3005
R264 GND.n22 GND.n21 9.3005
R265 GND.n23 GND.n15 9.3005
R266 GND.n25 GND.n24 9.3005
R267 GND.n26 GND.n14 9.3005
R268 GND.n28 GND.n27 9.3005
R269 GND.n29 GND.n13 9.3005
R270 GND.n43 GND.n42 9.3005
R271 GND.n41 GND.n12 9.3005
R272 GND.n40 GND.n39 9.3005
R273 GND.n38 GND.n30 9.3005
R274 GND.n37 GND.n36 9.3005
R275 GND.n35 GND.n31 9.3005
R276 GND.n34 GND.n33 9.3005
R277 GND.n32 GND.n0 9.3005
R278 GND.n18 GND.n17 7.25901
R279 GND.n20 GND.n15 6.77697
R280 GND.n50 GND.n49 6.77697
R281 GND.n17 GND 0.796776
R282 GND.n48 GND 0.200356
R283 GND.n51 GND.n48 0.14581
R284 GND.n53 GND.n11 0.120292
R285 GND.n57 GND.n11 0.120292
R286 GND.n58 GND.n57 0.120292
R287 GND.n59 GND.n9 0.120292
R288 GND.n63 GND.n9 0.120292
R289 GND.n65 GND.n7 0.120292
R290 GND.n69 GND.n7 0.120292
R291 GND.n71 GND.n70 0.120292
R292 GND.n71 GND.n5 0.120292
R293 GND.n22 GND.n16 0.120292
R294 GND.n23 GND.n22 0.120292
R295 GND.n24 GND.n14 0.120292
R296 GND.n28 GND.n14 0.120292
R297 GND.n29 GND.n28 0.120292
R298 GND.n41 GND.n40 0.120292
R299 GND.n40 GND.n30 0.120292
R300 GND.n36 GND.n35 0.120292
R301 GND.n35 GND.n34 0.120292
R302 GND.n52 GND 0.0603958
R303 GND.n53 GND 0.0603958
R304 GND.n59 GND 0.0603958
R305 GND.n64 GND 0.0603958
R306 GND.n65 GND 0.0603958
R307 GND.n70 GND 0.0603958
R308 GND GND.n4 0.0603958
R309 GND GND.n3 0.0603958
R310 GND GND.n16 0.0603958
R311 GND.n24 GND 0.0603958
R312 GND.n42 GND 0.0603958
R313 GND GND.n41 0.0603958
R314 GND.n36 GND 0.0603958
R315 GND GND.n32 0.0603958
R316 GND.n79 GND 0.0603958
R317 GND.n17 GND 0.0535408
R318 GND GND.n52 0.0330521
R319 GND GND.n64 0.0330521
R320 GND.n4 GND 0.0330521
R321 GND.n3 GND 0.0330521
R322 GND.n42 GND 0.0330521
R323 GND.n32 GND 0.0330521
R324 GND GND.n79 0.0330521
R325 GND GND.n63 0.0239375
R326 GND GND.n69 0.0239375
R327 GND.n5 GND 0.0239375
R328 GND GND.n30 0.0239375
R329 GND.n34 GND 0.0239375
R330 GND GND.n51 0.0226354
R331 GND GND.n23 0.0226354
R332 GND GND.n58 0.0213333
R333 GND GND.n29 0.0213333
R334 b[9].n1 b[9].t5 230.155
R335 b[9].n0 b[9].t1 229.369
R336 b[9].n5 b[9].t0 229.369
R337 b[9] b[9].n0 157.927
R338 b[9].n1 b[9].t2 157.856
R339 b[9].n0 b[9].t4 157.07
R340 b[9].n5 b[9].t3 157.07
R341 b[9].n2 b[9].n1 152
R342 b[9].n6 b[9].n5 152
R343 b[9].n3 b[9].n2 13.1513
R344 b[9].n6 b[9].n4 11.8414
R345 b[9].n4 b[9].n3 9.3005
R346 b[9].n3 b[9] 7.11161
R347 b[9].n4 b[9] 6.86887
R348 b[9] b[9].n6 4.39453
R349 b[9].n2 b[9] 2.3045
R350 x3.Y.n3 x3.Y.t4 230.363
R351 x3.Y.n5 x3.Y.n2 203.147
R352 x3.Y.n3 x3.Y.t3 158.064
R353 x3.Y.n4 x3.Y.n3 156.364
R354 x3.Y.n0 x3.Y.t1 132.067
R355 x3.Y.n2 x3.Y.t0 26.5955
R356 x3.Y.n2 x3.Y.t2 26.5955
R357 x3.Y x3.Y.n5 21.6304
R358 x3.Y.n5 x3.Y.n4 19.7021
R359 x3.Y.n1 x3.Y.n0 4.15748
R360 x3.Y x3.Y.n1 3.76521
R361 x3.Y.n4 x3.Y 2.32777
R362 x3.Y.n0 x3.Y 1.17559
R363 x3.Y.n1 x3.Y 0.921363
R364 BS[9].n2 BS[9].t1 274.793
R365 BS[9].n0 BS[9].t4 230.576
R366 BS[9].n2 BS[9].n1 205.28
R367 BS[9].n0 BS[9].t5 158.275
R368 BS[9].n4 BS[9].n0 153.067
R369 BS[9].n3 BS[9].t3 133.124
R370 BS[9] BS[9].n2 67.4857
R371 BS[9].n3 BS[9] 36.3299
R372 BS[9].n1 BS[9].t0 26.5955
R373 BS[9].n1 BS[9].t2 26.5955
R374 BS[9].n4 BS[9] 10.0554
R375 BS[9] BS[9].n3 9.93288
R376 BS[9] BS[9].n4 5.6005
R377 BSB[9] BSB[9].t1 230.518
R378 BSB[9] BSB[9].t0 159.29
R379 BSB[9].n0 BSB[9] 14.7483
R380 BSB[9] BSB[9].n0 7.23528
R381 BSB[9].n0 BSB[9] 5.04292
R382 x2.Y.t0 x2.Y 272.038
R383 x2.Y.n4 x2.Y.t0 258.846
R384 x2.Y.n1 x2.Y.t4 241.536
R385 x2.Y.n3 x2.Y.n0 195.704
R386 x2.Y.n1 x2.Y.t3 169.237
R387 x2.Y.n2 x2.Y.n1 154.514
R388 x2.Y x2.Y.n3 29.0733
R389 x2.Y.n0 x2.Y.t1 26.5955
R390 x2.Y.n0 x2.Y.t2 26.5955
R391 x2.Y.n3 x2.Y.n2 25.6543
R392 x2.Y.n5 x2.Y 3.76521
R393 x2.Y.n5 x2.Y.n4 3.03935
R394 x2.Y.n4 x2.Y 2.30266
R395 x2.Y x2.Y.n5 0.921363
R396 x2.Y.n2 x2.Y 0.229071
R397 bb[8].n0 bb[8].t1 230.363
R398 bb[8].n0 bb[8].t0 158.064
R399 bb[8].n1 bb[8].n0 152
R400 bb[8].n1 bb[8] 22.4019
R401 bb[8] bb[8].n1 3.2005
R402 a_6203_n3687.t0 a_6203_n3687.t1 49.8467
R403 x6.Y.n2 x6.Y.t0 268.077
R404 x6.Y.n2 x6.Y.t0 258.846
R405 x6.Y.n1 x6.Y.t3 241.536
R406 x6.Y x6.Y.n0 237.577
R407 x6.Y.n1 x6.Y.t4 169.237
R408 x6.Y x6.Y.n1 153.877
R409 x6.Y.n2 x6.Y 29.7595
R410 x6.Y.n0 x6.Y.t1 26.5955
R411 x6.Y.n0 x6.Y.t2 26.5955
R412 x6.Y.n3 x6.Y 16.5652
R413 x6.Y.n3 x6.Y 9.03579
R414 x6.Y.n3 x6.Y.n2 8.8386
R415 x6.Y x6.Y.n3 1.72748
R416 BS[8].n3 BS[8].t1 230.712
R417 BS[8].n0 BS[8].t4 230.576
R418 BS[8].n2 BS[8].n1 205.28
R419 BS[8] BS[8].t3 169.452
R420 BS[8].n0 BS[8].t5 158.275
R421 BS[8].n4 BS[8].n0 153.067
R422 BS[8].n2 BS[8] 67.4857
R423 BS[8].n3 BS[8].n2 44.0818
R424 BS[8].n1 BS[8].t2 26.5955
R425 BS[8].n1 BS[8].t0 26.5955
R426 BS[8].n4 BS[8] 9.79448
R427 BS[8] BS[8].n3 9.53757
R428 BS[8] BS[8].n4 5.6005
R429 x5.A.n1 x5.A.t0 274.793
R430 x5.A.n2 x5.A.t5 232.214
R431 x5.A.n1 x5.A.n0 205.28
R432 x5.A x5.A.t1 169.452
R433 x5.A.n2 x5.A.t4 159.915
R434 x5.A.n3 x5.A.n2 152
R435 x5.A.n4 x5.A.n1 58.4086
R436 x5.A.n0 x5.A.t2 26.5955
R437 x5.A.n0 x5.A.t3 26.5955
R438 x5.A.n4 x5.A.n3 23.9621
R439 x5.A x5.A.n4 9.07762
R440 x5.A.n3 x5.A 0.970197
R441 a_5559_n3687.t0 a_5559_n3687.t1 49.8467
R442 a_5643_n3687.t0 a_5643_n3687.t1 60.9236
R443 b[7].n1 b[7].t0 230.155
R444 b[7].n0 b[7].t1 229.369
R445 b[7].n1 b[7].t3 157.856
R446 b[7].n0 b[7].t2 157.07
R447 b[7].n4 b[7].n0 152.238
R448 b[7].n2 b[7].n1 152
R449 b[7].n3 b[7].n2 19.8154
R450 b[7].n4 b[7].n3 17.1483
R451 b[7] b[7].n4 5.68939
R452 b[7].n2 b[7] 4.39453
R453 b[7].n3 b[7] 0.15675
R454 bb[7].n0 bb[7].t1 241.536
R455 bb[7].n0 bb[7].t0 169.237
R456 bb[7] bb[7].n0 154.744
R457 a_6287_n3687.t0 a_6287_n3687.t1 60.9236
R458 a_4919_n2823.t0 a_4919_n2823.t1 49.8467
R459 x1.Y.n3 x1.Y.t4 232.214
R460 x1.Y.n5 x1.Y.n2 191.1
R461 x1.Y.n3 x1.Y.t3 159.915
R462 x1.Y.n4 x1.Y.n3 155.097
R463 x1.Y.n0 x1.Y.t1 132.067
R464 x1.Y x1.Y.n5 33.6787
R465 x1.Y.n5 x1.Y.n4 33.6331
R466 x1.Y.n2 x1.Y.t2 26.5955
R467 x1.Y.n2 x1.Y.t0 26.5955
R468 x1.Y.n1 x1.Y.n0 4.15748
R469 x1.Y x1.Y.n1 3.76521
R470 x1.Y.n4 x1.Y 1.65211
R471 x1.Y.n0 x1.Y 1.17559
R472 x1.Y.n1 x1.Y 0.921363
R473 a_5835_n2823.t0 a_5835_n2823.t1 49.8467
R474 a_5919_n2823.t0 a_5919_n2823.t1 60.9236
R475 b[8].n5 b[8].t2 230.155
R476 b[8].n1 b[8].t3 229.369
R477 b[8].n0 b[8].t5 229.369
R478 b[8] b[8].n0 157.927
R479 b[8].n5 b[8].t1 157.856
R480 b[8].n1 b[8].t0 157.07
R481 b[8].n0 b[8].t4 157.07
R482 b[8].n2 b[8].n1 153.423
R483 b[8].n6 b[8].n5 152
R484 b[8].n4 b[8].n3 17.3956
R485 b[8].n3 b[8].n2 15.3266
R486 b[8].n4 b[8] 13.1418
R487 b[8].n6 b[8].n4 7.9365
R488 b[8].n2 b[8] 4.5042
R489 b[8] b[8].n6 2.3045
R490 b[8].n3 b[8] 0.3755
R491 bb[6].n0 bb[6].t0 232.214
R492 bb[6].n0 bb[6].t1 159.915
R493 bb[6].n1 bb[6].n0 152
R494 bb[6].n1 bb[6] 19.2919
R495 bb[6] bb[6].n1 2.27147
R496 a_4919_n3687.t0 a_4919_n3687.t1 49.8467
R497 a_5563_n2823.t0 a_5563_n2823.t1 49.8467
R498 a_5195_n2823.t0 a_5195_n2823.t1 49.8467
R499 BSB[8].n0 BSB[8].t1 235.56
R500 BSB[8] BSB[8].t0 161.238
R501 BSB[8] BSB[8].n0 2.22659
R502 BSB[8].n0 BSB[8] 1.55202
C0 x1.Y BS[9] 0.21208f
C1 BSB[8] x5.A 0.04536f
C2 x3.Y x1.Y 0.01808f
C3 bb[6] x5.A 0.10573f
C4 b[9] b[6] 0.33349f
C5 x5.C x5.A 0.01033f
C6 x6.Y x5.A 0.10653f
C7 bb[8] VDD 0.45166f
C8 bb[7] x5.A 0.18679f
C9 BSB[9] VDD 0.15384f
C10 bb[6] a_6493_n3695# 0.02425f
C11 bb[8] BSB[8] 0.03453f
C12 bb[6] bb[8] 0.03693f
C13 x3.Y b[9] 0.05879f
C14 a_6493_n3151# VDD 0.04572f
C15 BS[8] VDD 0.54097f
C16 x3.Y BS[9] 0.09519f
C17 bb[7] bb[8] 1.1306f
C18 bb[6] a_6493_n3151# 0.0131f
C19 a_6493_n3429# VDD 0.03791f
C20 BSB[8] BS[8] 0.05836f
C21 a_6493_n3429# bb[6] 0.01008f
C22 VDD x2.Y 0.36565f
C23 x5.C BS[8] 0.08178f
C24 x6.Y BS[8] 0.19996f
C25 b[7] x2.Y 0.04684f
C26 a_6493_n3695# x5.A 0.01593f
C27 b[7] VDD 0.2427f
C28 BSB[9] BS[9] 0.06052f
C29 BSB[8] VDD 0.18859f
C30 x1.Y x2.Y 0.61284f
C31 bb[8] x5.A 0.20635f
C32 bb[6] VDD 0.18724f
C33 m2_7109_n3782# bb[8] 0.62241f
C34 x1.Y VDD 1.0624f
C35 x1.Y b[7] 0.04148f
C36 b[8] VDD 0.40233f
C37 x5.C VDD 0.33964f
C38 x6.Y VDD 0.28029f
C39 b[8] b[7] 1.00256f
C40 x6.Y b[7] 0.06263f
C41 bb[7] VDD 0.12669f
C42 b[6] x2.Y 0.17651f
C43 b[6] VDD 0.93409f
C44 b[8] x1.Y 0.05296f
C45 x5.A BS[8] 0.23849f
C46 bb[7] bb[6] 1.04818f
C47 b[9] x2.Y 0.13356f
C48 b[6] b[7] 0.74556f
C49 x5.C b[8] 0.0538f
C50 x6.Y b[8] 0.15112f
C51 a_6493_n3429# x5.A 0.02202f
C52 x5.C x6.Y 0.29614f
C53 b[9] VDD 0.42196f
C54 b[9] b[7] 0.71105f
C55 x1.Y b[6] 0.10858f
C56 BS[9] x2.Y 0.2128f
C57 x3.Y x2.Y 0.2455f
C58 b[8] b[6] 0.74843f
C59 x5.C b[6] 0.20914f
C60 x6.Y b[6] 0.041f
C61 BSB[9] a_6493_n3151# 0.0174f
C62 BS[9] VDD 0.52855f
C63 x3.Y VDD 0.33402f
C64 x1.Y b[9] 0.13525f
C65 BS[9] b[7] 0.01229f
C66 bb[8] BS[8] 0.03947f
C67 x5.A VDD 0.42019f
C68 x3.Y b[7] 0.26557f
C69 m2_7109_n3782# VDD 0.68104f
C70 b[8] b[9] 0.94215f
C71 x5.C b[9] 0.0149f
C72 a_6493_n3429# bb[8] 0.02963f
C73 BSB[9] a_6493_n2823# 0.01166f
C74 BSB[8] GND 0.12672f
C75 bb[6] GND 0.46132f
C76 bb[7] GND 0.26121f
C77 bb[8] GND 0.31166f
C78 BS[8] GND 0.37465f
C79 BSB[9] GND 0.15857f
C80 BS[9] GND 0.6073f
C81 b[7] GND 1.21269f
C82 b[6] GND 1.09514f
C83 b[9] GND 0.70667f
C84 b[8] GND 0.62706f
C85 VDD GND 6.64227f
C86 m2_7109_n3782# GND 0.10886f $ **FLOATING
C87 a_6493_n3695# GND 0.03465f $ **FLOATING
C88 x5.A GND 0.53369f
C89 x6.Y GND 0.71195f
C90 x5.C GND 0.37678f
C91 a_6493_n3151# GND 0.01647f $ **FLOATING
C92 a_6493_n2823# GND 0.03495f $ **FLOATING
C93 x1.Y GND 0.34394f
C94 x2.Y GND 0.31806f
C95 x3.Y GND 0.33953f
.ends

