magic
tech sky130A
magscale 1 2
timestamp 1743275510
<< pwell >>
rect -201 -671 201 671
<< psubdiff >>
rect -165 601 -69 635
rect 69 601 165 635
rect -165 539 -131 601
rect 131 539 165 601
rect -165 -601 -131 -539
rect 131 -601 165 -539
rect -165 -635 -69 -601
rect 69 -635 165 -601
<< psubdiffcont >>
rect -69 601 69 635
rect -165 -539 -131 539
rect 131 -539 165 539
rect -69 -635 69 -601
<< xpolycontact >>
rect -35 73 35 505
rect -35 -505 35 -73
<< xpolyres >>
rect -35 -73 35 73
<< locali >>
rect -165 601 -69 635
rect 69 601 165 635
rect -165 539 -131 601
rect 131 539 165 601
rect -165 -601 -131 -539
rect 131 -601 165 -539
rect -165 -635 -69 -601
rect 69 -635 165 -601
<< viali >>
rect -19 90 19 487
rect -19 -487 19 -90
<< metal1 >>
rect -25 487 25 499
rect -25 90 -19 487
rect 19 90 25 487
rect -25 78 25 90
rect -25 -90 25 -78
rect -25 -487 -19 -90
rect 19 -487 25 -90
rect -25 -499 25 -487
<< properties >>
string FIXED_BBOX -148 -618 148 618
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.889 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 6.155k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
