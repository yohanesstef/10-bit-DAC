magic
tech sky130A
magscale 1 2
timestamp 1749220931
<< error_p >>
rect -174 -140 -144 72
rect -108 -74 -78 6
rect 78 -74 108 6
rect -108 -78 108 -74
rect 144 -140 174 72
rect -174 -144 174 -140
<< nwell >>
rect -144 -140 144 106
<< mvpmos >>
rect -50 -78 50 6
<< mvpdiff >>
rect -108 -6 -50 6
rect -108 -66 -96 -6
rect -62 -66 -50 -6
rect -108 -78 -50 -66
rect 50 -6 108 6
rect 50 -66 62 -6
rect 96 -66 108 -6
rect 50 -78 108 -66
<< mvpdiffc >>
rect -96 -66 -62 -6
rect 62 -66 96 -6
<< poly >>
rect -50 87 50 103
rect -50 53 -34 87
rect 34 53 50 87
rect -50 6 50 53
rect -50 -104 50 -78
<< polycont >>
rect -34 53 34 87
<< locali >>
rect -50 53 -34 87
rect 34 53 50 87
rect -96 -6 -62 10
rect -96 -82 -62 -66
rect 62 -6 96 10
rect 62 -82 96 -66
<< viali >>
rect -34 53 34 87
rect -96 -66 -62 -6
rect 62 -66 96 -6
<< metal1 >>
rect -46 87 46 93
rect -46 53 -34 87
rect 34 53 46 87
rect -46 47 46 53
rect -102 -6 -56 6
rect -102 -66 -96 -6
rect -62 -66 -56 -6
rect -102 -78 -56 -66
rect 56 -6 102 6
rect 56 -66 62 -6
rect 96 -66 102 -6
rect 56 -78 102 -66
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 0.50 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
