magic
tech sky130A
magscale 1 2
timestamp 1750150351
<< nwell >>
rect 1 -1290 1691 1392
<< mvnsubdiffcont >>
rect 140 1279 1552 1313
rect 80 -1151 114 1253
rect 1578 -1151 1612 1253
rect 140 -1211 1552 -1177
<< viali >>
rect 80 1279 140 1313
rect 140 1279 1552 1313
rect 1552 1279 1612 1313
rect 80 1253 114 1279
rect 80 -1151 114 1253
rect 80 -1177 114 -1151
rect 1578 1253 1612 1279
rect 1578 -1151 1612 1253
rect 1578 -1177 1612 -1151
rect 80 -1211 140 -1177
rect 140 -1211 1552 -1177
rect 1552 -1211 1612 -1177
<< metal1 >>
rect 506 141 552 169
rect 1140 141 1186 169
rect 249 81 701 141
rect 989 81 1186 141
rect 249 -961 309 81
rect 249 -1027 309 -1021
rect 337 -39 701 21
rect 990 -39 1186 21
rect 337 -961 397 -39
rect 506 -67 552 -39
rect 1140 -67 1186 -39
rect 337 -1027 397 -1021
<< via1 >>
rect 249 -1021 309 -961
rect 337 -1021 397 -961
<< metal2 >>
rect 249 -961 309 -955
rect 249 -1224 309 -1021
rect 337 -961 397 -955
rect 337 -1224 397 -1021
use cross_pair  cross_pair_0
timestamp 1750150351
transform -1 0 37104 0 -1 1996
box 36114 1855 36403 2035
use fc_pmos1_2  fc_pmos1_2_0
timestamp 1750009003
transform -1 0 1251 0 1 113
box -440 -128 1250 1279
use fc_pmos1_2  fc_pmos1_2_1
timestamp 1750009003
transform -1 0 1251 0 -1 -11
box -440 -128 1250 1279
<< end >>
