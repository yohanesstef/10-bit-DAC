* PEX produced on Sun Mar 30 19:20:10 +07 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from res_seg_3.ext - technology: sky130A

.subckt res_seg_3-lay v8 v7 v6 v5 v4 v3 v2 v1 v0 gnd
X0 v6.t1 v5.t1 gnd.t6 sky130_fd_pr__res_xhigh_po_0p35 l=0.85
X1 v8.t0 v7.t1 gnd.t7 sky130_fd_pr__res_xhigh_po_0p35 l=0.95
X2 v4.t1 v5.t0 gnd.t3 sky130_fd_pr__res_xhigh_po_0p35 l=0.81
X3 v6.t0 v7.t0 gnd.t0 sky130_fd_pr__res_xhigh_po_0p35 l=0.89
X4 v4.t0 v3.t0 gnd.t1 sky130_fd_pr__res_xhigh_po_0p35 l=0.77
X5 v2.t0 v1.t0 gnd.t2 sky130_fd_pr__res_xhigh_po_0p35 l=0.72
X6 v2.t1 v3.t1 gnd.t4 sky130_fd_pr__res_xhigh_po_0p35 l=0.74
X7 v0.t0 v1.t1 gnd.t5 sky130_fd_pr__res_xhigh_po_0p35 l=0.69
R0 v6.n0 v6.t0 45.1448
R1 v6.n0 v6.t1 42.3691
R2 v6 v6.n0 0.0248056
R3 v5 v5.t1 45.0331
R4 v5 v5.t0 42.5516
R5 gnd.n33 gnd.n25 4374.56
R6 gnd.n29 gnd.n25 4374.56
R7 gnd.n33 gnd.n26 4374.56
R8 gnd.n40 gnd.n22 4339.79
R9 gnd.n36 gnd.n22 4339.79
R10 gnd.n40 gnd.n23 4339.79
R11 gnd.n36 gnd.n23 4339.79
R12 gnd.n47 gnd.n19 4316.62
R13 gnd.n43 gnd.n19 4316.62
R14 gnd.n47 gnd.n20 4316.62
R15 gnd.n43 gnd.n20 4316.62
R16 gnd.n54 gnd.n16 4293.44
R17 gnd.n50 gnd.n16 4293.44
R18 gnd.n54 gnd.n17 4293.44
R19 gnd.n50 gnd.n17 4293.44
R20 gnd.n61 gnd.n13 4270.26
R21 gnd.n57 gnd.n13 4270.26
R22 gnd.n61 gnd.n14 4270.26
R23 gnd.n57 gnd.n14 4270.26
R24 gnd.n68 gnd.n10 4252.88
R25 gnd.n64 gnd.n10 4252.88
R26 gnd.n68 gnd.n11 4252.88
R27 gnd.n64 gnd.n11 4252.88
R28 gnd.n75 gnd.n7 4241.29
R29 gnd.n71 gnd.n7 4241.29
R30 gnd.n75 gnd.n8 4241.29
R31 gnd.n71 gnd.n8 4241.29
R32 gnd.n78 gnd.n2 4223.91
R33 gnd.n5 gnd.n3 4223.91
R34 gnd.n78 gnd.n3 4223.91
R35 gnd.n77 gnd.t5 480.945
R36 gnd.n76 gnd.t2 480.945
R37 gnd.n70 gnd.t2 480.945
R38 gnd.n69 gnd.t4 480.945
R39 gnd.n63 gnd.t4 480.945
R40 gnd.n62 gnd.t1 480.945
R41 gnd.n56 gnd.t1 480.945
R42 gnd.n55 gnd.t3 480.945
R43 gnd.n49 gnd.t3 480.945
R44 gnd.n48 gnd.t6 480.945
R45 gnd.n42 gnd.t6 480.945
R46 gnd.n41 gnd.t0 480.945
R47 gnd.n35 gnd.t0 480.945
R48 gnd.n34 gnd.t7 480.945
R49 gnd.n29 gnd.n28 436.656
R50 gnd.n6 gnd.n5 436.07
R51 gnd.n77 gnd.n76 344.462
R52 gnd.n70 gnd.n69 344.462
R53 gnd.n63 gnd.n62 344.462
R54 gnd.n56 gnd.n55 344.462
R55 gnd.n49 gnd.n48 344.462
R56 gnd.n42 gnd.n41 344.462
R57 gnd.n35 gnd.n34 344.462
R58 gnd.n73 gnd.n8 292.5
R59 gnd.n8 gnd.t2 292.5
R60 gnd.n9 gnd.n7 292.5
R61 gnd.n7 gnd.t2 292.5
R62 gnd.n66 gnd.n11 292.5
R63 gnd.n11 gnd.t4 292.5
R64 gnd.n12 gnd.n10 292.5
R65 gnd.n10 gnd.t4 292.5
R66 gnd.n59 gnd.n14 292.5
R67 gnd.n14 gnd.t1 292.5
R68 gnd.n15 gnd.n13 292.5
R69 gnd.n13 gnd.t1 292.5
R70 gnd.n52 gnd.n17 292.5
R71 gnd.n17 gnd.t3 292.5
R72 gnd.n18 gnd.n16 292.5
R73 gnd.n16 gnd.t3 292.5
R74 gnd.n45 gnd.n20 292.5
R75 gnd.n20 gnd.t6 292.5
R76 gnd.n21 gnd.n19 292.5
R77 gnd.n19 gnd.t6 292.5
R78 gnd.n38 gnd.n23 292.5
R79 gnd.n23 gnd.t0 292.5
R80 gnd.n24 gnd.n22 292.5
R81 gnd.n22 gnd.t0 292.5
R82 gnd.n31 gnd.n26 292.5
R83 gnd.n27 gnd.n25 292.5
R84 gnd.n25 gnd.t7 292.5
R85 gnd.n3 gnd.n1 292.5
R86 gnd.t5 gnd.n3 292.5
R87 gnd.n2 gnd.n0 292.5
R88 gnd.n32 gnd.n27 284.236
R89 gnd.n30 gnd.n27 284.236
R90 gnd.n32 gnd.n31 284.236
R91 gnd.n31 gnd.n30 284.236
R92 gnd.n39 gnd.n24 281.976
R93 gnd.n37 gnd.n24 281.976
R94 gnd.n39 gnd.n38 281.976
R95 gnd.n38 gnd.n37 281.976
R96 gnd.n46 gnd.n21 280.471
R97 gnd.n44 gnd.n21 280.471
R98 gnd.n46 gnd.n45 280.471
R99 gnd.n45 gnd.n44 280.471
R100 gnd.n53 gnd.n18 278.966
R101 gnd.n51 gnd.n18 278.966
R102 gnd.n53 gnd.n52 278.966
R103 gnd.n52 gnd.n51 278.966
R104 gnd.n60 gnd.n15 277.459
R105 gnd.n58 gnd.n15 277.459
R106 gnd.n60 gnd.n59 277.459
R107 gnd.n59 gnd.n58 277.459
R108 gnd.n67 gnd.n12 276.329
R109 gnd.n65 gnd.n12 276.329
R110 gnd.n67 gnd.n66 276.329
R111 gnd.n66 gnd.n65 276.329
R112 gnd.n74 gnd.n9 275.577
R113 gnd.n72 gnd.n9 275.577
R114 gnd.n74 gnd.n73 275.577
R115 gnd.n73 gnd.n72 275.577
R116 gnd.n79 gnd.n1 274.447
R117 gnd.n4 gnd.n1 274.447
R118 gnd.n4 gnd.n0 274.447
R119 gnd gnd.n79 248.471
R120 gnd.n28 gnd.n26 246.803
R121 gnd.n6 gnd.n2 245.316
R122 gnd.n72 gnd.n71 39.0005
R123 gnd.n71 gnd.n70 39.0005
R124 gnd.n75 gnd.n74 39.0005
R125 gnd.n76 gnd.n75 39.0005
R126 gnd.n65 gnd.n64 39.0005
R127 gnd.n64 gnd.n63 39.0005
R128 gnd.n68 gnd.n67 39.0005
R129 gnd.n69 gnd.n68 39.0005
R130 gnd.n79 gnd.n78 39.0005
R131 gnd.n78 gnd.n77 39.0005
R132 gnd.n5 gnd.n4 39.0005
R133 gnd.n58 gnd.n57 36.563
R134 gnd.n57 gnd.n56 36.563
R135 gnd.n61 gnd.n60 36.563
R136 gnd.n62 gnd.n61 36.563
R137 gnd.n51 gnd.n50 36.563
R138 gnd.n50 gnd.n49 36.563
R139 gnd.n54 gnd.n53 36.563
R140 gnd.n55 gnd.n54 36.563
R141 gnd.n44 gnd.n43 36.563
R142 gnd.n43 gnd.n42 36.563
R143 gnd.n47 gnd.n46 36.563
R144 gnd.n48 gnd.n47 36.563
R145 gnd.n37 gnd.n36 36.563
R146 gnd.n36 gnd.n35 36.563
R147 gnd.n40 gnd.n39 36.563
R148 gnd.n41 gnd.n40 36.563
R149 gnd.n30 gnd.n29 36.563
R150 gnd.n33 gnd.n32 36.563
R151 gnd.n34 gnd.n33 36.563
R152 gnd.t5 gnd.n6 30.1982
R153 gnd.n28 gnd.t7 29.1975
R154 gnd gnd.n0 25.977
R155 v8 v8.t0 42.3816
R156 v7.n0 v7.t1 45.1181
R157 v7.n0 v7.t0 42.5516
R158 v7 v7.n0 0.0355
R159 v4 v4.t1 44.773
R160 v4 v4.t0 42.3916
R161 v3 v3.t0 44.9981
R162 v3 v3.t1 42.5566
R163 v2 v2.t1 44.763
R164 v2 v2.t0 42.3716
R165 v1 v1.t0 44.8731
R166 v1 v1.t1 42.5516
R167 v0 v0.t0 42.37
C0 v6 v8 0.04591f
C1 v6 v7 0.02147f
C2 v4 v5 0.02349f
C3 v7 v8 0.02005f
C4 v3 v2 0.02557f
C5 v1 v2 0.02625f
C6 v1 v3 0.04717f
C7 v6 v5 0.02243f
C8 v5 v7 0.04722f
C9 v3 v5 0.04717f
C10 v4 v6 0.04636f
C11 v0 v2 0.04659f
C12 v4 v2 0.04659f
C13 v4 v3 0.02463f
C14 v1 v0 0.02715f
C15 v0 gnd 0.53321f
C16 v1 gnd 1.18148f
C17 v2 gnd 1.13855f
C18 v3 gnd 1.13772f
C19 v4 gnd 1.14077f
C20 v5 gnd 1.13929f
C21 v6 gnd 1.14618f
C22 v7 gnd 1.19088f
C23 v8 gnd 0.53599f
.ends

