magic
tech sky130A
magscale 1 2
timestamp 1749033013
<< psubdiff >>
rect 991 5238 4501 5298
rect 991 -11001 1051 5238
rect 4441 -11001 4501 5238
rect 991 -11061 4501 -11001
<< metal3 >>
rect 4155 -11001 4355 -10905
<< properties >>
string FIXED_BBOX -254 -929 254 929
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 4 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 5.94k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
