magic
tech sky130A
magscale 1 2
timestamp 1750019162
<< error_s >>
rect 2557 1312 2584 1322
rect 2531 1252 2584 1312
rect 2557 1242 2584 1252
rect 2585 1312 2612 1322
rect 4062 1312 4089 1322
rect 2585 1252 2638 1312
rect 4036 1252 4089 1312
rect 2585 1242 2612 1252
rect 4062 1242 4089 1252
rect 4090 1312 4117 1322
rect 5567 1312 5594 1322
rect 4090 1252 4143 1312
rect 5541 1252 5594 1312
rect 4090 1242 4117 1252
rect 5567 1242 5594 1252
rect 5595 1312 5622 1322
rect 7072 1312 7099 1322
rect 5595 1252 5648 1312
rect 7046 1252 7099 1312
rect 5595 1242 5622 1252
rect 7072 1242 7099 1252
rect 7100 1312 7127 1322
rect 8577 1312 8604 1322
rect 7100 1252 7153 1312
rect 8551 1252 8604 1312
rect 7100 1242 7127 1252
rect 8577 1242 8604 1252
rect 8605 1312 8632 1322
rect 8605 1252 8658 1312
rect 8605 1242 8632 1252
rect 2557 1154 2584 1214
rect 2585 1154 2612 1214
rect 4062 1154 4089 1214
rect 4090 1154 4117 1214
rect 5567 1154 5594 1214
rect 5595 1154 5622 1214
rect 7072 1154 7099 1214
rect 7100 1154 7127 1214
rect 8577 1154 8604 1214
rect 8605 1154 8632 1214
rect 2557 226 2584 286
rect 2585 226 2612 286
rect 4062 226 4089 286
rect 4090 226 4117 286
rect 5567 226 5594 286
rect 5595 226 5622 286
rect 7072 226 7099 286
rect 7100 226 7127 286
rect 8577 226 8604 286
rect 8605 226 8632 286
rect 2557 188 2584 198
rect 2531 128 2584 188
rect 2557 118 2584 128
rect 2585 188 2612 198
rect 4062 188 4089 198
rect 2585 128 2638 188
rect 4036 128 4089 188
rect 2585 118 2612 128
rect 4062 118 4089 128
rect 4090 188 4117 198
rect 5567 188 5594 198
rect 4090 128 4143 188
rect 5541 128 5594 188
rect 4090 118 4117 128
rect 5567 118 5594 128
rect 5595 188 5622 198
rect 7072 188 7099 198
rect 5595 128 5648 188
rect 7046 128 7099 188
rect 5595 118 5622 128
rect 7072 118 7099 128
rect 7100 188 7127 198
rect 8577 188 8604 198
rect 7100 128 7153 188
rect 8551 128 8604 188
rect 7100 118 7127 128
rect 8577 118 8604 128
rect 8605 188 8632 198
rect 8605 128 8658 188
rect 8605 118 8632 128
rect 2557 30 2584 90
rect 2585 30 2612 90
rect 4062 30 4089 90
rect 4090 30 4117 90
rect 5567 30 5594 90
rect 5595 30 5622 90
rect 7072 30 7099 90
rect 7100 30 7127 90
rect 8577 30 8604 90
rect 8605 30 8632 90
rect 2557 -898 2584 -838
rect 2585 -898 2612 -838
rect 4062 -898 4089 -838
rect 4090 -898 4117 -838
rect 5567 -898 5594 -838
rect 5595 -898 5622 -838
rect 7072 -898 7099 -838
rect 7100 -898 7127 -838
rect 8577 -898 8604 -838
rect 8605 -898 8632 -838
rect 2557 -936 2584 -926
rect 2531 -969 2584 -936
rect 1091 -996 2584 -969
rect 1117 -1006 2584 -996
rect 2585 -936 2612 -926
rect 4062 -936 4089 -926
rect 2585 -969 2638 -936
rect 4036 -969 4089 -936
rect 2585 -1006 4089 -969
rect 4090 -936 4117 -926
rect 5567 -936 5594 -926
rect 4090 -969 4143 -936
rect 5541 -969 5594 -936
rect 4090 -1006 5594 -969
rect 5595 -936 5622 -926
rect 7072 -936 7099 -926
rect 5595 -969 5648 -936
rect 7046 -969 7099 -936
rect 5595 -1006 7099 -969
rect 7100 -936 7127 -926
rect 8577 -936 8604 -926
rect 7100 -969 7153 -936
rect 8551 -969 8604 -936
rect 7100 -1006 8604 -969
rect 8605 -936 8632 -926
rect 8605 -969 8658 -936
rect 8605 -1006 10109 -969
rect 1145 -1050 2649 -1013
rect 2596 -1083 2649 -1050
rect 2622 -1093 2649 -1083
rect 2650 -1050 4154 -1013
rect 2650 -1083 2703 -1050
rect 4101 -1083 4154 -1050
rect 2650 -1093 2677 -1083
rect 4127 -1093 4154 -1083
rect 4155 -1050 5659 -1013
rect 4155 -1083 4208 -1050
rect 5606 -1083 5659 -1050
rect 4155 -1093 4182 -1083
rect 5632 -1093 5659 -1083
rect 5660 -1050 7164 -1013
rect 5660 -1083 5713 -1050
rect 7111 -1083 7164 -1050
rect 5660 -1093 5687 -1083
rect 7137 -1093 7164 -1083
rect 7165 -1050 8669 -1013
rect 7165 -1083 7218 -1050
rect 8616 -1083 8669 -1050
rect 7165 -1093 7192 -1083
rect 8642 -1093 8669 -1083
rect 8670 -1023 10137 -1013
rect 8670 -1050 10163 -1023
rect 8670 -1083 8723 -1050
rect 8670 -1093 8697 -1083
rect 2622 -1181 2649 -1121
rect 2650 -1181 2677 -1121
rect 4127 -1181 4154 -1121
rect 4155 -1181 4182 -1121
rect 5632 -1181 5659 -1121
rect 5660 -1181 5687 -1121
rect 7137 -1181 7164 -1121
rect 7165 -1181 7192 -1121
rect 8642 -1181 8669 -1121
rect 8670 -1181 8697 -1121
rect 2622 -2109 2649 -2049
rect 2650 -2109 2677 -2049
rect 4127 -2109 4154 -2049
rect 4155 -2109 4182 -2049
rect 5632 -2109 5659 -2049
rect 5660 -2109 5687 -2049
rect 7137 -2109 7164 -2049
rect 7165 -2109 7192 -2049
rect 8642 -2109 8669 -2049
rect 8670 -2109 8697 -2049
rect 2622 -2147 2649 -2137
rect 2596 -2207 2649 -2147
rect 2622 -2217 2649 -2207
rect 2650 -2147 2677 -2137
rect 4127 -2147 4154 -2137
rect 2650 -2207 2703 -2147
rect 4101 -2207 4154 -2147
rect 2650 -2217 2677 -2207
rect 4127 -2217 4154 -2207
rect 4155 -2147 4182 -2137
rect 5632 -2147 5659 -2137
rect 4155 -2207 4208 -2147
rect 5606 -2207 5659 -2147
rect 4155 -2217 4182 -2207
rect 5632 -2217 5659 -2207
rect 5660 -2147 5687 -2137
rect 7137 -2147 7164 -2137
rect 5660 -2207 5713 -2147
rect 7111 -2207 7164 -2147
rect 5660 -2217 5687 -2207
rect 7137 -2217 7164 -2207
rect 7165 -2147 7192 -2137
rect 8642 -2147 8669 -2137
rect 7165 -2207 7218 -2147
rect 8616 -2207 8669 -2147
rect 7165 -2217 7192 -2207
rect 8642 -2217 8669 -2207
rect 8670 -2147 8697 -2137
rect 8670 -2207 8723 -2147
rect 8670 -2217 8697 -2207
rect 2622 -2305 2649 -2245
rect 2650 -2305 2677 -2245
rect 4127 -2305 4154 -2245
rect 4155 -2305 4182 -2245
rect 5632 -2305 5659 -2245
rect 5660 -2305 5687 -2245
rect 7137 -2305 7164 -2245
rect 7165 -2305 7192 -2245
rect 8642 -2305 8669 -2245
rect 8670 -2305 8697 -2245
rect 2622 -3199 2649 -3173
rect 2650 -3199 2677 -3173
rect 4127 -3199 4154 -3173
rect 4155 -3199 4182 -3173
rect 5632 -3199 5659 -3173
rect 5660 -3199 5687 -3173
rect 7137 -3199 7164 -3173
rect 7165 -3199 7192 -3173
rect 8642 -3199 8669 -3173
rect 8670 -3199 8697 -3173
rect 2622 -3209 2679 -3199
rect 4127 -3209 4184 -3199
rect 5632 -3209 5689 -3199
rect 7137 -3209 7194 -3199
rect 8642 -3209 8699 -3199
rect 1222 -3217 1455 -3209
rect 1598 -3217 1831 -3209
rect 1974 -3217 2207 -3209
rect 2350 -3217 2583 -3209
rect 2598 -3217 2705 -3209
rect 2727 -3217 2960 -3209
rect 3103 -3217 3336 -3209
rect 3479 -3217 3712 -3209
rect 3855 -3217 4088 -3209
rect 4103 -3217 4210 -3209
rect 4232 -3217 4465 -3209
rect 4608 -3217 4841 -3209
rect 4984 -3217 5217 -3209
rect 5360 -3217 5593 -3209
rect 5608 -3217 5715 -3209
rect 5737 -3217 5970 -3209
rect 6113 -3217 6346 -3209
rect 6489 -3217 6722 -3209
rect 6865 -3217 7098 -3209
rect 7113 -3217 7220 -3209
rect 7242 -3217 7475 -3209
rect 7618 -3217 7851 -3209
rect 7994 -3217 8227 -3209
rect 8370 -3217 8603 -3209
rect 8618 -3217 8725 -3209
rect 8747 -3217 8980 -3209
rect 9123 -3217 9356 -3209
rect 9499 -3217 9732 -3209
rect 9875 -3217 10108 -3209
rect 1147 -3233 10176 -3217
rect 1147 -3251 2651 -3233
rect 2652 -3251 4156 -3233
rect 4157 -3251 5661 -3233
rect 5662 -3251 7166 -3233
rect 7167 -3251 8671 -3233
rect 8672 -3251 10176 -3233
rect 1147 -3261 10176 -3251
rect 1147 -3269 2651 -3261
rect 2652 -3269 4156 -3261
rect 4157 -3269 5661 -3261
rect 5662 -3269 7166 -3261
rect 7167 -3269 8671 -3261
rect 8672 -3269 10176 -3261
rect 1145 -3307 2649 -3271
rect 2650 -3307 4154 -3271
rect 4155 -3307 5659 -3271
rect 5660 -3307 7164 -3271
rect 7165 -3307 8669 -3271
rect 8670 -3307 10174 -3271
rect 1145 -3323 10174 -3307
rect 1224 -3331 1457 -3323
rect 1600 -3331 1833 -3323
rect 1976 -3331 2209 -3323
rect 2352 -3331 2585 -3323
rect 2596 -3331 2703 -3323
rect 2729 -3331 2962 -3323
rect 3105 -3331 3338 -3323
rect 3481 -3331 3714 -3323
rect 3857 -3331 4090 -3323
rect 4101 -3331 4208 -3323
rect 4234 -3331 4467 -3323
rect 4610 -3331 4843 -3323
rect 4986 -3331 5219 -3323
rect 5362 -3331 5595 -3323
rect 5606 -3331 5713 -3323
rect 5739 -3331 5972 -3323
rect 6115 -3331 6348 -3323
rect 6491 -3331 6724 -3323
rect 6867 -3331 7100 -3323
rect 7111 -3331 7218 -3323
rect 7244 -3331 7477 -3323
rect 7620 -3331 7853 -3323
rect 7996 -3331 8229 -3323
rect 8372 -3331 8605 -3323
rect 8616 -3331 8723 -3323
rect 8749 -3331 8982 -3323
rect 9125 -3331 9358 -3323
rect 9501 -3331 9734 -3323
rect 9877 -3331 10110 -3323
rect 2622 -3341 2679 -3331
rect 4127 -3341 4184 -3331
rect 5632 -3341 5689 -3331
rect 7137 -3341 7194 -3331
rect 8642 -3341 8699 -3331
rect 2624 -3367 2651 -3341
rect 2652 -3367 2679 -3341
rect 4129 -3367 4156 -3341
rect 4157 -3367 4184 -3341
rect 5634 -3367 5661 -3341
rect 5662 -3367 5689 -3341
rect 7139 -3367 7166 -3341
rect 7167 -3367 7194 -3341
rect 8644 -3367 8671 -3341
rect 8672 -3367 8699 -3341
rect 2624 -4295 2651 -4235
rect 2652 -4295 2679 -4235
rect 4129 -4295 4156 -4235
rect 4157 -4295 4184 -4235
rect 5634 -4295 5661 -4235
rect 5662 -4295 5689 -4235
rect 7139 -4295 7166 -4235
rect 7167 -4295 7194 -4235
rect 8644 -4295 8671 -4235
rect 8672 -4295 8699 -4235
rect 2624 -4333 2651 -4323
rect 2598 -4393 2651 -4333
rect 2624 -4403 2651 -4393
rect 2652 -4333 2679 -4323
rect 4129 -4333 4156 -4323
rect 2652 -4393 2705 -4333
rect 4103 -4393 4156 -4333
rect 2652 -4403 2679 -4393
rect 4129 -4403 4156 -4393
rect 4157 -4333 4184 -4323
rect 5634 -4333 5661 -4323
rect 4157 -4393 4210 -4333
rect 5608 -4393 5661 -4333
rect 4157 -4403 4184 -4393
rect 5634 -4403 5661 -4393
rect 5662 -4333 5689 -4323
rect 7139 -4333 7166 -4323
rect 5662 -4393 5715 -4333
rect 7113 -4393 7166 -4333
rect 5662 -4403 5689 -4393
rect 7139 -4403 7166 -4393
rect 7167 -4333 7194 -4323
rect 8644 -4333 8671 -4323
rect 7167 -4393 7220 -4333
rect 8618 -4393 8671 -4333
rect 7167 -4403 7194 -4393
rect 8644 -4403 8671 -4393
rect 8672 -4333 8699 -4323
rect 8672 -4393 8725 -4333
rect 8672 -4403 8699 -4393
rect 2624 -4491 2651 -4431
rect 2652 -4491 2679 -4431
rect 4129 -4491 4156 -4431
rect 4157 -4491 4184 -4431
rect 5634 -4491 5661 -4431
rect 5662 -4491 5689 -4431
rect 7139 -4491 7166 -4431
rect 7167 -4491 7194 -4431
rect 8644 -4491 8671 -4431
rect 8672 -4491 8699 -4431
rect 2624 -5419 2651 -5359
rect 2652 -5419 2679 -5359
rect 4129 -5419 4156 -5359
rect 4157 -5419 4184 -5359
rect 5634 -5419 5661 -5359
rect 5662 -5419 5689 -5359
rect 7139 -5419 7166 -5359
rect 7167 -5419 7194 -5359
rect 8644 -5419 8671 -5359
rect 8672 -5419 8699 -5359
rect 2624 -5457 2651 -5447
rect 2598 -5517 2651 -5457
rect 2624 -5527 2651 -5517
rect 2652 -5457 2679 -5447
rect 4129 -5457 4156 -5447
rect 2652 -5517 2705 -5457
rect 4103 -5517 4156 -5457
rect 2652 -5527 2679 -5517
rect 4129 -5527 4156 -5517
rect 4157 -5457 4184 -5447
rect 5634 -5457 5661 -5447
rect 4157 -5517 4210 -5457
rect 5608 -5517 5661 -5457
rect 4157 -5527 4184 -5517
rect 5634 -5527 5661 -5517
rect 5662 -5457 5689 -5447
rect 7139 -5457 7166 -5447
rect 5662 -5517 5715 -5457
rect 7113 -5517 7166 -5457
rect 5662 -5527 5689 -5517
rect 7139 -5527 7166 -5517
rect 7167 -5457 7194 -5447
rect 8644 -5457 8671 -5447
rect 7167 -5517 7220 -5457
rect 8618 -5517 8671 -5457
rect 7167 -5527 7194 -5517
rect 8644 -5527 8671 -5517
rect 8672 -5457 8699 -5447
rect 8672 -5517 8725 -5457
rect 8672 -5527 8699 -5517
use cm_pcell1_4_4  cm_pcell1_4_4_6
timestamp 1749895928
transform 1 0 -12 0 1 -462
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_7
timestamp 1749895928
transform 1 0 1493 0 1 -462
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_8
timestamp 1749895928
transform 1 0 2998 0 1 -462
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_9
timestamp 1749895928
transform 1 0 4503 0 1 -462
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_10
timestamp 1749895928
transform 1 0 6008 0 1 -462
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_11
timestamp 1749895928
transform 1 0 7513 0 1 -462
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_12
timestamp 1749895928
transform 1 0 53 0 1 -2797
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_13
timestamp 1749895928
transform 1 0 1558 0 1 -2797
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_14
timestamp 1749895928
transform 1 0 3063 0 1 -2797
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_15
timestamp 1749895928
transform 1 0 4568 0 1 -2797
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_16
timestamp 1749895928
transform 1 0 6073 0 1 -2797
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_17
timestamp 1749895928
transform 1 0 7578 0 1 -2797
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_18
timestamp 1749895928
transform 1 0 55 0 1 -4983
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_19
timestamp 1749895928
transform 1 0 1560 0 1 -4983
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_20
timestamp 1749895928
transform 1 0 3065 0 1 -4983
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_21
timestamp 1749895928
transform 1 0 4570 0 1 -4983
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_22
timestamp 1749895928
transform 1 0 6075 0 1 -4983
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_23
timestamp 1749895928
transform 1 0 7580 0 1 -4983
box 1026 -600 2672 1840
<< end >>
