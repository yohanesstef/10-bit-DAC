magic
tech sky130A
magscale 1 2
timestamp 1749147130
<< pwell >>
rect -307 -730 307 730
<< psubdiff >>
rect -271 660 -175 694
rect 175 660 271 694
rect -271 598 -237 660
rect 237 598 271 660
rect -271 -660 -237 -598
rect 237 -660 271 -598
rect -271 -694 -175 -660
rect 175 -694 271 -660
<< psubdiffcont >>
rect -175 660 175 694
rect -271 -598 -237 598
rect 237 -598 271 598
rect -175 -694 175 -660
<< xpolycontact >>
rect -141 132 141 564
rect -141 -564 141 -132
<< xpolyres >>
rect -141 -132 141 132
<< locali >>
rect -271 660 -175 694
rect 175 660 271 694
rect -271 598 -237 660
rect 237 598 271 660
rect -271 -660 -237 -598
rect 237 -660 271 -598
rect -271 -694 -175 -660
rect 175 -694 271 -660
<< viali >>
rect -125 149 125 546
rect -125 -546 125 -149
<< metal1 >>
rect -131 546 131 558
rect -131 149 -125 546
rect 125 149 131 546
rect -131 137 131 149
rect -131 -149 131 -137
rect -131 -546 -125 -149
rect 125 -546 131 -149
rect -131 -558 131 -546
<< properties >>
string FIXED_BBOX -254 -677 254 677
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.476 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 2.36k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
