magic
tech sky130A
magscale 1 2
timestamp 1750867770
<< metal1 >>
rect 20864 2133 20870 2281
rect 21070 2133 22559 2281
rect 10756 1313 10762 1513
rect 10938 1313 11752 1513
rect 11928 1313 12742 1513
rect 12918 1313 13732 1513
rect 13908 1313 14722 1513
rect 14898 1313 15712 1513
rect 15888 1313 16702 1513
rect 16878 1313 17692 1513
rect 17868 1313 18682 1513
rect 18858 1313 19672 1513
rect 19848 1313 21142 1513
rect 9046 1081 9832 1109
rect 9045 1001 9744 1029
rect 8206 173 9656 201
rect 9056 141 9656 173
rect 9046 85 9304 113
rect 9056 53 9304 85
rect 9046 -3 9062 25
rect 9056 -35 9062 -3
rect 9122 -35 9128 25
rect 9046 -91 9216 -63
rect 9056 -123 9216 -91
rect 9056 -651 9062 -591
rect 9122 -651 9128 -591
rect 9056 -827 9062 -767
rect 9122 -827 9128 -767
rect 9056 -1059 9062 -1027
rect 9028 -1087 9062 -1059
rect 9122 -1087 9128 -1027
rect 9056 -1147 9062 -1115
rect 9027 -1175 9062 -1147
rect 9122 -1175 9128 -1115
rect 9156 -1471 9216 -123
rect 9156 -1537 9216 -1531
rect 9244 -1559 9304 53
rect 9508 25 9568 31
rect 9332 -591 9392 -585
rect 9332 -1295 9392 -651
rect 9332 -1361 9392 -1355
rect 9420 -767 9480 -761
rect 9420 -1383 9480 -827
rect 9508 -1207 9568 -35
rect 9596 -1119 9656 141
rect 9684 -1031 9744 1001
rect 9772 -943 9832 1081
rect 20697 942 20870 1090
rect 21070 942 21076 1090
rect 25348 1072 25408 1132
rect 25348 -267 25408 -207
rect 20750 -888 20870 -828
rect 21070 -888 21076 -828
rect 9772 -1009 9832 -1003
rect 9684 -1097 9744 -1091
rect 9596 -1185 9656 -1179
rect 9508 -1273 9568 -1267
rect 9420 -1449 9480 -1443
rect 9028 -1658 9062 -1598
rect 9122 -1658 9128 -1598
rect 9244 -1625 9304 -1619
rect 9028 -1663 9128 -1658
rect 9027 -1719 9062 -1691
rect 9056 -1751 9062 -1719
rect 9122 -1751 9128 -1691
rect 9784 -1779 9860 -1747
rect 9028 -1807 9860 -1779
rect 9028 -1843 9971 -1807
rect 8865 -1875 9971 -1843
rect 9860 -1876 9971 -1875
rect 5748 -2019 8596 -1959
rect 8660 -2019 12930 -1959
rect 12990 -2019 23644 -1959
rect 5754 -2107 6030 -2047
rect 6094 -2107 13018 -2047
rect 13078 -2107 23644 -2047
rect 5754 -2195 8504 -2135
rect 8568 -2195 13574 -2135
rect 13634 -2195 23644 -2135
rect 5754 -2283 5938 -2223
rect 6002 -2283 13662 -2223
rect 13722 -2283 23644 -2223
rect 5754 -2371 8412 -2311
rect 8476 -2371 14218 -2311
rect 14278 -2371 23026 -2311
rect 23086 -2371 23644 -2311
rect 5754 -2459 5846 -2399
rect 5910 -2459 14306 -2399
rect 14366 -2459 23546 -2399
rect 23606 -2459 23644 -2399
rect 5754 -2547 8320 -2487
rect 8384 -2547 14862 -2487
rect 14922 -2547 20133 -2487
rect 20193 -2547 22938 -2487
rect 22998 -2547 23644 -2487
rect 5748 -2635 5754 -2575
rect 5818 -2635 14950 -2575
rect 15010 -2635 20317 -2575
rect 20377 -2635 23224 -2575
rect 23284 -2635 23644 -2575
rect 9226 -2723 15506 -2663
rect 15566 -2723 19143 -2663
rect 19203 -2723 21602 -2663
rect 21662 -2723 23644 -2663
rect 9226 -2811 15594 -2751
rect 15654 -2811 19327 -2751
rect 19387 -2811 22122 -2751
rect 22182 -2811 23644 -2751
rect 9226 -2899 16150 -2839
rect 16210 -2899 18153 -2839
rect 18213 -2899 21514 -2839
rect 21574 -2899 23644 -2839
rect 9226 -2987 16238 -2927
rect 16298 -2987 18337 -2927
rect 18397 -2987 21800 -2927
rect 21860 -2987 23644 -2927
rect 9226 -3075 16794 -3015
rect 16854 -3075 17163 -3015
rect 17223 -3075 23644 -3015
rect 9226 -3163 16882 -3103
rect 16942 -3163 17251 -3103
rect 17311 -3163 23644 -3103
rect 9226 -3251 15974 -3191
rect 16034 -3251 17438 -3191
rect 17498 -3251 23644 -3191
rect 9226 -3339 16414 -3279
rect 16474 -3339 17526 -3279
rect 17586 -3339 23644 -3279
rect 9226 -3427 15183 -3367
rect 15243 -3427 18082 -3367
rect 18142 -3427 23644 -3367
rect 9226 -3515 15367 -3455
rect 15427 -3515 18170 -3455
rect 18230 -3515 23644 -3455
rect 9226 -3603 14042 -3543
rect 14102 -3603 18726 -3543
rect 18786 -3603 23644 -3543
rect 9226 -3691 14482 -3631
rect 14542 -3691 18814 -3631
rect 18874 -3691 23644 -3631
rect 5366 -3807 24077 -3743
rect 5366 -3903 5386 -3807
rect 5542 -3903 8688 -3807
rect 8844 -3903 22539 -3807
rect 22635 -3903 23975 -3807
rect 24071 -3903 24077 -3807
rect 5564 -4447 5570 -4351
rect 5726 -4447 8872 -4351
rect 9028 -4447 20870 -4351
rect 21070 -4447 21235 -4351
rect 21331 -4447 25275 -4351
rect 25371 -4447 25377 -4351
rect 5564 -4551 25377 -4447
<< via1 >>
rect 20870 2133 21070 2281
rect 10762 1313 10938 1513
rect 11752 1313 11928 1513
rect 12742 1313 12918 1513
rect 13732 1313 13908 1513
rect 14722 1313 14898 1513
rect 15712 1313 15888 1513
rect 16702 1313 16878 1513
rect 17692 1313 17868 1513
rect 18682 1313 18858 1513
rect 19672 1313 19848 1513
rect 9062 -35 9122 25
rect 9062 -651 9122 -591
rect 9062 -827 9122 -767
rect 9062 -1087 9122 -1027
rect 9062 -1175 9122 -1115
rect 9156 -1531 9216 -1471
rect 9508 -35 9568 25
rect 9332 -651 9392 -591
rect 9332 -1355 9392 -1295
rect 9420 -827 9480 -767
rect 20870 942 21070 1090
rect 10762 278 10938 378
rect 11752 278 11928 378
rect 12742 278 12918 378
rect 13732 278 13908 378
rect 14722 278 14898 378
rect 15712 278 15888 378
rect 16702 278 16878 378
rect 17692 278 17868 378
rect 18682 278 18858 378
rect 19672 278 19848 378
rect 20870 -888 21070 -828
rect 9772 -1003 9832 -943
rect 9684 -1091 9744 -1031
rect 9596 -1179 9656 -1119
rect 9508 -1267 9568 -1207
rect 21235 -1299 21331 -1203
rect 25275 -1299 25371 -1203
rect 9420 -1443 9480 -1383
rect 9062 -1658 9122 -1598
rect 9244 -1619 9304 -1559
rect 9062 -1751 9122 -1691
rect 22539 -1843 22635 -1747
rect 23975 -1843 24071 -1747
rect 8596 -2019 8660 -1959
rect 12930 -2019 12990 -1959
rect 6030 -2107 6094 -2047
rect 13018 -2107 13078 -2047
rect 8504 -2195 8568 -2135
rect 13574 -2195 13634 -2135
rect 5938 -2283 6002 -2223
rect 13662 -2283 13722 -2223
rect 8412 -2371 8476 -2311
rect 14218 -2371 14278 -2311
rect 23026 -2371 23086 -2311
rect 5846 -2459 5910 -2399
rect 14306 -2459 14366 -2399
rect 23546 -2459 23606 -2399
rect 8320 -2547 8384 -2487
rect 14862 -2547 14922 -2487
rect 20133 -2547 20193 -2487
rect 22938 -2547 22998 -2487
rect 5754 -2635 5818 -2575
rect 14950 -2635 15010 -2575
rect 20317 -2635 20377 -2575
rect 23224 -2635 23284 -2575
rect 15506 -2723 15566 -2663
rect 19143 -2723 19203 -2663
rect 21602 -2723 21662 -2663
rect 15594 -2811 15654 -2751
rect 19327 -2811 19387 -2751
rect 22122 -2811 22182 -2751
rect 16150 -2899 16210 -2839
rect 18153 -2899 18213 -2839
rect 21514 -2899 21574 -2839
rect 16238 -2987 16298 -2927
rect 18337 -2987 18397 -2927
rect 21800 -2987 21860 -2927
rect 16794 -3075 16854 -3015
rect 17163 -3075 17223 -3015
rect 16882 -3163 16942 -3103
rect 17251 -3163 17311 -3103
rect 15974 -3251 16034 -3191
rect 17438 -3251 17498 -3191
rect 16414 -3339 16474 -3279
rect 17526 -3339 17586 -3279
rect 15183 -3427 15243 -3367
rect 18082 -3427 18142 -3367
rect 15367 -3515 15427 -3455
rect 18170 -3515 18230 -3455
rect 14042 -3603 14102 -3543
rect 18726 -3603 18786 -3543
rect 14482 -3691 14542 -3631
rect 18814 -3691 18874 -3631
rect 5386 -3903 5542 -3807
rect 8688 -3903 8844 -3807
rect 22539 -3903 22635 -3807
rect 23975 -3903 24071 -3807
rect 5570 -4447 5726 -4351
rect 8872 -4447 9028 -4351
rect 20870 -4447 21070 -4351
rect 21235 -4447 21331 -4351
rect 25275 -4447 25371 -4351
<< metal2 >>
rect 20870 2281 21070 2287
rect 21354 2221 21414 2281
rect 21442 2221 21502 2281
rect 21696 2221 21756 2281
rect 21784 2221 21844 2281
rect 22038 2221 22098 2281
rect 22126 2221 22186 2281
rect 22380 2221 22440 2281
rect 22468 2221 22528 2281
rect 10762 1513 10938 1519
rect 10417 1030 10477 1090
rect 10762 378 10938 1313
rect 11752 1513 11928 1519
rect 11407 1030 11467 1090
rect 10762 272 10938 278
rect 11752 378 11928 1313
rect 12742 1513 12918 1519
rect 12397 1030 12457 1090
rect 11752 272 11928 278
rect 12742 378 12918 1313
rect 13732 1513 13908 1519
rect 13387 1030 13447 1090
rect 12742 272 12918 278
rect 13732 378 13908 1313
rect 14722 1513 14898 1519
rect 14432 1030 14492 1090
rect 14520 1030 14580 1090
rect 13732 272 13908 278
rect 14722 378 14898 1313
rect 15712 1513 15888 1519
rect 15422 1030 15482 1090
rect 15510 1030 15570 1090
rect 14722 272 14898 278
rect 15712 378 15888 1313
rect 16702 1513 16878 1519
rect 16412 1030 16472 1090
rect 16500 1030 16560 1090
rect 15712 272 15888 278
rect 16702 378 16878 1313
rect 17692 1513 17868 1519
rect 17402 1030 17462 1090
rect 17490 1030 17550 1090
rect 16702 272 16878 278
rect 17692 378 17868 1313
rect 18682 1513 18858 1519
rect 18392 1030 18452 1090
rect 18480 1030 18540 1090
rect 17692 272 17868 278
rect 18682 378 18858 1313
rect 19672 1513 19848 1519
rect 19382 1030 19442 1090
rect 19470 1030 19530 1090
rect 18682 272 18858 278
rect 19672 378 19848 1313
rect 20870 1090 21070 2133
rect 22806 1379 22866 1439
rect 23148 1379 23208 1439
rect 23490 1379 23550 1439
rect 23832 1379 23892 1439
rect 24230 1379 24290 1439
rect 24572 1379 24632 1439
rect 24914 1379 24974 1439
rect 25256 1379 25316 1439
rect 20372 1030 20432 1090
rect 20460 1030 20520 1090
rect 19672 272 19848 278
rect 9056 -35 9062 25
rect 9122 -35 9508 25
rect 9568 -35 9574 25
rect 9056 -651 9062 -591
rect 9122 -651 9332 -591
rect 9392 -651 9398 -591
rect 9056 -827 9062 -767
rect 9122 -827 9420 -767
rect 9480 -827 9486 -767
rect 20690 -794 20750 -734
rect 20870 -828 21070 942
rect 9766 -1003 9772 -943
rect 9832 -1003 13447 -943
rect 9056 -1087 9062 -1027
rect 9122 -1032 9156 -1027
rect 9122 -1087 9166 -1032
rect 9156 -1088 9166 -1087
rect 9222 -1088 9232 -1032
rect 9678 -1091 9684 -1031
rect 9744 -1091 13263 -1031
rect 9056 -1175 9062 -1115
rect 9122 -1175 9128 -1115
rect 9068 -1219 9128 -1175
rect 9590 -1179 9596 -1119
rect 9656 -1179 12457 -1119
rect 9068 -1275 9166 -1219
rect 9222 -1275 9232 -1219
rect 9502 -1267 9508 -1207
rect 9568 -1267 12273 -1207
rect 9326 -1355 9332 -1295
rect 9392 -1355 11467 -1295
rect 9414 -1443 9420 -1383
rect 9480 -1443 11283 -1383
rect 9150 -1531 9156 -1471
rect 9216 -1531 10477 -1471
rect 9056 -1658 9062 -1598
rect 9122 -1602 9128 -1598
rect 9165 -1658 9175 -1602
rect 9238 -1619 9244 -1559
rect 9304 -1619 10293 -1559
rect 10233 -1647 10293 -1619
rect 9056 -1663 9128 -1658
rect 10417 -1665 10477 -1531
rect 11223 -1647 11283 -1443
rect 11407 -1647 11467 -1355
rect 12213 -1648 12273 -1267
rect 12397 -1647 12457 -1179
rect 13203 -1647 13263 -1091
rect 13387 -1647 13447 -1003
rect 5386 -3807 5542 -1843
rect 5386 -3909 5542 -3903
rect 5570 -4351 5726 -1843
rect 5754 -2575 5818 -1843
rect 5846 -2399 5910 -1843
rect 5938 -2223 6002 -1843
rect 6030 -2047 6094 -1843
rect 6030 -2113 6094 -2107
rect 5938 -2289 6002 -2283
rect 5846 -2465 5910 -2459
rect 8320 -2487 8384 -1843
rect 8412 -2311 8476 -1843
rect 8504 -2135 8568 -1843
rect 8596 -1959 8660 -1843
rect 8596 -2025 8660 -2019
rect 8504 -2201 8568 -2195
rect 8412 -2377 8476 -2371
rect 8320 -2553 8384 -2547
rect 5754 -2641 5818 -2635
rect 8688 -3807 8844 -1731
rect 9056 -1751 9062 -1691
rect 9122 -1728 9128 -1691
rect 9056 -1784 9108 -1751
rect 9164 -1784 9174 -1728
rect 14042 -1843 14193 -1783
rect 14437 -1843 14542 -1783
rect 8688 -3909 8844 -3903
rect 5570 -4453 5726 -4447
rect 8872 -4351 9028 -1843
rect 12930 -1959 12990 -1953
rect 12930 -3807 12990 -2019
rect 13018 -2047 13078 -2041
rect 13018 -3807 13078 -2107
rect 13574 -2135 13634 -2129
rect 13574 -3807 13634 -2195
rect 13662 -2223 13722 -2217
rect 13662 -3807 13722 -2283
rect 14042 -3543 14102 -1843
rect 14042 -3609 14102 -3603
rect 14218 -2311 14278 -2305
rect 14218 -3807 14278 -2371
rect 14306 -2399 14366 -2393
rect 14306 -3807 14366 -2459
rect 14482 -3631 14542 -1843
rect 14482 -3697 14542 -3691
rect 14862 -2487 14922 -2481
rect 14862 -3807 14922 -2547
rect 14950 -2575 15010 -2569
rect 14950 -3807 15010 -2635
rect 15183 -3367 15243 -1695
rect 15183 -3433 15243 -3427
rect 15367 -3455 15427 -1695
rect 15974 -1843 16209 -1783
rect 15367 -3521 15427 -3515
rect 15506 -2663 15566 -2657
rect 15506 -3807 15566 -2723
rect 15594 -2751 15654 -2745
rect 15594 -3807 15654 -2811
rect 15974 -3191 16034 -1843
rect 15974 -3257 16034 -3251
rect 16150 -2839 16210 -2833
rect 16150 -3807 16210 -2899
rect 16238 -2927 16298 -2921
rect 16238 -3807 16298 -2987
rect 16414 -3279 16474 -1783
rect 17251 -1843 17371 -1783
rect 16414 -3345 16474 -3339
rect 16794 -3015 16854 -3009
rect 16794 -3807 16854 -3075
rect 17163 -3015 17223 -1843
rect 17163 -3081 17223 -3075
rect 16882 -3103 16942 -3097
rect 16882 -3807 16942 -3163
rect 17251 -3103 17311 -1843
rect 18153 -2839 18213 -1843
rect 18153 -2905 18213 -2899
rect 18337 -2927 18397 -1843
rect 19143 -2663 19203 -1843
rect 19143 -2729 19203 -2723
rect 19327 -2751 19387 -1843
rect 20133 -2487 20193 -1843
rect 20133 -2553 20193 -2547
rect 20317 -2575 20377 -1843
rect 20317 -2641 20377 -2635
rect 19327 -2817 19387 -2811
rect 18337 -2993 18397 -2987
rect 17251 -3169 17311 -3163
rect 17438 -3191 17498 -3185
rect 17438 -3807 17498 -3251
rect 17526 -3279 17586 -3273
rect 17526 -3807 17586 -3339
rect 18082 -3367 18142 -3361
rect 18082 -3807 18142 -3427
rect 18170 -3455 18230 -3449
rect 18170 -3807 18230 -3515
rect 18726 -3543 18786 -3537
rect 18726 -3807 18786 -3603
rect 18814 -3631 18874 -3625
rect 18814 -3807 18874 -3691
rect 8872 -4453 9028 -4447
rect 20870 -4351 21070 -888
rect 24336 -1093 24392 -1083
rect 24392 -1149 24396 -1145
rect 20870 -4453 21070 -4447
rect 21235 -1203 21331 -1197
rect 21235 -4351 21331 -1299
rect 24336 -1343 24396 -1149
rect 25275 -1203 25371 -1197
rect 24970 -1214 25026 -1209
rect 24970 -1219 25030 -1214
rect 25026 -1275 25030 -1219
rect 24336 -1393 24510 -1343
rect 24450 -1529 24510 -1393
rect 24970 -1458 25030 -1275
rect 24362 -1602 24418 -1592
rect 24362 -1668 24418 -1658
rect 24648 -1728 24704 -1718
rect 22539 -1747 22635 -1741
rect 23975 -1747 24071 -1741
rect 24648 -1794 24704 -1784
rect 21514 -2839 21574 -1843
rect 21602 -2663 21662 -1843
rect 21602 -2729 21662 -2723
rect 21514 -2905 21574 -2899
rect 21800 -2927 21860 -1843
rect 22122 -2751 22182 -1843
rect 22122 -2817 22182 -2811
rect 21800 -2993 21860 -2987
rect 22539 -3807 22635 -1843
rect 22938 -2487 22998 -1843
rect 23026 -2311 23086 -1843
rect 23026 -2377 23086 -2371
rect 22938 -2553 22998 -2547
rect 23224 -2575 23284 -1843
rect 23546 -2399 23606 -1843
rect 23546 -2465 23606 -2459
rect 23224 -2641 23284 -2635
rect 22539 -3909 22635 -3903
rect 23975 -3807 24071 -1843
rect 23975 -3909 24071 -3903
rect 21235 -4453 21331 -4447
rect 25275 -4351 25371 -1299
rect 25275 -4453 25371 -4447
<< via2 >>
rect 9166 -1088 9222 -1032
rect 9166 -1275 9222 -1219
rect 9109 -1658 9122 -1602
rect 9122 -1658 9165 -1602
rect 9108 -1751 9122 -1728
rect 9122 -1751 9164 -1728
rect 9108 -1784 9164 -1751
rect 24336 -1149 24392 -1093
rect 24970 -1275 25026 -1219
rect 24362 -1658 24418 -1602
rect 24648 -1784 24704 -1728
<< metal3 >>
rect 9156 -1032 9232 -1027
rect 9156 -1088 9166 -1032
rect 9222 -1088 9232 -1032
rect 9156 -1094 9232 -1088
rect 24326 -1093 24402 -1088
rect 24326 -1094 24336 -1093
rect 9156 -1149 24336 -1094
rect 24392 -1149 24402 -1093
rect 9156 -1154 24402 -1149
rect 9156 -1219 25036 -1214
rect 9156 -1275 9166 -1219
rect 9222 -1274 24970 -1219
rect 9222 -1275 9232 -1274
rect 9156 -1280 9232 -1275
rect 24960 -1275 24970 -1274
rect 25026 -1275 25036 -1219
rect 24960 -1280 25036 -1275
rect 9099 -1602 9175 -1597
rect 9099 -1658 9109 -1602
rect 9165 -1603 9175 -1602
rect 24352 -1602 24428 -1597
rect 24352 -1603 24362 -1602
rect 9165 -1658 24362 -1603
rect 24418 -1658 24428 -1602
rect 9099 -1663 24428 -1658
rect 9098 -1728 24714 -1723
rect 9098 -1784 9108 -1728
rect 9164 -1783 24648 -1728
rect 9164 -1784 9174 -1783
rect 9098 -1789 9174 -1784
rect 24638 -1784 24648 -1783
rect 24704 -1784 24714 -1728
rect 24638 -1789 24714 -1784
use buffer_bus  buffer_bus_0
timestamp 1750863581
transform 1 0 11354 0 1 4262
box 1252 -8709 7768 -8069
use dcell_lv  dcell_lv_0
timestamp 1750867770
transform 1 0 5395 0 1 -747
box -9 -1096 3665 1886
use decoder_3  decoder_3_0
timestamp 1750842002
transform 1 0 19667 0 1 -1841
box 1403 -2 5807 4142
use lvsf_7bit  lvsf_7bit_0
timestamp 1750828667
transform 1 0 13803 0 1 -1683
box -49 -160 7013 2793
use seg_selector_lvsf  seg_selector_lvsf_0
timestamp 1750828667
transform 1 0 9839 0 1 -1829
box -45 -14 4047 2939
<< labels >>
flabel metal2 s 18461 -4447 18521 -4387 0 FreeSans 320 0 0 0 DIN0
port 0 nsew
flabel metal2 s 17817 -4447 17877 -4387 0 FreeSans 320 0 0 0 DIN1
port 1 nsew
flabel metal2 s 17173 -4447 17233 -4387 0 FreeSans 320 0 0 0 DIN2
port 2 nsew
flabel metal2 s 15885 -4447 15945 -4387 0 FreeSans 320 0 0 0 DIN4
port 4 nsew
flabel metal2 s 15241 -4447 15301 -4387 0 FreeSans 320 0 0 0 DIN5
port 5 nsew
flabel metal2 s 14597 -4447 14657 -4387 0 FreeSans 320 0 0 0 DIN6
port 6 nsew
flabel metal2 s 13953 -4447 14013 -4387 0 FreeSans 320 0 0 0 DIN7
port 7 nsew
flabel metal2 s 13309 -4447 13369 -4387 0 FreeSans 320 0 0 0 DIN8
port 8 nsew
flabel metal2 s 12665 -4447 12725 -4387 0 FreeSans 320 0 0 0 DIN9
port 9 nsew
flabel metal2 s 20690 34 20750 94 0 FreeSans 320 0 0 0 VBPLV
port 10 nsew
flabel metal2 s 20690 -794 20750 -734 0 FreeSans 320 0 0 0 VBNLV
port 11 nsew
flabel metal1 s 25348 1072 25408 1132 0 FreeSans 320 0 0 0 VBPDEC
port 12 nsew
flabel metal1 s 25348 -267 25408 -207 0 FreeSans 320 0 0 0 VBNDEC
port 13 nsew
flabel metal2 s 14520 1030 14580 1090 0 FreeSans 160 0 0 0 b[0]
port 14 nsew
flabel metal2 s 14432 1030 14492 1090 0 FreeSans 160 0 0 0 bb[0]
port 21 nsew
flabel metal2 s 15422 1030 15482 1090 0 FreeSans 160 0 0 0 bb[1]
port 22 nsew
flabel metal2 s 15510 1030 15570 1090 0 FreeSans 160 0 0 0 b[1]
port 15 nsew
flabel metal2 s 16500 1030 16560 1090 0 FreeSans 160 0 0 0 b[2]
port 16 nsew
flabel metal2 s 16412 1030 16472 1090 0 FreeSans 160 0 0 0 bb[2]
port 23 nsew
flabel metal2 s 17402 1030 17462 1090 0 FreeSans 160 0 0 0 bb[3]
port 24 nsew
flabel metal2 s 17490 1030 17550 1090 0 FreeSans 160 0 0 0 b[3]
port 17 nsew
flabel metal2 s 18392 1030 18452 1090 0 FreeSans 160 0 0 0 bb[4]
port 25 nsew
flabel metal2 s 18480 1030 18540 1090 0 FreeSans 160 0 0 0 b[4]
port 18 nsew
flabel metal2 s 19382 1030 19442 1090 0 FreeSans 160 0 0 0 bb[5]
port 26 nsew
flabel metal2 s 19470 1030 19530 1090 0 FreeSans 160 0 0 0 b[5]
port 19 nsew
flabel metal2 s 20372 1030 20432 1090 0 FreeSans 160 0 0 0 bb[6]
port 27 nsew
flabel metal2 s 20460 1030 20520 1090 0 FreeSans 160 0 0 0 b[6]
port 20 nsew
flabel metal2 s 10417 1030 10477 1090 0 FreeSans 320 180 0 0 SH[1]
port 44 nsew
flabel metal2 s 11407 1030 11467 1090 0 FreeSans 320 180 0 0 SH[2]
port 45 nsew
flabel metal2 s 12397 1030 12457 1090 0 FreeSans 320 180 0 0 SH[3]
port 46 nsew
flabel metal2 s 13387 1030 13447 1090 0 FreeSans 320 180 0 0 SH[4]
port 47 nsew
flabel metal1 s 5851 -3903 6076 -3743 0 FreeSans 1600 0 0 0 VDD
port 48 nsew
flabel metal1 s 10938 1313 11243 1513 0 FreeSans 1600 0 0 0 VDDH
port 49 nsew
flabel metal1 s 6512 -4551 6817 -4351 0 FreeSans 1600 0 0 0 GND
port 50 nsew
flabel metal2 s 16547 -4428 16572 -4409 0 FreeSans 320 0 0 0 DIN3
port 3 nsew
flabel metal2 s 24230 1379 24290 1439 0 FreeSans 320 180 0 0 dec0[0]
port 28 nsew
flabel metal2 s 24572 1379 24632 1439 0 FreeSans 320 180 0 0 dec0[1]
port 29 nsew
flabel metal2 s 24914 1379 24974 1439 0 FreeSans 320 180 0 0 dec0[2]
port 30 nsew
flabel metal2 s 25256 1379 25316 1439 0 FreeSans 320 180 0 0 dec0[3]
port 31 nsew
flabel metal2 s 22806 1379 22866 1439 0 FreeSans 320 0 0 0 dec1[0]
port 32 nsew
flabel metal2 s 23148 1379 23208 1439 0 FreeSans 320 0 0 0 dec1[1]
port 33 nsew
flabel metal2 s 23490 1379 23550 1439 0 FreeSans 320 0 0 0 dec1[2]
port 34 nsew
flabel metal2 s 23832 1379 23892 1439 0 FreeSans 320 0 0 0 dec1[3]
port 35 nsew
flabel metal2 s 21442 2221 21502 2281 0 FreeSans 320 90 0 0 dec2[0]
port 36 nsew
flabel metal2 s 21354 2221 21414 2281 0 FreeSans 320 270 0 0 dec2b[0]
port 40 nsew
flabel metal2 s 21696 2221 21756 2281 0 FreeSans 320 270 0 0 dec2b[1]
port 41 nsew
flabel metal2 s 21784 2221 21844 2281 0 FreeSans 320 90 0 0 dec2[1]
port 37 nsew
flabel metal2 s 22126 2221 22186 2281 0 FreeSans 320 90 0 0 dec2[2]
port 38 nsew
flabel metal2 s 22038 2221 22098 2281 0 FreeSans 320 270 0 0 dec2b[2]
port 42 nsew
flabel metal2 s 22380 2221 22440 2281 0 FreeSans 320 270 0 0 dec2b[3]
port 43 nsew
flabel metal2 s 22468 2221 22528 2281 0 FreeSans 320 90 0 0 dec2[3]
port 39 nsew
<< end >>
