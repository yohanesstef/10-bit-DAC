magic
tech sky130A
timestamp 1749714889
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 595 0 1 -1180
box -19 -24 65 296
use sky130_fd_sc_hd__nand4_1  x1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1749714889
transform 1 0 641 0 1 -1180
box -19 -24 249 296
use sky130_fd_sc_hd__nand4_1  x2
timestamp 1749714889
transform 1 0 365 0 1 -1180
box -19 -24 249 296
use sky130_fd_sc_hd__nand2_1  x3 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 871 0 1 -1180
box -19 -24 157 296
<< end >>
