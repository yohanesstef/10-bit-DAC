magic
tech sky130A
magscale 1 2
timestamp 1749057406
<< pwell >>
rect -307 -935 307 935
<< psubdiff >>
rect -271 865 -175 899
rect 175 865 271 899
rect -271 803 -237 865
rect 237 803 271 865
rect -271 -865 -237 -803
rect 237 -865 271 -803
rect -271 -899 -175 -865
rect 175 -899 271 -865
<< psubdiffcont >>
rect -175 865 175 899
rect -271 -803 -237 803
rect 237 -803 271 803
rect -175 -899 175 -865
<< xpolycontact >>
rect -141 337 141 769
rect -141 -769 141 -337
<< xpolyres >>
rect -141 -337 141 337
<< locali >>
rect -271 865 -175 899
rect 175 865 271 899
rect -271 803 -237 865
rect 237 803 271 865
rect -271 -865 -237 -803
rect 237 -865 271 -803
rect -271 -899 -175 -865
rect 175 -899 271 -865
<< viali >>
rect -125 354 125 751
rect -125 -751 125 -354
<< metal1 >>
rect -131 751 131 763
rect -131 354 -125 751
rect 125 354 131 751
rect -131 342 131 354
rect -131 -354 131 -342
rect -131 -751 -125 -354
rect 125 -751 131 -354
rect -131 -763 131 -751
<< properties >>
string FIXED_BBOX -254 -882 254 882
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 3.527 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 5.269k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
