magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -848 307 848
<< psubdiff >>
rect -271 778 -175 812
rect 175 778 271 812
rect -271 716 -237 778
rect 237 716 271 778
rect -271 -778 -237 -716
rect 237 -778 271 -716
rect -271 -812 -175 -778
rect 175 -812 271 -778
<< psubdiffcont >>
rect -175 778 175 812
rect -271 -716 -237 716
rect 237 -716 271 716
rect -175 -812 175 -778
<< xpolycontact >>
rect -141 250 141 682
rect -141 -682 141 -250
<< xpolyres >>
rect -141 -250 141 250
<< locali >>
rect -271 778 -175 812
rect 175 778 271 812
rect -271 716 -237 778
rect 237 716 271 778
rect -271 -778 -237 -716
rect 237 -778 271 -716
rect -271 -812 -175 -778
rect 175 -812 271 -778
<< viali >>
rect -125 267 125 664
rect -125 -664 125 -267
<< metal1 >>
rect -131 664 131 676
rect -131 267 -125 664
rect 125 267 131 664
rect -131 255 131 267
rect -131 -267 131 -255
rect -131 -664 -125 -267
rect 125 -664 131 -267
rect -131 -676 131 -664
<< properties >>
string FIXED_BBOX -254 -795 254 795
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 2.655 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 4.032k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
