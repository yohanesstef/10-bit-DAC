magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1099 307 1099
<< psubdiff >>
rect -271 1029 -175 1063
rect 175 1029 271 1063
rect -271 967 -237 1029
rect 237 967 271 1029
rect -271 -1029 -237 -967
rect 237 -1029 271 -967
rect -271 -1063 -175 -1029
rect 175 -1063 271 -1029
<< psubdiffcont >>
rect -175 1029 175 1063
rect -271 -967 -237 967
rect 237 -967 271 967
rect -175 -1063 175 -1029
<< xpolycontact >>
rect -141 501 141 933
rect -141 -933 141 -501
<< xpolyres >>
rect -141 -501 141 501
<< locali >>
rect -271 1029 -175 1063
rect 175 1029 271 1063
rect -271 967 -237 1029
rect 237 967 271 1029
rect -271 -1029 -237 -967
rect 237 -1029 271 -967
rect -271 -1063 -175 -1029
rect 175 -1063 271 -1029
<< viali >>
rect -125 518 125 915
rect -125 -915 125 -518
<< metal1 >>
rect -131 915 131 927
rect -131 518 -125 915
rect 125 518 131 915
rect -131 506 131 518
rect -131 -518 131 -506
rect -131 -915 -125 -518
rect 125 -915 131 -518
rect -131 -927 131 -915
<< properties >>
string FIXED_BBOX -254 -1046 254 1046
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 5.167 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 7.596k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
