magic
tech sky130A
magscale 1 2
timestamp 1749896124
<< error_s >>
rect 808 1711 814 1717
rect 862 1711 868 1717
rect 1450 1711 1456 1717
rect 1504 1711 1510 1717
rect 2312 1711 2318 1717
rect 2366 1711 2372 1717
rect 2954 1711 2960 1717
rect 3008 1711 3014 1717
rect 802 1705 808 1711
rect 868 1705 874 1711
rect 1444 1705 1450 1711
rect 1510 1705 1516 1711
rect 2306 1705 2312 1711
rect 2372 1705 2378 1711
rect 2948 1705 2954 1711
rect 3014 1705 3020 1711
rect 802 1651 808 1657
rect 868 1651 874 1657
rect 1444 1651 1450 1657
rect 1510 1651 1516 1657
rect 2306 1651 2312 1657
rect 2372 1651 2378 1657
rect 2948 1651 2954 1657
rect 3014 1651 3020 1657
rect 808 1645 814 1651
rect 862 1645 868 1651
rect 1450 1645 1456 1651
rect 1504 1645 1510 1651
rect 2312 1645 2318 1651
rect 2366 1645 2372 1651
rect 2954 1645 2960 1651
rect 3008 1645 3014 1651
rect 56 1623 62 1629
rect 110 1623 116 1629
rect 698 1623 704 1629
rect 752 1623 758 1629
rect 1560 1623 1566 1629
rect 1614 1623 1620 1629
rect 2202 1623 2208 1629
rect 2256 1623 2262 1629
rect 3064 1623 3070 1629
rect 3118 1623 3124 1629
rect 3706 1623 3712 1629
rect 3760 1623 3766 1629
rect 50 1617 56 1623
rect 116 1617 122 1623
rect 692 1617 698 1623
rect 758 1617 764 1623
rect 1554 1617 1560 1623
rect 1620 1617 1626 1623
rect 2196 1617 2202 1623
rect 2262 1617 2268 1623
rect 3058 1617 3064 1623
rect 3124 1617 3130 1623
rect 3700 1617 3706 1623
rect 3766 1617 3772 1623
rect 50 1563 56 1569
rect 116 1563 122 1569
rect 692 1563 698 1569
rect 758 1563 764 1569
rect 1554 1563 1560 1569
rect 1620 1563 1626 1569
rect 2196 1563 2202 1569
rect 2262 1563 2268 1569
rect 3058 1563 3064 1569
rect 3124 1563 3130 1569
rect 3700 1563 3706 1569
rect 3766 1563 3772 1569
rect 56 1557 62 1563
rect 110 1557 116 1563
rect 698 1557 704 1563
rect 752 1557 758 1563
rect 1560 1557 1566 1563
rect 1614 1557 1620 1563
rect 2202 1557 2208 1563
rect 2256 1557 2262 1563
rect 3064 1557 3070 1563
rect 3118 1557 3124 1563
rect 3706 1557 3712 1563
rect 3760 1557 3766 1563
rect 1129 1447 1135 1453
rect 1183 1447 1189 1453
rect 2633 1447 2639 1453
rect 2687 1447 2693 1453
rect 1123 1441 1129 1447
rect 1189 1441 1195 1447
rect 2627 1441 2633 1447
rect 2693 1441 2699 1447
rect 1123 1387 1129 1393
rect 1189 1387 1195 1393
rect 2627 1387 2633 1393
rect 2693 1387 2699 1393
rect 1129 1381 1135 1387
rect 1183 1381 1189 1387
rect 2633 1381 2639 1387
rect 2687 1381 2693 1387
rect 377 1359 383 1365
rect 431 1359 437 1365
rect 1881 1359 1887 1365
rect 1935 1359 1941 1365
rect 3385 1359 3391 1365
rect 3439 1359 3445 1365
rect 371 1353 377 1359
rect 437 1353 443 1359
rect 1875 1353 1881 1359
rect 1941 1353 1947 1359
rect 3379 1353 3385 1359
rect 3445 1353 3451 1359
rect 371 1299 377 1305
rect 437 1299 443 1305
rect 1875 1299 1881 1305
rect 1941 1299 1947 1305
rect 3379 1299 3385 1305
rect 3445 1299 3451 1305
rect 377 1293 383 1299
rect 431 1293 437 1299
rect 1881 1293 1887 1299
rect 1935 1293 1941 1299
rect 3385 1293 3391 1299
rect 3439 1293 3445 1299
rect 237 1271 243 1277
rect 291 1271 297 1277
rect 231 1265 237 1271
rect 297 1265 303 1271
rect 231 1211 237 1217
rect 297 1211 303 1217
rect 237 1205 243 1211
rect 291 1205 297 1211
rect 60 1095 66 1101
rect 114 1095 120 1101
rect 54 1089 60 1095
rect 120 1089 126 1095
rect 54 1035 60 1041
rect 120 1035 126 1041
rect 60 1029 66 1035
rect 114 1029 120 1035
rect 436 919 442 925
rect 490 919 496 925
rect 1070 919 1076 925
rect 1124 919 1130 925
rect 430 913 436 919
rect 496 913 502 919
rect 1064 913 1070 919
rect 1130 913 1136 919
rect 430 859 436 865
rect 496 859 502 865
rect 1064 859 1070 865
rect 1130 859 1136 865
rect 436 853 442 859
rect 490 853 496 859
rect 1070 853 1076 859
rect 1124 853 1130 859
rect 2692 831 2698 837
rect 2746 831 2752 837
rect 3326 831 3332 837
rect 3380 831 3386 837
rect 2686 825 2692 831
rect 2752 825 2758 831
rect 3320 825 3326 831
rect 3386 825 3392 831
rect 2686 771 2692 777
rect 2752 771 2758 777
rect 3320 771 3326 777
rect 3386 771 3392 777
rect 2692 765 2698 771
rect 2746 765 2752 771
rect 3326 765 3332 771
rect 3380 765 3386 771
rect 753 743 759 749
rect 807 743 813 749
rect 747 737 753 743
rect 813 737 819 743
rect 747 683 753 689
rect 813 683 819 689
rect 753 677 759 683
rect 807 677 813 683
rect 3009 655 3015 661
rect 3063 655 3069 661
rect 3003 649 3009 655
rect 3069 649 3075 655
rect 3003 595 3009 601
rect 3069 595 3075 601
rect 3009 589 3015 595
rect 3063 589 3069 595
rect 1505 567 1511 573
rect 1559 567 1565 573
rect 1499 561 1505 567
rect 1565 561 1571 567
rect 1499 507 1505 513
rect 1565 507 1571 513
rect 1505 501 1511 507
rect 1559 501 1565 507
rect 2257 479 2263 485
rect 2311 479 2317 485
rect 3702 479 3708 485
rect 3756 479 3762 485
rect 2251 473 2257 479
rect 2317 473 2323 479
rect 3696 473 3702 479
rect 3762 473 3768 479
rect 2251 419 2257 425
rect 2317 419 2323 425
rect 3696 419 3702 425
rect 3762 419 3768 425
rect 2257 413 2263 419
rect 2311 413 2317 419
rect 3702 413 3708 419
rect 3756 413 3762 419
rect 1936 303 1942 309
rect 1990 303 1996 309
rect 2578 303 2584 309
rect 2632 303 2638 309
rect 3440 303 3446 309
rect 3494 303 3500 309
rect 1930 297 1936 303
rect 1996 297 2002 303
rect 2572 297 2578 303
rect 2638 297 2644 303
rect 3434 297 3440 303
rect 3500 297 3506 303
rect 1930 243 1936 249
rect 1996 243 2002 249
rect 2572 243 2578 249
rect 2638 243 2644 249
rect 3434 243 3440 249
rect 3500 243 3506 249
rect 1936 237 1942 243
rect 1990 237 1996 243
rect 2578 237 2584 243
rect 2632 237 2638 243
rect 3440 237 3446 243
rect 3494 237 3500 243
rect 1184 215 1190 221
rect 1238 215 1244 221
rect 1826 215 1832 221
rect 1880 215 1886 221
rect 1178 209 1184 215
rect 1244 209 1250 215
rect 1820 209 1826 215
rect 1886 209 1892 215
rect 1178 155 1184 161
rect 1244 155 1250 161
rect 1820 155 1826 161
rect 1886 155 1892 161
rect 1184 149 1190 155
rect 1238 149 1244 155
rect 1826 149 1832 155
rect 1880 149 1886 155
<< metal1 >>
rect 802 1651 808 1711
rect 868 1651 874 1711
rect 1444 1651 1450 1711
rect 1510 1651 1516 1711
rect 2306 1651 2312 1711
rect 2372 1651 2378 1711
rect 2948 1651 2954 1711
rect 3014 1651 3020 1711
rect 50 1563 56 1623
rect 116 1563 122 1623
rect 692 1563 698 1623
rect 758 1563 764 1623
rect 56 1130 116 1563
rect 237 1271 297 1277
rect 54 1035 60 1095
rect 120 1035 126 1095
rect 60 460 120 1035
rect 237 736 297 1211
rect 698 1130 758 1563
rect 808 1130 868 1651
rect 1450 1130 1510 1651
rect 1554 1563 1560 1623
rect 1620 1563 1626 1623
rect 2196 1563 2202 1623
rect 2262 1563 2268 1623
rect 1560 1130 1620 1563
rect 2202 1130 2262 1563
rect 2312 1130 2372 1651
rect 2954 1130 3014 1651
rect 3058 1563 3064 1623
rect 3124 1563 3130 1623
rect 3700 1563 3706 1623
rect 3766 1563 3772 1623
rect 3064 1130 3124 1563
rect 3706 1130 3766 1563
rect 430 859 436 919
rect 496 859 502 919
rect 1064 859 1070 919
rect 1130 859 1136 919
rect 237 676 325 736
rect 436 460 496 859
rect 701 730 753 743
rect 813 730 865 743
rect 1070 460 1130 859
rect 2686 771 2692 831
rect 2752 771 2758 831
rect 3320 771 3326 831
rect 3386 771 3392 831
rect 1184 215 1244 736
rect 1826 215 1886 736
rect 1936 303 1996 736
rect 2205 419 2257 479
rect 2317 419 2369 479
rect 2578 303 2638 736
rect 2692 460 2752 771
rect 3326 460 3386 771
rect 3440 303 3500 736
rect 3696 419 3702 479
rect 3762 419 3768 479
rect 1930 243 1936 303
rect 1996 243 2002 303
rect 2572 243 2578 303
rect 2638 243 2644 303
rect 3434 243 3440 303
rect 3500 243 3506 303
rect 1178 155 1184 215
rect 1244 155 1250 215
rect 1820 155 1826 215
rect 1886 155 1892 215
<< via1 >>
rect 808 1651 868 1711
rect 1450 1651 1510 1711
rect 2312 1651 2372 1711
rect 2954 1651 3014 1711
rect 56 1563 116 1623
rect 698 1563 758 1623
rect 377 1299 437 1359
rect 237 1211 297 1271
rect 60 1035 120 1095
rect 1129 1387 1189 1447
rect 1560 1563 1620 1623
rect 2202 1563 2262 1623
rect 1881 1299 1941 1359
rect 2633 1387 2693 1447
rect 3064 1563 3124 1623
rect 3706 1563 3766 1623
rect 3385 1299 3445 1359
rect 436 859 496 919
rect 1070 859 1130 919
rect 753 683 813 743
rect 2692 771 2752 831
rect 3326 771 3386 831
rect 1505 507 1565 567
rect 2257 419 2317 479
rect 3009 595 3069 655
rect 3702 419 3762 479
rect 1936 243 1996 303
rect 2578 243 2638 303
rect 3440 243 3500 303
rect 1184 155 1244 215
rect 1826 155 1886 215
use cm_pcell2_cell  cm_pcell2_cell_0
timestamp 1749896124
transform 1 0 -3459 0 1 -1741
box 3424 1732 8172 3616
<< end >>
