magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1053 307 1053
<< psubdiff >>
rect -271 983 -175 1017
rect 175 983 271 1017
rect -271 921 -237 983
rect 237 921 271 983
rect -271 -983 -237 -921
rect 237 -983 271 -921
rect -271 -1017 -175 -983
rect 175 -1017 271 -983
<< psubdiffcont >>
rect -175 983 175 1017
rect -271 -921 -237 921
rect 237 -921 271 921
rect -175 -1017 175 -983
<< xpolycontact >>
rect -141 455 141 887
rect -141 -887 141 -455
<< xpolyres >>
rect -141 -455 141 455
<< locali >>
rect -271 983 -175 1017
rect 175 983 271 1017
rect -271 921 -237 983
rect 237 921 271 983
rect -271 -983 -237 -921
rect 237 -983 271 -921
rect -271 -1017 -175 -983
rect 175 -1017 271 -983
<< viali >>
rect -125 472 125 869
rect -125 -869 125 -472
<< metal1 >>
rect -131 869 131 881
rect -131 472 -125 869
rect 125 472 131 869
rect -131 460 131 472
rect -131 -472 131 -460
rect -131 -869 -125 -472
rect 125 -869 131 -472
rect -131 -881 131 -869
<< properties >>
string FIXED_BBOX -254 -1000 254 1000
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 4.705 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 6.94k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
