magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -684 307 684
<< psubdiff >>
rect -271 614 -175 648
rect 175 614 271 648
rect -271 552 -237 614
rect 237 552 271 614
rect -271 -614 -237 -552
rect 237 -614 271 -552
rect -271 -648 -175 -614
rect 175 -648 271 -614
<< psubdiffcont >>
rect -175 614 175 648
rect -271 -552 -237 552
rect 237 -552 271 552
rect -175 -648 175 -614
<< xpolycontact >>
rect -141 86 141 518
rect -141 -518 141 -86
<< xpolyres >>
rect -141 -86 141 86
<< locali >>
rect -271 614 -175 648
rect 175 614 271 648
rect -271 552 -237 614
rect 237 552 271 614
rect -271 -614 -237 -552
rect 237 -614 271 -552
rect -271 -648 -175 -614
rect 175 -648 271 -614
<< viali >>
rect -125 103 125 500
rect -125 -500 125 -103
<< metal1 >>
rect -131 500 131 512
rect -131 103 -125 500
rect 125 103 131 500
rect -131 91 131 103
rect -131 -103 131 -91
rect -131 -500 -125 -103
rect 125 -500 131 -103
rect -131 -512 131 -500
<< properties >>
string FIXED_BBOX -254 -631 254 631
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.015 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 1.706k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
