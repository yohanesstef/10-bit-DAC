magic
tech sky130A
magscale 1 2
timestamp 1749842112
<< nwell >>
rect -358 -762 358 762
<< mvpmos >>
rect -100 -536 100 464
<< mvpdiff >>
rect -158 452 -100 464
rect -158 -524 -146 452
rect -112 -524 -100 452
rect -158 -536 -100 -524
rect 100 452 158 464
rect 100 -524 112 452
rect 146 -524 158 452
rect 100 -536 158 -524
<< mvpdiffc >>
rect -146 -524 -112 452
rect 112 -524 146 452
<< mvnsubdiff >>
rect -292 684 292 696
rect -292 650 -184 684
rect 184 650 292 684
rect -292 638 292 650
rect -292 588 -234 638
rect -292 -588 -280 588
rect -246 -588 -234 588
rect 234 588 292 638
rect -292 -638 -234 -588
rect 234 -588 246 588
rect 280 -588 292 588
rect 234 -638 292 -588
rect -292 -650 292 -638
rect -292 -684 -184 -650
rect 184 -684 292 -650
rect -292 -696 292 -684
<< mvnsubdiffcont >>
rect -184 650 184 684
rect -280 -588 -246 588
rect 246 -588 280 588
rect -184 -684 184 -650
<< poly >>
rect -100 545 100 561
rect -100 511 -84 545
rect 84 511 100 545
rect -100 464 100 511
rect -100 -562 100 -536
<< polycont >>
rect -84 511 84 545
<< locali >>
rect -280 650 -184 684
rect 184 650 280 684
rect -280 588 -246 650
rect 246 588 280 650
rect -100 511 -84 545
rect 84 511 100 545
rect -146 452 -112 468
rect -146 -540 -112 -524
rect 112 452 146 468
rect 112 -540 146 -524
rect -280 -650 -246 -588
rect 246 -650 280 -588
rect -280 -684 -184 -650
rect 184 -684 280 -650
<< viali >>
rect -63 511 63 545
rect -146 -402 -112 330
rect 112 -402 146 330
<< metal1 >>
rect -75 545 75 551
rect -75 511 -63 545
rect 63 511 75 545
rect -75 505 75 511
rect -152 330 -106 342
rect -152 -402 -146 330
rect -112 -402 -106 330
rect -152 -414 -106 -402
rect 106 330 152 342
rect 106 -402 112 330
rect 146 -402 152 330
rect 106 -414 152 -402
<< properties >>
string FIXED_BBOX -263 -667 263 667
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 75 viadrn 75 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
