magic
tech sky130A
magscale 1 2
timestamp 1749624948
<< error_p >>
rect -313 -198 -283 130
rect -247 -132 -217 64
rect 217 -132 247 64
rect -247 -136 247 -132
rect 283 -198 313 130
rect -313 -202 313 -198
<< nwell >>
rect -283 -198 283 164
<< mvpmos >>
rect -189 -136 -29 64
rect 29 -136 189 64
<< mvpdiff >>
rect -247 52 -189 64
rect -247 -124 -235 52
rect -201 -124 -189 52
rect -247 -136 -189 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 189 52 247 64
rect 189 -124 201 52
rect 235 -124 247 52
rect 189 -136 247 -124
<< mvpdiffc >>
rect -235 -124 -201 52
rect -17 -124 17 52
rect 201 -124 235 52
<< poly >>
rect -189 145 -29 161
rect -189 111 -173 145
rect -45 111 -29 145
rect -189 64 -29 111
rect 29 145 189 161
rect 29 111 45 145
rect 173 111 189 145
rect 29 64 189 111
rect -189 -162 -29 -136
rect 29 -162 189 -136
<< polycont >>
rect -173 111 -45 145
rect 45 111 173 145
<< locali >>
rect -189 111 -173 145
rect -45 111 -29 145
rect 29 111 45 145
rect 173 111 189 145
rect -235 52 -201 68
rect -235 -140 -201 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 201 52 235 68
rect 201 -140 235 -124
<< viali >>
rect -173 111 -45 145
rect 45 111 173 145
rect -235 -124 -201 52
rect -17 -124 17 52
rect 201 -124 235 52
<< metal1 >>
rect -185 145 -33 151
rect -185 111 -173 145
rect -45 111 -33 145
rect -185 105 -33 111
rect 33 145 185 151
rect 33 111 45 145
rect 173 111 185 145
rect 33 105 185 111
rect -241 52 -195 64
rect -241 -124 -235 52
rect -201 -124 -195 52
rect -241 -136 -195 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 195 52 241 64
rect 195 -124 201 52
rect 235 -124 241 52
rect 195 -136 241 -124
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.8 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
