magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1504 307 1504
<< psubdiff >>
rect -271 1434 -175 1468
rect 175 1434 271 1468
rect -271 1372 -237 1434
rect 237 1372 271 1434
rect -271 -1434 -237 -1372
rect 237 -1434 271 -1372
rect -271 -1468 -175 -1434
rect 175 -1468 271 -1434
<< psubdiffcont >>
rect -175 1434 175 1468
rect -271 -1372 -237 1372
rect 237 -1372 271 1372
rect -175 -1468 175 -1434
<< xpolycontact >>
rect -141 906 141 1338
rect -141 -1338 141 -906
<< xpolyres >>
rect -141 -906 141 906
<< locali >>
rect -271 1434 -175 1468
rect 175 1434 271 1468
rect -271 1372 -237 1434
rect 237 1372 271 1434
rect -271 -1434 -237 -1372
rect 237 -1434 271 -1372
rect -271 -1468 -175 -1434
rect 175 -1468 271 -1434
<< viali >>
rect -125 923 125 1320
rect -125 -1320 125 -923
<< metal1 >>
rect -131 1320 131 1332
rect -131 923 -125 1320
rect 125 923 131 1320
rect -131 911 131 923
rect -131 -923 131 -911
rect -131 -1320 -125 -923
rect 125 -1320 131 -923
rect -131 -1332 131 -1320
<< properties >>
string FIXED_BBOX -254 -1451 254 1451
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 9.216 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 13.339k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
