magic
tech sky130A
magscale 1 2
timestamp 1749147130
<< pwell >>
rect -307 -745 307 745
<< psubdiff >>
rect -271 675 -175 709
rect 175 675 271 709
rect -271 613 -237 675
rect 237 613 271 675
rect -271 -675 -237 -613
rect 237 -675 271 -613
rect -271 -709 -175 -675
rect 175 -709 271 -675
<< psubdiffcont >>
rect -175 675 175 709
rect -271 -613 -237 613
rect 237 -613 271 613
rect -175 -709 175 -675
<< xpolycontact >>
rect -141 147 141 579
rect -141 -579 141 -147
<< xpolyres >>
rect -141 -147 141 147
<< locali >>
rect -271 675 -175 709
rect 175 675 271 709
rect -271 613 -237 675
rect 237 613 271 675
rect -271 -675 -237 -613
rect 237 -675 271 -613
rect -271 -709 -175 -675
rect 175 -709 271 -675
<< viali >>
rect -125 164 125 561
rect -125 -561 125 -164
<< metal1 >>
rect -131 561 131 573
rect -131 164 -125 561
rect 125 164 131 561
rect -131 152 131 164
rect -131 -164 131 -152
rect -131 -561 -125 -164
rect 125 -561 131 -164
rect -131 -573 131 -561
<< properties >>
string FIXED_BBOX -254 -692 254 692
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.63 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 2.579k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
