magic
tech sky130A
magscale 1 2
timestamp 1749479990
<< error_s >>
rect 474 344 477 362
rect 502 328 505 334
<< locali >>
rect -185 26 2061 116
<< metal1 >>
rect -793 325 -764 522
rect -511 473 -483 514
rect 161 473 189 507
rect -534 424 198 473
rect 449 468 477 527
rect 1138 468 1166 500
rect 1421 471 1449 487
rect 2126 471 2154 530
rect -511 331 -483 424
rect 161 324 189 424
rect 449 419 1192 468
rect 1421 422 2155 471
rect 449 344 477 419
rect 1138 317 1166 419
rect 1421 304 1449 422
rect 2126 347 2154 422
rect 2411 361 2439 544
rect -623 -149 -595 79
rect -339 -59 -311 112
rect -359 -111 -353 -59
rect -301 -111 -295 -59
rect -636 -201 -630 -149
rect -578 -201 -572 -149
rect -623 -237 -595 -201
rect -339 -204 -311 -111
rect 333 -149 361 104
rect 615 -56 643 122
rect 597 -108 603 -56
rect 655 -108 661 -56
rect 312 -201 318 -149
rect 370 -201 376 -149
rect 615 -194 643 -108
rect 1306 -148 1334 117
rect 1590 -55 1618 109
rect 1574 -107 1580 -55
rect 1632 -107 1638 -55
rect 1289 -200 1295 -148
rect 1347 -200 1353 -148
rect 333 -212 361 -201
rect 1590 -207 1618 -107
rect 2298 -148 2326 147
rect 2580 -51 2608 147
rect 2562 -103 2568 -51
rect 2620 -103 2626 -51
rect 2280 -200 2286 -148
rect 2338 -200 2344 -148
rect 2580 -169 2608 -103
<< via1 >>
rect -353 -111 -301 -59
rect -630 -201 -578 -149
rect 603 -108 655 -56
rect 318 -201 370 -149
rect 1580 -107 1632 -55
rect 1295 -200 1347 -148
rect 2568 -103 2620 -51
rect 2286 -200 2338 -148
<< metal2 >>
rect -359 -62 -353 -59
rect -717 -109 -353 -62
rect -359 -111 -353 -109
rect -301 -62 -295 -59
rect 597 -62 603 -56
rect -301 -108 603 -62
rect 655 -62 661 -56
rect 1574 -62 1580 -55
rect 655 -107 1580 -62
rect 1632 -62 1638 -55
rect 2562 -59 2568 -51
rect 1717 -62 2568 -59
rect 1632 -103 2568 -62
rect 2620 -59 2626 -51
rect 2620 -103 4178 -59
rect 1632 -106 4178 -103
rect 1632 -107 1744 -106
rect 655 -108 1744 -107
rect -301 -109 1744 -108
rect -301 -111 -295 -109
rect 1289 -149 1295 -148
rect -718 -196 -630 -149
rect -636 -201 -630 -196
rect -578 -196 318 -149
rect -578 -201 -572 -196
rect 312 -201 318 -196
rect 370 -196 1295 -149
rect 370 -201 376 -196
rect 1289 -200 1295 -196
rect 1347 -149 1353 -148
rect 1347 -152 1743 -149
rect 2280 -152 2286 -148
rect 1347 -196 2286 -152
rect 1347 -200 1353 -196
rect 1695 -199 2286 -196
rect 2280 -200 2286 -199
rect 2338 -152 2344 -148
rect 2338 -199 4156 -152
rect 2338 -200 2344 -199
use nswitch_2  nswitch_2_0
timestamp 1749479165
transform 1 0 144 0 1 150
box -150 -174 682 364
use nswitch_2  nswitch_2_1
timestamp 1749479165
transform 1 0 1120 0 1 138
box -150 -174 682 364
use nswitch_2  nswitch_2_2
timestamp 1749479165
transform 1 0 -812 0 1 150
box -150 -174 682 364
use nswitch_2  nswitch_2_3
timestamp 1749479165
transform 1 0 2112 0 1 178
box -150 -174 682 364
<< labels >>
flabel metal1 s -792 518 -792 518 4 FreeSans 320 0 0 0 vin[0]
port 0 se
flabel metal2 s -808 303 -808 303 4 FreeSans 320 0 0 0 dec[0]
port 1 se
flabel metal2 s -485 -91 -485 -91 4 FreeSans 320 0 0 0 VH
port 2 se
flabel metal2 s -449 -165 -449 -165 4 FreeSans 320 0 0 0 VL
port 3 se
flabel locali s -890 37 -890 37 4 FreeSans 320 0 0 0 VNB
port 4 se
<< end >>
