magic
tech sky130A
magscale 1 2
timestamp 1749386853
<< error_s >>
rect -133 1037 1043 1041
rect -133 825 -103 1037
rect -67 971 149 975
rect 209 971 425 975
rect 485 971 701 975
rect 761 971 977 975
rect -67 891 -37 971
rect 947 891 977 971
rect 1013 825 1043 1037
rect 695 -167 725 45
rect 761 -101 791 -21
rect 1775 -101 1805 -21
rect 761 -105 977 -101
rect 1037 -105 1253 -101
rect 1313 -105 1529 -101
rect 1589 -105 1805 -101
rect 1841 -167 1871 45
rect 695 -171 1871 -167
<< metal1 >>
rect -369 597 -309 975
rect -93 685 -33 975
rect 183 773 243 975
rect 459 773 519 975
rect 183 713 338 773
rect -93 625 250 685
rect -369 537 162 597
rect 102 -375 162 537
rect 190 -375 250 625
rect 278 -375 338 713
rect 366 713 519 773
rect 366 449 425 713
rect 366 -375 426 449
rect 454 -375 514 -21
rect 667 -105 727 157
rect 943 -105 1003 247
rect 1219 -105 1279 331
rect 1495 -105 1555 425
rect 760 -375 820 -105
rect 1036 -375 1096 -105
rect 1312 -375 1372 -105
use hpmos_4  hpmos_4_0
timestamp 1749384553
transform 1 0 317 0 1 -202
box 378 31 1554 281
use hpmos_4  hpmos_4_1
timestamp 1749384553
transform 1 0 -511 0 -1 1072
box 378 31 1554 281
<< end >>
