magic
tech sky130A
magscale 1 2
timestamp 1749289931
<< metal1 >>
rect 10045 -15802 10105 -15478
rect 10032 -16388 10105 -15802
rect 10133 -16450 10193 -15478
rect 10058 -17036 10193 -16450
rect 10221 -17098 10281 -15478
rect 10099 -17684 10281 -17098
<< end >>
