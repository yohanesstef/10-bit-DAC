* PEX produced on Tue Jun 17 16:16:41 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from top_buffer_opamp.ext - technology: sky130A

.subckt op_amp_posim P_IN[0] P_IN[1] P_IN[2] P_IN[3] P_IN[4] N_IN VOUT ROUT VDDA
+ GNDA
X0 VDDA.t252 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t22 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t3 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t39 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t4 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t13 VDDA.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t28 VOUT.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t19 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t39 VDDA.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t19 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t9 GNDA.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t23 VDDA.t251 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X6 GNDA.t83 opa_folded_cascode_0.monticelli_top_0.B.t6 VOUT.t2 GNDA.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t20 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t38 VDDA.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X8 GNDA.t77 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t22 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t31 GNDA.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X9 VDDA.t250 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t19 VDDA.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t0 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t37 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t24 VOUT.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 GNDA.t296 GNDA.t294 GNDA.t295 GNDA.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X13 a_n9736_226.t8 N_IN.t0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t15 GNDA.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t36 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t1 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X15 opa_folded_cascode_0.monticelli_top_0.A.t5 opa_folded_cascode_0.VB2.t12 opa_folded_cascode_0.monticelli_top_0.B.t5 GNDA.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X16 VDDA.t249 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t25 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t18 VDDA.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t25 VOUT.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 GNDA.t76 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t23 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t37 GNDA.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X19 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t15 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t5 a_n11789_1598.t15 GNDA.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X20 a_n9736_226.t4 P_IN[2].t0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t5 GNDA.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t12 N_IN.t1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t3 VDDA.t261 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X22 GNDA.t292 GNDA.t293 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t3 P_IN[4].t0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t5 VDDA.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X24 VDDA.t248 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t26 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t14 VDDA.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t8 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t18 GNDA.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X26 VDDA.t247 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t13 VDDA.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X27 VDDA.t246 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t12 VDDA.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X28 VDDA.t262 a_n4822_n1462.t2 a_n4822_n1462.t3 VDDA.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=0.696 ps=5.09 w=4.8 l=1
X29 GNDA.t75 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t15 GNDA.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X30 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t9 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t38 VDDA.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X31 GNDA.t291 GNDA.t289 GNDA.t290 GNDA.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X32 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t14 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t7 a_n11789_1598.t14 GNDA.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X33 GNDA.t103 opa_folded_cascode_0.monticelli_top_0.Bx.t6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t23 GNDA.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X34 VDDA.t245 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t29 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t11 VDDA.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X35 GNDA.t272 GNDA.t273 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t15 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t25 GNDA.t70 GNDA.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X37 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t21 N_IN.t2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t7 VDDA.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X38 VDDA.t244 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t30 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t19 VDDA.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X39 VDDA.t239 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t31 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t18 VDDA.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X40 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t37 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t10 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t8 VDDA.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X41 VDDA.t170 VDDA.t168 VDDA.t169 VDDA.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X42 GNDA.t288 GNDA.t287 GNDA.t288 GNDA.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0 ps=0 w=1.6 l=1
X43 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t12 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t35 VDDA.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X44 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t8 opa_folded_cascode_0.monticelli_top_0.Bx.t1 GNDA.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X45 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t35 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t26 GNDA.t74 GNDA.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X46 a_n9242_n890.t5 P_IN[1].t0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t10 GNDA.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X47 VDDA.t167 VDDA.t165 VDDA.t166 VDDA.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X48 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t13 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t34 VDDA.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X49 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t32 VDDA.t243 VDDA.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X50 a_n9242_n890.t9 N_IN.t3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t4 GNDA.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X51 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t18 P_IN[0].t0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t5 VDDA.t260 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X52 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t33 VDDA.t242 VDDA.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X53 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t30 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t27 GNDA.t73 GNDA.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X54 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t6 N_IN.t4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t20 VDDA.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X55 VDDA.t164 VDDA.t162 VDDA.t163 VDDA.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X56 VDDA.t241 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t34 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t17 VDDA.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X57 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t7 N_IN.t5 a_n9242_n890.t8 GNDA.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X58 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t35 VDDA.t240 VDDA.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X59 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t36 VDDA.t238 VDDA.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X60 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t33 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t16 VDDA.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X61 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t29 VOUT.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 GNDA.t270 GNDA.t271 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t26 VOUT.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 opa_folded_cascode_0.monticelli_top_0.B.t1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t16 GNDA.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X65 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t12 P_IN[1].t1 a_n9242_n890.t4 GNDA.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X66 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t20 opa_folded_cascode_0.monticelli_top_0.Ax.t6 VDDA.t266 VDDA.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X67 VDDA.t237 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t37 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t6 VDDA.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X68 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t32 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t17 VDDA.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X69 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t13 N_IN.t6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t3 VDDA.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X70 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t27 VOUT.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 a_n9242_n890.t7 N_IN.t7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t10 GNDA.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X72 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t26 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t23 VDDA.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X73 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t14 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t28 GNDA.t72 GNDA.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X74 opa_folded_cascode_0.monticelli_top_0.A.t2 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t14 VDDA.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X75 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t5 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t36 VDDA.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X76 GNDA.t71 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t29 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t7 GNDA.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X77 a_n9242_n890.t3 P_IN[1].t2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t18 GNDA.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X78 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t2 N_IN.t8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t16 VDDA.t265 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X79 GNDA.t69 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t30 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t30 GNDA.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X80 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t7 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t17 GNDA.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X81 GNDA.t268 GNDA.t269 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 VDDA.t236 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t38 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t5 VDDA.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X83 GNDA.t286 GNDA.t284 GNDA.t286 GNDA.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0 ps=0 w=1.6 l=1
X84 VDDA.t235 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t39 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t15 VDDA.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X85 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t30 VOUT.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t11 P_IN[1].t3 a_n9242_n890.t2 GNDA.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X87 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t3 N_IN.t9 a_n10488_226.t14 GNDA.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X88 opa_folded_cascode_0.VB1.t11 opa_folded_cascode_0.VB1.t10 a_n4822_n1462.t4 VDDA.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=0.696 ps=5.09 w=4.8 l=1
X89 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t3 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t9 VDDA.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X90 GNDA.t68 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t31 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t29 GNDA.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X91 a_n9736_226.t1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t3 GNDA.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X92 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t9 P_IN[3].t0 a_n10488_226.t15 GNDA.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X93 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t28 VOUT.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t6 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t16 GNDA.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X95 GNDA.t283 GNDA.t281 GNDA.t282 GNDA.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X96 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t6 N_IN.t10 a_n9242_n890.t6 GNDA.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X97 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t40 VDDA.t234 VDDA.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X98 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t22 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t22 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X99 GNDA.t279 GNDA.t280 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t28 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t32 GNDA.t67 GNDA.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X101 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t19 N_IN.t11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t5 VDDA.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X102 GNDA.t277 GNDA.t278 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t27 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t33 GNDA.t66 GNDA.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X104 opa_folded_cascode_0.VB2.t4 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t20 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t15 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X105 a_n4822_464.t5 opa_folded_cascode_0.VB2.t8 opa_folded_cascode_0.VB2.t9 GNDA.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.464 ps=3.78 w=1.6 l=1
X106 GNDA.t276 GNDA.t274 GNDA.t275 GNDA.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X107 GNDA.t266 GNDA.t267 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 GNDA.t65 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t34 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t26 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X109 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t31 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t21 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t7 VDDA.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X110 a_n7784_12197.t3 ROUT.t2 ROUT.t3 VDDA.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X111 a_n10488_226.t7 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t2 GNDA.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X112 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t23 opa_folded_cascode_0.monticelli_top_0.Ax.t7 VDDA.t263 VDDA.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X113 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t3 P_IN[1].t4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t14 VDDA.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X114 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t28 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t35 GNDA.t64 GNDA.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X115 GNDA.t63 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t36 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t27 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X116 VDDA.t161 VDDA.t159 VDDA.t160 VDDA.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X117 a_n11843_11539.t3 a_n11843_11539.t2 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t0 VDDA.t253 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X118 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t2 a_n11843_11539.t0 a_n11843_11539.t1 VDDA.t257 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X119 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t3 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t3 GNDA.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.087 ps=0.89 w=0.6 l=20
X120 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t5 N_IN.t12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t7 VDDA.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X121 VDDA.t233 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t41 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t9 VDDA.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X122 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t14 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t22 opa_folded_cascode_0.VB2.t0 VDDA.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X123 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t7 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t4 VDDA.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X124 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t31 VOUT.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t18 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t30 VDDA.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X126 GNDA.t264 GNDA.t265 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t13 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t25 opa_folded_cascode_0.VB2.t5 VDDA.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X128 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t15 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t14 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t19 GNDA.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X129 a_n9242_226.t9 N_IN.t13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t19 GNDA.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X130 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t11 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t26 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t15 VDDA.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X131 opa_folded_cascode_0.monticelli_top_0.Bx.t0 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t0 GNDA.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X132 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t6 N_IN.t14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t3 VDDA.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X133 GNDA.t262 GNDA.t263 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 opa_folded_cascode_0.VB1.t7 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t16 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t6 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X135 a_n9242_226.t5 P_IN[0].t1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t16 GNDA.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X136 opa_folded_cascode_0.monticelli_top_0.B.t2 opa_folded_cascode_0.VB1.t12 opa_folded_cascode_0.monticelli_top_0.A.t0 VDDA.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X137 GNDA.t261 GNDA.t259 GNDA.t260 GNDA.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X138 GNDA.t62 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t37 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t14 GNDA.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X139 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t32 VOUT.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t38 GNDA.t61 GNDA.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X141 a_n9736_226.t9 P_IN[2].t1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t8 GNDA.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X142 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t21 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t18 VDDA.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X143 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t17 a_n9242_n890.t1 GNDA.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X144 opa_folded_cascode_0.monticelli_top_0.Ax.t5 opa_folded_cascode_0.VB2.t13 opa_folded_cascode_0.monticelli_top_0.Bx.t5 GNDA.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X145 GNDA.t222 GNDA.t223 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t5 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t18 opa_folded_cascode_0.VB1.t6 GNDA.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X147 a_n9736_226.t7 N_IN.t15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t17 GNDA.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X148 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t10 P_IN[1].t5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t2 VDDA.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X149 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t8 N_IN.t16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t3 VDDA.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X150 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t6 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t6 VDDA.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X151 GNDA.t258 GNDA.t256 GNDA.t257 GNDA.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X152 VOUT.t42 opa_folded_cascode_0.monticelli_top_0.B.t7 GNDA.t299 GNDA.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X153 VDDA.t158 VDDA.t156 VDDA.t157 VDDA.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X154 GNDA.t255 GNDA.t253 GNDA.t254 GNDA.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0 ps=0 w=1.6 l=1
X155 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t7 P_IN[3].t1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t2 VDDA.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X156 GNDA.t252 GNDA.t250 GNDA.t251 GNDA.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X157 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t33 VOUT.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t11 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t19 a_n11789_1598.t13 GNDA.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X159 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t16 N_IN.t17 a_n9736_226.t6 GNDA.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X160 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t5 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t29 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t5 VDDA.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X161 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t12 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t30 opa_folded_cascode_0.VB2.t3 VDDA.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X162 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t26 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t39 GNDA.t60 GNDA.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X163 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t18 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t20 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t14 GNDA.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X164 GNDA.t249 GNDA.t247 GNDA.t248 GNDA.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X165 a_n11789_1598.t12 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t21 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t10 GNDA.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X166 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t13 P_IN[2].t2 a_n9736_226.t10 GNDA.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X167 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t18 N_IN.t18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t2 VDDA.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X168 GNDA.t115 opa_folded_cascode_0.monticelli_top_0.B.t8 VOUT.t15 GNDA.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X169 a_n10488_226.t6 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t22 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t4 GNDA.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X170 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t40 GNDA.t59 GNDA.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X171 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t41 GNDA.t58 GNDA.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X172 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t3 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t23 opa_folded_cascode_0.VB1.t5 GNDA.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X173 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t6 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t31 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t29 VDDA.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X174 GNDA.t242 GNDA.t243 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 GNDA.t240 GNDA.t241 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t2 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t0 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t1 GNDA.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.087 pd=0.89 as=0.174 ps=1.78 w=0.6 l=20
X177 GNDA.t57 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t42 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t13 GNDA.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X178 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t43 GNDA.t56 GNDA.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X179 VDDA.t232 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t42 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t8 VDDA.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X180 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t7 opa_folded_cascode_0.monticelli_top_0.Bx.t7 GNDA.t90 GNDA.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X181 a_n11789_1598.t11 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t5 GNDA.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X182 GNDA.t246 GNDA.t244 GNDA.t245 GNDA.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X183 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t43 VDDA.t231 VDDA.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X184 VDDA.t155 VDDA.t152 VDDA.t154 VDDA.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X185 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t19 opa_folded_cascode_0.monticelli_top_0.Bx.t8 GNDA.t300 GNDA.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X186 opa_folded_cascode_0.monticelli_top_0.A.t3 opa_folded_cascode_0.VB1.t13 opa_folded_cascode_0.monticelli_top_0.B.t3 VDDA.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X187 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t15 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t32 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t35 VDDA.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X188 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t20 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t33 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t23 VDDA.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X189 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t44 VDDA.t230 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X190 GNDA.t239 GNDA.t237 GNDA.t238 GNDA.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X191 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t17 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t13 GNDA.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X192 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t2 N_IN.t19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t11 VDDA.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X193 VDDA.t229 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t45 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t12 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X194 GNDA.t236 GNDA.t233 GNDA.t235 GNDA.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0 ps=0 w=1.6 l=1
X195 a_n11789_1598.t10 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t26 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t4 GNDA.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X196 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t46 VDDA.t228 VDDA.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X197 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t44 GNDA.t55 GNDA.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X198 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t7 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t27 a_n11789_1598.t9 GNDA.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X199 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t3 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t28 a_n10488_226.t5 GNDA.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X200 VDDA.t227 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t47 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t15 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X201 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t29 VOUT.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t16 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t29 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t12 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X203 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t22 P_IN[0].t2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t9 VDDA.t261 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X204 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t11 P_IN[2].t3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t11 VDDA.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X205 VDDA.t151 VDDA.t149 VDDA.t150 VDDA.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X206 opa_folded_cascode_0.VB1.t4 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t30 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t1 GNDA.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X207 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t34 VOUT.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t4 N_IN.t20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t22 VDDA.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X209 VDDA.t226 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t48 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t14 VDDA.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X210 GNDA.t220 GNDA.t221 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 GNDA.t107 opa_folded_cascode_0.monticelli_top_0.Bx.t9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t13 GNDA.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X212 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t2 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t34 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t28 VDDA.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X213 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t49 VDDA.t225 VDDA.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X214 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t30 VOUT.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 a_n4822_n1462.t5 opa_folded_cascode_0.VB1.t8 opa_folded_cascode_0.VB1.t9 VDDA.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.696 pd=5.09 as=1.392 ps=10.18 w=4.8 l=1
X216 a_n11789_1598.t8 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t31 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t6 GNDA.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X217 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t14 N_IN.t21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t1 VDDA.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X218 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t50 VDDA.t224 VDDA.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X219 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t25 opa_folded_cascode_0.monticelli_top_0.Bx.t10 GNDA.t109 GNDA.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X220 GNDA.t218 GNDA.t219 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 GNDA.t54 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t45 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t12 GNDA.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X222 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t9 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t32 a_n11789_1598.t7 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X223 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t31 VOUT.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t51 VDDA.t223 VDDA.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X225 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t8 P_IN[4].t1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t2 VDDA.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X226 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t26 opa_folded_cascode_0.monticelli_top_0.Bx.t11 GNDA.t298 GNDA.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X227 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t29 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t46 GNDA.t53 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X228 a_n10488_226.t10 P_IN[3].t2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t2 GNDA.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X229 VDDA.t222 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t52 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t3 VDDA.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X230 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t35 VOUT.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 a_n10488_226.t13 N_IN.t22 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t0 GNDA.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X232 GNDA.t232 GNDA.t230 GNDA.t231 GNDA.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X233 GNDA.t229 GNDA.t227 GNDA.t228 GNDA.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X234 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t10 N_IN.t23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t0 VDDA.t260 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X235 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t53 VDDA.t221 VDDA.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X236 GNDA.t216 GNDA.t217 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 VDDA.t220 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t54 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t8 VDDA.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X238 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t1 P_IN[4].t2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t23 VDDA.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X239 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t14 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t35 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t34 VDDA.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X240 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t47 GNDA.t52 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X241 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t36 VOUT.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t32 VOUT.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 VDDA.t219 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t55 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t7 VDDA.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X244 VDDA.t148 VDDA.t146 VDDA.t147 VDDA.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X245 a_n4822_464.t3 a_n4822_464.t2 GNDA.t95 GNDA.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.464 ps=3.78 w=1.6 l=1
X246 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t56 VDDA.t218 VDDA.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X247 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t33 VOUT.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t57 VDDA.t217 VDDA.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X249 GNDA.t303 opa_folded_cascode_0.monticelli_top_0.Bx.t12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t27 GNDA.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X250 VDDA.t216 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t58 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t6 VDDA.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X251 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t59 VDDA.t215 VDDA.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X252 VDDA.t214 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t60 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t11 VDDA.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X253 opa_folded_cascode_0.monticelli_top_0.Bx.t4 opa_folded_cascode_0.VB2.t14 opa_folded_cascode_0.monticelli_top_0.Ax.t4 GNDA.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X254 VDDA.t145 VDDA.t143 VDDA.t144 VDDA.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X255 GNDA.t226 GNDA.t224 GNDA.t225 GNDA.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X256 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t61 VDDA.t213 VDDA.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X257 VDDA.t142 VDDA.t140 VDDA.t141 VDDA.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X258 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t10 P_IN[2].t4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t24 VDDA.t265 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X259 opa_folded_cascode_0.monticelli_top_0.Ax.t3 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t36 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t21 VDDA.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X260 VDDA.t139 VDDA.t137 VDDA.t138 VDDA.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X261 GNDA.t215 GNDA.t213 GNDA.t214 GNDA.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X262 VDDA.t212 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t62 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t6 VDDA.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X263 GNDA.t142 GNDA.t143 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 VDDA.t136 VDDA.t134 VDDA.t135 VDDA.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X265 VDDA.t133 VDDA.t131 VDDA.t132 VDDA.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X266 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t24 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t37 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t19 VDDA.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X267 a_n4822_n1462.t1 a_n4822_n1462.t0 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.696 pd=5.09 as=1.392 ps=10.18 w=4.8 l=1
X268 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t48 GNDA.t51 GNDA.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X269 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t23 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t38 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t33 VDDA.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X270 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t49 GNDA.t50 GNDA.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X271 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t3 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t33 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t11 GNDA.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X272 VDDA.t211 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t63 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t5 VDDA.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X273 opa_folded_cascode_0.VB2.t2 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t39 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t11 VDDA.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X274 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t37 VOUT.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t6 P_IN[3].t3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t1 VDDA.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X276 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t64 VDDA.t210 VDDA.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X277 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t5 N_IN.t24 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t4 VDDA.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X278 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t10 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t40 opa_folded_cascode_0.VB2.t7 VDDA.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X279 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t14 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t41 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t10 VDDA.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X280 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t65 VDDA.t209 VDDA.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X281 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t34 VOUT.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 VOUT.t12 opa_folded_cascode_0.monticelli_top_0.A.t6 VDDA.t255 VDDA.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X283 GNDA.t211 GNDA.t212 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t34 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t10 GNDA.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X285 GNDA.t209 GNDA.t210 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 VDDA.t130 VDDA.t128 VDDA.t129 VDDA.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X287 GNDA.t49 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t50 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t10 GNDA.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X288 GNDA.t208 GNDA.t206 GNDA.t207 GNDA.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X289 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t27 P_IN[1].t6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t1 VDDA.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X290 ROUT.t1 ROUT.t0 a_n7784_12197.t2 VDDA.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X291 a_n9242_226.t4 P_IN[0].t3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t6 GNDA.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X292 VDDA.t127 VDDA.t125 VDDA.t126 VDDA.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X293 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t22 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t42 opa_folded_cascode_0.monticelli_top_0.Ax.t2 VDDA.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X294 a_n9242_226.t8 N_IN.t25 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t9 GNDA.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X295 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t38 VOUT.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 VDDA.t264 opa_folded_cascode_0.monticelli_top_0.A.t7 VOUT.t45 VDDA.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X297 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t0 P_IN[1].t7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t6 VDDA.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X298 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t66 VDDA.t208 VDDA.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X299 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t0 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t43 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t13 VDDA.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X300 GNDA.t204 GNDA.t205 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 GNDA.t203 GNDA.t201 GNDA.t202 GNDA.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X302 VDDA.t124 VDDA.t121 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X303 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t39 VOUT.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 GNDA.t48 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t51 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t11 GNDA.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X305 GNDA.t200 GNDA.t197 GNDA.t199 GNDA.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X306 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t67 VDDA.t207 VDDA.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X307 VDDA.t120 VDDA.t118 VDDA.t119 VDDA.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X308 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t18 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t44 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t17 VDDA.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X309 GNDA.t195 GNDA.t196 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t35 a_n9736_226.t0 GNDA.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X311 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t68 VDDA.t206 VDDA.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X312 GNDA.t193 GNDA.t194 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t6 N_IN.t26 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t4 VDDA.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X314 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t0 P_IN[3].t4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t5 VDDA.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X315 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t8 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t45 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t2 VDDA.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X316 GNDA.t192 GNDA.t190 GNDA.t191 GNDA.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X317 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t7 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t36 a_n10488_226.t4 GNDA.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X318 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t27 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t46 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t15 VDDA.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X319 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t52 GNDA.t47 GNDA.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X320 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t69 VDDA.t205 VDDA.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X321 VDDA.t117 VDDA.t115 VDDA.t116 VDDA.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X322 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t20 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t47 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t32 VDDA.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X323 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t26 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t48 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t11 VDDA.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X324 a_n11789_1598.t6 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t37 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t8 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X325 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t5 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t38 a_n10488_226.t3 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X326 GNDA.t177 GNDA.t178 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 GNDA.t97 a_n4822_464.t0 a_n4822_464.t1 GNDA.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.232 ps=1.89 w=1.6 l=1
X328 VDDA.t114 VDDA.t112 VDDA.t113 VDDA.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X329 a_n11789_1598.t5 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t39 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t3 GNDA.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X330 GNDA.t175 GNDA.t176 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 VDDA.t111 VDDA.t109 VDDA.t110 VDDA.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X332 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t40 VOUT.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 GNDA.t46 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t53 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t20 GNDA.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X334 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t27 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t49 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t17 VDDA.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X335 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t7 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t50 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t4 VDDA.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X336 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t54 GNDA.t45 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X337 GNDA.t173 GNDA.t174 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t70 VDDA.t204 VDDA.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X339 VDDA.t108 VDDA.t106 VDDA.t107 VDDA.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X340 VDDA.t105 VDDA.t103 VDDA.t104 VDDA.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X341 GNDA.t93 opa_folded_cascode_0.monticelli_top_0.Bx.t13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t2 GNDA.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X342 a_n11789_1598.t4 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t40 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t2 GNDA.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X343 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t8 P_IN[0].t4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t21 VDDA.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X344 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t12 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t41 opa_folded_cascode_0.monticelli_top_0.B.t0 GNDA.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X345 a_n9736_226.t2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t42 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t1 GNDA.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X346 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t16 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t51 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t29 VDDA.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X347 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t71 VDDA.t203 VDDA.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X348 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t55 GNDA.t44 GNDA.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X349 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t15 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t43 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t9 GNDA.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X350 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t35 VOUT.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 opa_folded_cascode_0.monticelli_top_0.Ax.t1 opa_folded_cascode_0.VB1.t14 opa_folded_cascode_0.monticelli_top_0.Bx.t3 VDDA.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X352 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t4 P_IN[0].t5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t17 VDDA.t256 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X353 GNDA.t189 GNDA.t187 GNDA.t188 GNDA.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X354 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t25 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t52 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t10 VDDA.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X355 GNDA.t185 GNDA.t186 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t6 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t44 a_n10488_226.t2 GNDA.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X357 VDDA.t102 VDDA.t99 VDDA.t101 VDDA.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X358 VDDA.t202 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t72 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t6 VDDA.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X359 opa_folded_cascode_0.VB2.t11 opa_folded_cascode_0.VB2.t10 a_n4822_464.t4 GNDA.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.232 ps=1.89 w=1.6 l=1
X360 GNDA.t184 GNDA.t182 GNDA.t183 GNDA.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X361 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t56 GNDA.t43 GNDA.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X362 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t24 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t53 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t5 VDDA.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X363 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t0 N_IN.t27 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t7 VDDA.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X364 GNDA.t42 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t57 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t23 GNDA.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X365 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t73 VDDA.t194 VDDA.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X366 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t36 VOUT.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t3 a_n11843_11539.t6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t21 VDDA.t257 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X368 GNDA.t181 GNDA.t179 GNDA.t180 GNDA.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X369 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t23 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t58 GNDA.t41 GNDA.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X370 VDDA.t98 VDDA.t96 VDDA.t97 VDDA.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X371 VDDA.t201 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t74 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t3 VDDA.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X372 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t75 VDDA.t200 VDDA.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X373 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t1 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t21 GNDA.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.087 pd=0.89 as=0.174 ps=1.78 w=0.6 l=20
X374 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t31 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t54 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t19 VDDA.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X375 GNDA.t40 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t59 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t22 GNDA.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X376 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t9 P_IN[2].t5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t9 VDDA.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X377 GNDA.t172 GNDA.t170 GNDA.t171 GNDA.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X378 GNDA.t140 GNDA.t141 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 GNDA.t39 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t60 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t21 GNDA.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X380 GNDA.t302 opa_folded_cascode_0.monticelli_top_0.Bx.t14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t25 GNDA.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X381 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t30 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t55 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t4 VDDA.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X382 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t4 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t56 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t23 VDDA.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X383 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t8 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t45 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t14 GNDA.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X384 VDDA.t95 VDDA.t93 VDDA.t94 VDDA.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X385 VDDA.t259 opa_folded_cascode_0.monticelli_top_0.Ax.t8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t20 VDDA.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X386 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t76 VDDA.t199 VDDA.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X387 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t29 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t57 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t22 VDDA.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X388 GNDA.t138 GNDA.t139 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 VDDA.t92 VDDA.t90 VDDA.t91 VDDA.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X390 VDDA.t89 VDDA.t87 VDDA.t88 VDDA.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X391 VDDA.t86 VDDA.t84 VDDA.t85 VDDA.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X392 GNDA.t33 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t61 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t3 GNDA.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X393 GNDA.t37 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t62 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t22 GNDA.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X394 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t46 a_n11789_1598.t3 GNDA.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X395 VDDA.t83 VDDA.t81 VDDA.t82 VDDA.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X396 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t22 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t58 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t9 VDDA.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X397 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t38 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t63 GNDA.t38 GNDA.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X398 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t7 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t47 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t1 GNDA.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X399 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t17 P_IN[2].t6 a_n9736_226.t11 GNDA.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X400 GNDA.t36 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t64 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t39 GNDA.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X401 a_n11843_11539.t5 ROUT.t4 a_n7784_12197.t0 VDDA.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X402 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t77 VDDA.t198 VDDA.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X403 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t41 VOUT.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 GNDA.t136 GNDA.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t78 VDDA.t197 VDDA.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X406 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t21 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t65 GNDA.t35 GNDA.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X407 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t18 N_IN.t28 a_n9736_226.t5 GNDA.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X408 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t66 GNDA.t34 GNDA.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X409 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t79 VDDA.t196 VDDA.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X410 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t42 VOUT.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VDDA.t80 VDDA.t78 VDDA.t79 VDDA.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X412 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t37 VOUT.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t28 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t59 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t21 VDDA.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X414 GNDA.t32 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t67 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t20 GNDA.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X415 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t8 a_n11843_11539.t7 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t1 VDDA.t253 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X416 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t80 VDDA.t195 VDDA.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X417 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t27 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t60 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t18 VDDA.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X418 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t38 VOUT.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 VDDA.t267 opa_folded_cascode_0.monticelli_top_0.Ax.t9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t21 VDDA.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X420 GNDA.t31 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t68 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t31 GNDA.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X421 GNDA.t30 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t69 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t8 GNDA.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X422 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t22 P_IN[4].t3 a_n11789_1598.t23 GNDA.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X423 VDDA.t193 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t81 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t0 VDDA.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X424 GNDA.t163 GNDA.t164 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t70 GNDA.t29 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X426 VDDA.t192 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t82 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t3 VDDA.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X427 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t83 VDDA.t191 VDDA.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X428 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t13 N_IN.t29 a_n11789_1598.t20 GNDA.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X429 VDDA.t190 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t84 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t3 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X430 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t43 VOUT.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 GNDA.t161 GNDA.t162 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t39 VOUT.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t85 VDDA.t189 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X434 VDDA.t77 VDDA.t75 VDDA.t76 VDDA.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X435 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t1 N_IN.t30 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t15 VDDA.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X436 VDDA.t188 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t86 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t2 VDDA.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X437 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t21 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t61 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t3 VDDA.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X438 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t40 VOUT.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t87 VDDA.t187 VDDA.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X440 VDDA.t74 VDDA.t72 VDDA.t73 VDDA.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X441 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t15 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t62 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t28 VDDA.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X442 GNDA.t28 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t71 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t8 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X443 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t26 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t63 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t17 VDDA.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X444 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t30 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t64 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t14 VDDA.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X445 VDDA.t186 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t88 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t1 VDDA.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X446 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t13 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t65 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t21 VDDA.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X447 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t26 P_IN[2].t7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t8 VDDA.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X448 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t24 opa_folded_cascode_0.monticelli_top_0.Bx.t15 GNDA.t105 GNDA.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X449 GNDA.t168 GNDA.t169 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 a_n9242_n890.t0 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t48 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t0 GNDA.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X451 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t15 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t66 opa_folded_cascode_0.monticelli_top_0.A.t1 VDDA.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X452 VDDA.t185 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t89 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t0 VDDA.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X453 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t3 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t67 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t7 VDDA.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X454 VDDA.t71 VDDA.t69 VDDA.t70 VDDA.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X455 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t90 VDDA.t184 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X456 VDDA.t183 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t91 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t7 VDDA.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X457 GNDA.t167 GNDA.t165 GNDA.t166 GNDA.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X458 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t0 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t49 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t6 GNDA.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X459 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t9 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t68 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t12 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X460 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t20 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t25 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t0 GNDA.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.087 ps=0.89 w=0.6 l=20
X461 GNDA.t160 GNDA.t158 GNDA.t159 GNDA.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X462 VDDA.t68 VDDA.t66 VDDA.t67 VDDA.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X463 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t12 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t69 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t16 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X464 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t5 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t50 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t11 GNDA.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X465 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t0 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t51 opa_folded_cascode_0.VB1.t3 GNDA.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X466 GNDA.t27 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t72 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t33 GNDA.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X467 GNDA.t157 GNDA.t154 GNDA.t156 GNDA.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X468 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t4 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t52 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t10 GNDA.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X469 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t92 VDDA.t182 VDDA.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X470 GNDA.t152 GNDA.t153 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t44 VOUT.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 a_n10488_226.t12 N_IN.t31 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t1 GNDA.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X473 VDDA.t181 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t93 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t1 VDDA.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X474 GNDA.t26 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t73 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t2 GNDA.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X475 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t94 VDDA.t180 VDDA.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X476 VDDA.t65 VDDA.t62 VDDA.t64 VDDA.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X477 a_n10488_226.t9 P_IN[3].t5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t1 GNDA.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X478 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t3 P_IN[4].t4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t0 VDDA.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X479 GNDA.t25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t74 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t19 GNDA.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X480 VDDA.t61 VDDA.t59 VDDA.t60 VDDA.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X481 GNDA.t151 GNDA.t148 GNDA.t150 GNDA.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X482 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t45 VOUT.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 GNDA.t24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t75 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t34 GNDA.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X484 VDDA.t178 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t95 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t0 VDDA.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X485 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t11 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t70 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t12 VDDA.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X486 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t46 VOUT.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t0 P_IN[3].t6 a_n10488_226.t8 GNDA.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X488 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t31 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t71 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t11 VDDA.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X489 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t3 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t53 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t13 GNDA.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X490 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t6 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t72 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t2 VDDA.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X491 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t2 N_IN.t32 a_n10488_226.t11 GNDA.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X492 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t20 opa_folded_cascode_0.monticelli_top_0.Bx.t16 GNDA.t301 GNDA.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X493 GNDA.t134 GNDA.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 opa_folded_cascode_0.monticelli_top_0.B.t4 opa_folded_cascode_0.VB2.t15 opa_folded_cascode_0.monticelli_top_0.A.t4 GNDA.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X495 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t20 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t73 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t10 VDDA.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X496 GNDA.t23 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t76 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t18 GNDA.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X497 VDDA.t58 VDDA.t55 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X498 opa_folded_cascode_0.VB1.t2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t54 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t7 GNDA.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X499 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t55 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t12 GNDA.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X500 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t19 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t74 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t9 VDDA.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X501 a_n11789_1598.t2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t56 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t0 GNDA.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X502 GNDA.t147 GNDA.t144 GNDA.t146 GNDA.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X503 GNDA.t132 GNDA.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t47 VOUT.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t57 a_n9242_226.t0 GNDA.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X506 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t1 N_IN.t33 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t9 VDDA.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X507 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t16 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t75 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t25 VDDA.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X508 opa_folded_cascode_0.VB2.t6 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t76 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t9 VDDA.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X509 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t13 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t58 a_n11789_1598.t1 GNDA.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X510 GNDA.t131 GNDA.t129 GNDA.t130 GNDA.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X511 opa_folded_cascode_0.monticelli_top_0.Bx.t2 opa_folded_cascode_0.VB1.t15 opa_folded_cascode_0.monticelli_top_0.Ax.t0 VDDA.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X512 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t96 VDDA.t177 VDDA.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X513 GNDA.t127 GNDA.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t10 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t77 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t24 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X515 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t10 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t78 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t14 VDDA.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X516 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t9 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t79 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t15 VDDA.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X517 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t23 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t80 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t7 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X518 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t59 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t5 GNDA.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X519 opa_folded_cascode_0.VB1.t1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t60 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t4 GNDA.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X520 VDDA.t54 VDDA.t51 VDDA.t53 VDDA.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X521 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t13 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t81 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t8 VDDA.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X522 VOUT.t9 opa_folded_cascode_0.monticelli_top_0.A.t8 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X523 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t5 N_IN.t34 a_n9242_226.t7 GNDA.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X524 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t17 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t77 GNDA.t22 GNDA.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X525 a_n10488_226.t1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t61 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t0 GNDA.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X526 a_n11789_1598.t21 P_IN[4].t5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t7 GNDA.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X527 opa_folded_cascode_0.VB2.t1 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t82 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t8 VDDA.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X528 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t12 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t62 a_n11789_1598.t0 GNDA.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X529 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t3 P_IN[0].t6 a_n9242_226.t3 GNDA.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X530 VDDA.t176 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t97 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t2 VDDA.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X531 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t41 VOUT.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t63 opa_folded_cascode_0.VB1.t0 GNDA.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X533 a_n11789_1598.t19 N_IN.t35 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t12 GNDA.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X534 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t0 N_IN.t36 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t17 VDDA.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X535 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t32 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t78 GNDA.t21 GNDA.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X536 VDDA.t175 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t98 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t1 VDDA.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X537 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t99 VDDA.t174 VDDA.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X538 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t14 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t83 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t20 VDDA.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X539 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t0 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t64 a_n9736_226.t3 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X540 VDDA.t173 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t100 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t0 VDDA.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X541 GNDA.t125 GNDA.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t16 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t79 GNDA.t20 GNDA.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X543 VDDA.t1 opa_folded_cascode_0.monticelli_top_0.A.t9 VOUT.t0 VDDA.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X544 a_n7784_12197.t1 ROUT.t5 a_n11843_11539.t4 VDDA.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X545 GNDA.t19 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t80 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t4 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X546 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t11 N_IN.t37 a_n11789_1598.t18 GNDA.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X547 GNDA.t123 GNDA.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t6 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t84 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t22 VDDA.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X549 GNDA.t121 GNDA.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 a_n10488_226.t0 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t65 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t1 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X551 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t4 P_IN[3].t7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t4 VDDA.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X552 VDDA.t50 VDDA.t47 VDDA.t49 VDDA.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X553 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t19 P_IN[4].t6 a_n11789_1598.t22 GNDA.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X554 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t36 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t81 GNDA.t18 GNDA.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X555 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t11 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t85 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t21 VDDA.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X556 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t8 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t86 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t25 VDDA.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X557 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t42 VOUT.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X558 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t23 P_IN[0].t7 a_n9242_226.t2 GNDA.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X559 VDDA.t46 VDDA.t43 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X560 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t0 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t66 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t4 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X561 VOUT.t16 opa_folded_cascode_0.monticelli_top_0.B.t9 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X562 a_n11789_1598.t17 N_IN.t38 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t14 GNDA.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X563 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t8 N_IN.t39 a_n9242_226.t6 GNDA.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X564 GNDA.t111 opa_folded_cascode_0.monticelli_top_0.Bx.t17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t15 GNDA.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X565 VDDA.t172 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t101 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t0 VDDA.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X566 a_n11789_1598.t16 P_IN[4].t7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t4 GNDA.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X567 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t20 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t87 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t12 VDDA.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X568 a_n9242_226.t1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t67 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t0 GNDA.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X569 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t43 VOUT.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n90 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t8 151.631
R1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t32 142.488
R2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t48 142.488
R3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n30 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t27 142.488
R4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t96 142.488
R5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n50 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t42 142.488
R6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n39 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t40 142.488
R7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n70 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t70 142.488
R8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n59 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t63 142.488
R9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t82 141.704
R10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t69 141.704
R11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t47 141.704
R12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t77 141.704
R13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t39 141.704
R14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t90 141.704
R15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t98 141.704
R16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t53 141.704
R17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t30 141.704
R18 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t71 141.704
R19 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t72 141.704
R20 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t61 141.704
R21 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t93 141.704
R22 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t67 141.704
R23 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t60 141.704
R24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t36 141.704
R25 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t86 141.704
R26 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t46 141.704
R27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n30 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t56 141.704
R28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n31 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t58 141.704
R29 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n32 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t85 141.704
R30 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n33 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t88 141.704
R31 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n34 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t59 141.704
R32 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n35 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t84 141.704
R33 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n36 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t66 141.704
R34 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t38 141.704
R35 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t65 141.704
R36 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t81 141.704
R37 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t94 141.704
R38 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t95 141.704
R39 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t64 141.704
R40 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t91 141.704
R41 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t92 141.704
R42 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t41 141.704
R43 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t68 141.704
R44 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t89 141.704
R45 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n50 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t73 141.704
R46 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n51 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t74 141.704
R47 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n52 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t23 141.704
R48 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n53 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t26 141.704
R49 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n54 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t75 141.704
R50 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n55 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t22 141.704
R51 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n56 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t83 141.704
R52 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n49 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t52 141.704
R53 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n48 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t79 141.704
R54 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n47 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t101 141.704
R55 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n46 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t35 141.704
R56 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n45 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t37 141.704
R57 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n44 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t78 141.704
R58 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n43 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t29 141.704
R59 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n42 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t33 141.704
R60 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n41 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t62 141.704
R61 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n40 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t87 141.704
R62 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n39 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t28 141.704
R63 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n70 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t97 141.704
R64 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n71 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t99 141.704
R65 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n72 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t45 141.704
R66 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n73 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t49 141.704
R67 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n74 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t100 141.704
R68 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n75 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t44 141.704
R69 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n76 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t31 141.704
R70 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n69 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t76 141.704
R71 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n68 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t25 141.704
R72 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n67 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t43 141.704
R73 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n66 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t55 141.704
R74 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n65 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t57 141.704
R75 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n64 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t24 141.704
R76 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n63 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t51 141.704
R77 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n62 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t54 141.704
R78 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n61 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t80 141.704
R79 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n60 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t34 141.704
R80 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n59 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t50 141.704
R81 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n90 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t21 134.811
R82 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n92 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t3 134.712
R83 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n94 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t4 134.712
R84 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n94 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t1 134.712
R85 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n82 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t19 134.712
R86 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n82 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t17 134.712
R87 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n80 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t13 134.712
R88 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n80 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t16 134.712
R89 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n79 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t12 134.712
R90 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n79 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t7 134.712
R91 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n99 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t14 134.712
R92 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n99 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t11 134.712
R93 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n97 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t18 134.712
R94 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n97 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t15 134.712
R95 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n88 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t6 134.712
R96 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n88 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t5 134.712
R97 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n86 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t20 134.712
R98 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n86 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t10 134.712
R99 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n85 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t2 134.712
R100 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n85 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t9 134.712
R101 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n92 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t0 134.712
R102 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n96 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n91 9.92246
R103 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n96 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n95 9.18808
R104 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n81 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n79 7.7474
R105 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n87 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n85 7.7474
R106 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n98 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n96 5.72717
R107 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n102 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n84 5.30474
R108 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n95 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n94 4.61407
R109 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n83 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n82 4.61407
R110 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n81 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n80 4.61407
R111 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n100 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n99 4.61407
R112 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n98 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n97 4.61407
R113 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n89 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n88 4.61407
R114 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n87 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n86 4.61407
R115 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n93 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n92 4.61407
R116 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n38 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n18 4.07135
R117 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n102 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n101 3.4105
R118 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n78 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n77 3.4105
R119 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n58 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n57 3.4105
R120 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n38 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n37 3.4105
R121 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n89 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n87 3.13383
R122 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n100 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n98 3.13383
R123 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n83 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n81 3.13383
R124 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n95 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n93 3.13383
R125 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n101 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n100 2.73592
R126 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n84 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n83 1.96508
R127 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n91 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n90 1.87758
R128 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n93 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n84 1.16925
R129 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n0 0.783833
R130 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n1 0.783833
R131 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n2 0.783833
R132 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n3 0.783833
R133 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n4 0.783833
R134 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n5 0.783833
R135 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n6 0.783833
R136 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n7 0.783833
R137 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n8 0.783833
R138 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n9 0.783833
R139 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n16 0.783833
R140 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n15 0.783833
R141 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n14 0.783833
R142 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n13 0.783833
R143 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n12 0.783833
R144 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n11 0.783833
R145 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n19 0.783833
R146 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n20 0.783833
R147 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n21 0.783833
R148 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n22 0.783833
R149 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n23 0.783833
R150 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n24 0.783833
R151 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n25 0.783833
R152 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n26 0.783833
R153 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n27 0.783833
R154 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n28 0.783833
R155 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n36 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n35 0.783833
R156 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n35 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n34 0.783833
R157 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n34 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n33 0.783833
R158 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n33 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n32 0.783833
R159 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n32 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n31 0.783833
R160 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n31 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n30 0.783833
R161 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n40 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n39 0.783833
R162 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n41 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n40 0.783833
R163 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n42 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n41 0.783833
R164 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n43 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n42 0.783833
R165 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n44 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n43 0.783833
R166 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n45 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n44 0.783833
R167 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n46 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n45 0.783833
R168 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n47 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n46 0.783833
R169 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n48 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n47 0.783833
R170 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n49 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n48 0.783833
R171 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n56 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n55 0.783833
R172 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n55 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n54 0.783833
R173 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n54 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n53 0.783833
R174 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n53 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n52 0.783833
R175 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n52 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n51 0.783833
R176 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n51 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n50 0.783833
R177 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n60 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n59 0.783833
R178 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n61 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n60 0.783833
R179 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n62 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n61 0.783833
R180 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n63 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n62 0.783833
R181 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n64 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n63 0.783833
R182 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n65 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n64 0.783833
R183 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n66 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n65 0.783833
R184 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n67 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n66 0.783833
R185 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n68 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n67 0.783833
R186 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n69 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n68 0.783833
R187 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n76 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n75 0.783833
R188 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n75 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n74 0.783833
R189 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n74 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n73 0.783833
R190 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n73 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n72 0.783833
R191 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n72 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n71 0.783833
R192 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n71 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n70 0.783833
R193 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n17 0.777583
R194 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n37 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n36 0.777583
R195 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n57 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n56 0.777583
R196 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n77 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n76 0.777583
R197 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n78 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n58 0.661348
R198 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n101 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n89 0.398417
R199 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n102 0.236924
R200 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n58 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n38 0.140076
R201 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n78 0.0916515
R202 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n91 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 0.0755
R203 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n10 0.00675
R204 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n37 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n29 0.00675
R205 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n57 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n49 0.00675
R206 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n77 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n69 0.00675
R207 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t14 141.399
R208 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t11 141.399
R209 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t10 141.399
R210 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t13 141.399
R211 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t12 140.061
R212 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t9 140.061
R213 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t15 140.061
R214 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t0 140.061
R215 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t4 134.732
R216 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t5 134.732
R217 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t1 134.732
R218 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t6 134.732
R219 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t2 134.712
R220 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t7 134.712
R221 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t8 134.712
R222 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t3 134.712
R223 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n4 8.29542
R224 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n0 6.98292
R225 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n1 6.72342
R226 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n3 5.41092
R227 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n2 3.89759
R228 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n9 3.55008
R229 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n5 3.4105
R230 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n12 3.4105
R231 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n8 3.12133
R232 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n10 1.80883
R233 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n11 1.55467
R234 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n13 1.11426
R235 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n6 0.578742
R236 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n7 0.242167
R237 VDDA.n328 VDDA.n70 10828.8
R238 VDDA.n328 VDDA.n327 10828.8
R239 VDDA.n90 VDDA.n68 10344.7
R240 VDDA.n205 VDDA.n90 10344.7
R241 VDDA.n129 VDDA.n45 9916.1
R242 VDDA.n146 VDDA.n79 9916.1
R243 VDDA.n78 VDDA.n45 9914.2
R244 VDDA.n320 VDDA.n79 9914.2
R245 VDDA.n213 VDDA.n53 9786.51
R246 VDDA.n332 VDDA.n53 9786.51
R247 VDDA.n316 VDDA.n88 8757.1
R248 VDDA.n316 VDDA.n80 8755.2
R249 VDDA.n206 VDDA.n89 8715.3
R250 VDDA.n89 VDDA.n69 8715.3
R251 VDDA.n313 VDDA.n91 8715.3
R252 VDDA.n313 VDDA.n66 8715.3
R253 VDDA.n211 VDDA.n63 8715.3
R254 VDDA.n65 VDDA.n63 8715.3
R255 VDDA.n376 VDDA.n54 7193.6
R256 VDDA.n64 VDDA.n54 7193.6
R257 VDDA.n25 VDDA.n12 4035.6
R258 VDDA.n35 VDDA.n12 4035.6
R259 VDDA.n395 VDDA.n14 3731.6
R260 VDDA.n395 VDDA.n15 3731.6
R261 VDDA.n272 VDDA.n127 3420
R262 VDDA.n216 VDDA.n127 3420
R263 VDDA.n323 VDDA.n76 3420
R264 VDDA.n77 VDDA.n76 3420
R265 VDDA.n111 VDDA.n110 2996.3
R266 VDDA.n114 VDDA.n111 2996.3
R267 VDDA.n114 VDDA.n112 2996.3
R268 VDDA.n112 VDDA.n110 2996.3
R269 VDDA.n35 VDDA.n33 2612.5
R270 VDDA.n27 VDDA.n24 2612.5
R271 VDDA.n27 VDDA.n26 2612.5
R272 VDDA.n26 VDDA.n25 2612.5
R273 VDDA.n37 VDDA.n32 2612.5
R274 VDDA.n37 VDDA.n33 2612.5
R275 VDDA.n32 VDDA.n15 2308.5
R276 VDDA.n24 VDDA.n14 2308.5
R277 VDDA.n5 VDDA.n3 2283.8
R278 VDDA.n398 VDDA.n5 2283.8
R279 VDDA.n398 VDDA.n9 2283.8
R280 VDDA.n9 VDDA.n3 2283.8
R281 VDDA.n381 VDDA.n380 1964.8
R282 VDDA.n144 VDDA.n130 1964.8
R283 VDDA.n130 VDDA.n81 1964.42
R284 VDDA.n377 VDDA.n376 1932.23
R285 VDDA.n377 VDDA.n52 1932.05
R286 VDDA.n255 VDDA.n237 1778.4
R287 VDDA.n255 VDDA.n239 1778.4
R288 VDDA.n223 VDDA.n221 1778.4
R289 VDDA.n223 VDDA.n220 1778.4
R290 VDDA.n269 VDDA.n128 1778.4
R291 VDDA.n269 VDDA.n217 1778.4
R292 VDDA.n245 VDDA.n75 1778.4
R293 VDDA.n245 VDDA.n243 1778.4
R294 VDDA.n317 VDDA.n84 1735.15
R295 VDDA.n380 VDDA.n46 1734.78
R296 VDDA.n318 VDDA.n317 1734.78
R297 VDDA.n312 VDDA.n311 1726.88
R298 VDDA.n208 VDDA.n72 1726.87
R299 VDDA.n329 VDDA.n72 1726.87
R300 VDDA.n312 VDDA.n92 1726.87
R301 VDDA.n337 VDDA.n62 1726.87
R302 VDDA.n337 VDDA.n336 1726.87
R303 VDDA.n272 VDDA.n128 1641.6
R304 VDDA.n263 VDDA.n128 1641.6
R305 VDDA.n263 VDDA.n221 1641.6
R306 VDDA.n258 VDDA.n221 1641.6
R307 VDDA.n258 VDDA.n237 1641.6
R308 VDDA.n249 VDDA.n237 1641.6
R309 VDDA.n249 VDDA.n75 1641.6
R310 VDDA.n323 VDDA.n75 1641.6
R311 VDDA.n217 VDDA.n216 1641.6
R312 VDDA.n265 VDDA.n217 1641.6
R313 VDDA.n265 VDDA.n220 1641.6
R314 VDDA.n238 VDDA.n220 1641.6
R315 VDDA.n239 VDDA.n238 1641.6
R316 VDDA.n251 VDDA.n239 1641.6
R317 VDDA.n251 VDDA.n243 1641.6
R318 VDDA.n243 VDDA.n77 1641.6
R319 VDDA.n331 VDDA.n66 1629.41
R320 VDDA.n210 VDDA.n91 1629.41
R321 VDDA.n331 VDDA.n69 1578.31
R322 VDDA.n69 VDDA.n68 1578.31
R323 VDDA.n206 VDDA.n205 1578.31
R324 VDDA.n210 VDDA.n206 1578.31
R325 VDDA.n26 VDDA.n13 1423.1
R326 VDDA.n33 VDDA.n13 1423.1
R327 VDDA.n24 VDDA.n11 1423.1
R328 VDDA.n32 VDDA.n11 1423.1
R329 VDDA.n129 VDDA.n88 1109.6
R330 VDDA.n320 VDDA.n80 1109.6
R331 VDDA.n80 VDDA.n78 1109.6
R332 VDDA.n146 VDDA.n88 1109.6
R333 VDDA.n204 VDDA.n91 1071.21
R334 VDDA.n334 VDDA.n66 1071.21
R335 VDDA.n211 VDDA.n204 1020.1
R336 VDDA.n332 VDDA.n65 1020.1
R337 VDDA.n334 VDDA.n65 1020.1
R338 VDDA.n213 VDDA.n211 1020.1
R339 VDDA.n34 VDDA.n4 756.33
R340 VDDA.n394 VDDA.n16 744.283
R341 VDDA.n394 VDDA.n17 744.283
R342 VDDA.n241 VDDA.n74 682.542
R343 VDDA.n218 VDDA.n125 682.542
R344 VDDA.n120 VDDA.n109 598.588
R345 VDDA.n120 VDDA.n119 598.588
R346 VDDA.n115 VDDA.n109 598.588
R347 VDDA.n119 VDDA.n115 598.588
R348 VDDA.n23 VDDA.n22 528.759
R349 VDDA.n34 VDDA.n31 522.542
R350 VDDA.n29 VDDA.n23 522.542
R351 VDDA.n28 VDDA.n20 522.542
R352 VDDA.n29 VDDA.n28 522.542
R353 VDDA.n39 VDDA.n38 522.542
R354 VDDA.n38 VDDA.n31 522.542
R355 VDDA.n275 VDDA.n274 507.824
R356 VDDA.n20 VDDA.n16 462.307
R357 VDDA.n39 VDDA.n17 462.307
R358 VDDA.n400 VDDA.n399 457.413
R359 VDDA.n399 VDDA.n6 457.413
R360 VDDA.n247 VDDA.n246 357.272
R361 VDDA.n246 VDDA.n242 357.272
R362 VDDA.n254 VDDA.n236 357.272
R363 VDDA.n254 VDDA.n253 357.272
R364 VDDA.n261 VDDA.n224 357.272
R365 VDDA.n224 VDDA.n219 357.272
R366 VDDA.n268 VDDA.n126 357.272
R367 VDDA.n268 VDDA.n267 357.272
R368 VDDA.n325 VDDA.n74 357.272
R369 VDDA.n274 VDDA.n125 357.272
R370 VDDA.n267 VDDA.n218 325.272
R371 VDDA.n267 VDDA.n266 325.272
R372 VDDA.n266 VDDA.n219 325.272
R373 VDDA.n240 VDDA.n219 325.272
R374 VDDA.n253 VDDA.n240 325.272
R375 VDDA.n253 VDDA.n252 325.272
R376 VDDA.n252 VDDA.n242 325.272
R377 VDDA.n242 VDDA.n241 325.272
R378 VDDA.n330 VDDA.n329 316.51
R379 VDDA.n329 VDDA.n71 316.51
R380 VDDA.n311 VDDA.n70 312.279
R381 VDDA.n327 VDDA.n326 312.24
R382 VDDA.n207 VDDA.n92 312.094
R383 VDDA.n209 VDDA.n208 307.2
R384 VDDA.n208 VDDA.n124 307.2
R385 VDDA.n401 VDDA.n400 301.748
R386 VDDA.n6 VDDA.n2 301.748
R387 VDDA.n30 VDDA.n29 281.976
R388 VDDA.n31 VDDA.n30 281.976
R389 VDDA.n40 VDDA.n20 281.976
R390 VDDA.n40 VDDA.n39 281.976
R391 VDDA.n22 VDDA.n21 275.2
R392 VDDA.n82 VDDA.n46 229.648
R393 VDDA.n84 VDDA.n44 224.754
R394 VDDA.n319 VDDA.n318 224.754
R395 VDDA.n318 VDDA.n83 224.754
R396 VDDA.n145 VDDA.n84 224.754
R397 VDDA.n336 VDDA.n55 206.352
R398 VDDA.n336 VDDA.n335 206.352
R399 VDDA.n311 VDDA.n64 205.362
R400 VDDA.n202 VDDA.n92 205.177
R401 VDDA.n203 VDDA.n62 200.282
R402 VDDA.n212 VDDA.n62 200.282
R403 VDDA.t0 VDDA.n9 174.853
R404 VDDA.t28 VDDA.n5 174.853
R405 VDDA.n402 VDDA.n2 155.107
R406 VDDA.n402 VDDA.n401 155.107
R407 VDDA.n189 VDDA.t159 139.454
R408 VDDA.n175 VDDA.t118 139.454
R409 VDDA.n189 VDDA.t140 139.454
R410 VDDA.n175 VDDA.t75 139.454
R411 VDDA.n194 VDDA.t84 139.454
R412 VDDA.n193 VDDA.t149 139.454
R413 VDDA.n170 VDDA.t55 139.454
R414 VDDA.n161 VDDA.t115 139.454
R415 VDDA.n372 VDDA.t59 139.454
R416 VDDA.n369 VDDA.t96 139.454
R417 VDDA.n371 VDDA.t62 139.454
R418 VDDA.n357 VDDA.t137 139.454
R419 VDDA.n355 VDDA.t131 139.454
R420 VDDA.n357 VDDA.t93 139.454
R421 VDDA.n355 VDDA.t90 139.454
R422 VDDA.n136 VDDA.t143 139.454
R423 VDDA.n140 VDDA.t162 139.454
R424 VDDA.n85 VDDA.t152 139.454
R425 VDDA.n86 VDDA.t168 139.454
R426 VDDA.n131 VDDA.t99 139.454
R427 VDDA.n132 VDDA.t146 139.454
R428 VDDA.n302 VDDA.t47 139.454
R429 VDDA.n304 VDDA.t43 139.454
R430 VDDA.n158 VDDA.t78 139.454
R431 VDDA.n103 VDDA.t106 139.454
R432 VDDA.n102 VDDA.t109 139.454
R433 VDDA.n231 VDDA.t81 139.454
R434 VDDA.n230 VDDA.t87 139.454
R435 VDDA.n226 VDDA.t72 139.454
R436 VDDA.n225 VDDA.t134 139.454
R437 VDDA.n198 VDDA.t165 139.454
R438 VDDA.n283 VDDA.t103 139.454
R439 VDDA.n282 VDDA.t156 139.454
R440 VDDA.n279 VDDA.t51 139.454
R441 VDDA.n278 VDDA.t112 139.454
R442 VDDA.n293 VDDA.t125 139.454
R443 VDDA.n292 VDDA.t128 139.454
R444 VDDA.n289 VDDA.t66 139.454
R445 VDDA.n288 VDDA.t69 139.454
R446 VDDA.n160 VDDA.t121 139.454
R447 VDDA.n194 VDDA.t85 135.662
R448 VDDA.n193 VDDA.t151 135.662
R449 VDDA.n103 VDDA.t107 135.662
R450 VDDA.n102 VDDA.t111 135.662
R451 VDDA.n231 VDDA.t82 135.662
R452 VDDA.n230 VDDA.t89 135.662
R453 VDDA.n226 VDDA.t73 135.662
R454 VDDA.n225 VDDA.t136 135.662
R455 VDDA.n283 VDDA.t104 135.662
R456 VDDA.n282 VDDA.t158 135.662
R457 VDDA.n279 VDDA.t53 135.662
R458 VDDA.n278 VDDA.t114 135.662
R459 VDDA.n293 VDDA.t126 135.662
R460 VDDA.n292 VDDA.t130 135.662
R461 VDDA.n289 VDDA.t67 135.662
R462 VDDA.n288 VDDA.t71 135.662
R463 VDDA.n174 VDDA.t76 135.312
R464 VDDA.n174 VDDA.t119 135.312
R465 VDDA.n373 VDDA.t61 135.312
R466 VDDA.n301 VDDA.t50 135.312
R467 VDDA.n199 VDDA.t166 135.312
R468 VDDA.n354 VDDA.t91 135.312
R469 VDDA.n354 VDDA.t132 135.312
R470 VDDA.n356 VDDA.t95 135.312
R471 VDDA.n356 VDDA.t139 135.312
R472 VDDA.n159 VDDA.t116 135.312
R473 VDDA.n188 VDDA.t142 135.312
R474 VDDA.n188 VDDA.t161 135.312
R475 VDDA.n371 VDDA.t65 135.127
R476 VDDA.n371 VDDA.t64 135.127
R477 VDDA.n85 VDDA.t155 135.127
R478 VDDA.n85 VDDA.t154 135.127
R479 VDDA.n86 VDDA.t170 135.127
R480 VDDA.n86 VDDA.t169 135.127
R481 VDDA.n131 VDDA.t102 135.127
R482 VDDA.n131 VDDA.t101 135.127
R483 VDDA.n132 VDDA.t148 135.127
R484 VDDA.n132 VDDA.t147 135.127
R485 VDDA.n160 VDDA.t124 135.127
R486 VDDA.n160 VDDA.t123 135.127
R487 VDDA.n137 VDDA.t144 135.026
R488 VDDA.n135 VDDA.t145 135.026
R489 VDDA.n139 VDDA.t164 135.026
R490 VDDA.n141 VDDA.t163 135.026
R491 VDDA.n191 VDDA.t141 134.712
R492 VDDA.n191 VDDA.t77 134.712
R493 VDDA.n192 VDDA.t79 134.712
R494 VDDA.n192 VDDA.t167 134.712
R495 VDDA.n195 VDDA.t150 134.712
R496 VDDA.n195 VDDA.t86 134.712
R497 VDDA.n172 VDDA.t57 134.712
R498 VDDA.n172 VDDA.t117 134.712
R499 VDDA.n173 VDDA.t160 134.712
R500 VDDA.n173 VDDA.t120 134.712
R501 VDDA.n49 VDDA.t244 134.712
R502 VDDA.n49 VDDA.t203 134.712
R503 VDDA.n360 VDDA.t60 134.712
R504 VDDA.n360 VDDA.t98 134.712
R505 VDDA.n359 VDDA.t138 134.712
R506 VDDA.n359 VDDA.t133 134.712
R507 VDDA.n100 VDDA.t45 134.712
R508 VDDA.n100 VDDA.t204 134.712
R509 VDDA.n150 VDDA.t211 134.712
R510 VDDA.n150 VDDA.t80 134.712
R511 VDDA.n151 VDDA.t241 134.712
R512 VDDA.n151 VDDA.t224 134.712
R513 VDDA.n152 VDDA.t220 134.712
R514 VDDA.n152 VDDA.t195 134.712
R515 VDDA.n153 VDDA.t250 134.712
R516 VDDA.n153 VDDA.t223 134.712
R517 VDDA.n93 VDDA.t219 134.712
R518 VDDA.n93 VDDA.t217 134.712
R519 VDDA.n95 VDDA.t249 134.712
R520 VDDA.n95 VDDA.t231 134.712
R521 VDDA.n96 VDDA.t239 134.712
R522 VDDA.n96 VDDA.t199 134.712
R523 VDDA.n97 VDDA.t173 134.712
R524 VDDA.n97 VDDA.t230 134.712
R525 VDDA.n98 VDDA.t229 134.712
R526 VDDA.n98 VDDA.t225 134.712
R527 VDDA.n99 VDDA.t176 134.712
R528 VDDA.n99 VDDA.t174 134.712
R529 VDDA.n58 VDDA.t94 134.712
R530 VDDA.n58 VDDA.t92 134.712
R531 VDDA.n101 VDDA.t49 134.712
R532 VDDA.n101 VDDA.t46 134.712
R533 VDDA.n104 VDDA.t110 134.712
R534 VDDA.n104 VDDA.t108 134.712
R535 VDDA.n232 VDDA.t88 134.712
R536 VDDA.n232 VDDA.t83 134.712
R537 VDDA.n227 VDDA.t135 134.712
R538 VDDA.n227 VDDA.t74 134.712
R539 VDDA.n280 VDDA.t113 134.712
R540 VDDA.n280 VDDA.t54 134.712
R541 VDDA.n284 VDDA.t157 134.712
R542 VDDA.n284 VDDA.t105 134.712
R543 VDDA.n290 VDDA.t70 134.712
R544 VDDA.n290 VDDA.t68 134.712
R545 VDDA.n294 VDDA.t129 134.712
R546 VDDA.n294 VDDA.t127 134.712
R547 VDDA.n176 VDDA.t185 134.712
R548 VDDA.n176 VDDA.t177 134.712
R549 VDDA.n177 VDDA.t246 134.712
R550 VDDA.n177 VDDA.t234 134.712
R551 VDDA.n178 VDDA.t233 134.712
R552 VDDA.n178 VDDA.t206 134.712
R553 VDDA.n179 VDDA.t212 134.712
R554 VDDA.n179 VDDA.t187 134.712
R555 VDDA.n180 VDDA.t183 134.712
R556 VDDA.n180 VDDA.t182 134.712
R557 VDDA.n181 VDDA.t245 134.712
R558 VDDA.n181 VDDA.t242 134.712
R559 VDDA.n182 VDDA.t178 134.712
R560 VDDA.n182 VDDA.t210 134.712
R561 VDDA.n183 VDDA.t237 134.712
R562 VDDA.n183 VDDA.t197 134.712
R563 VDDA.n59 VDDA.t193 134.712
R564 VDDA.n59 VDDA.t180 134.712
R565 VDDA.n60 VDDA.t172 134.712
R566 VDDA.n60 VDDA.t240 134.712
R567 VDDA.n339 VDDA.t236 134.712
R568 VDDA.n339 VDDA.t209 134.712
R569 VDDA.n340 VDDA.t222 134.712
R570 VDDA.n340 VDDA.t196 134.712
R571 VDDA.n342 VDDA.t190 134.712
R572 VDDA.n342 VDDA.t208 134.712
R573 VDDA.n343 VDDA.t252 134.712
R574 VDDA.n343 VDDA.t191 134.712
R575 VDDA.n345 VDDA.t186 134.712
R576 VDDA.n345 VDDA.t215 134.712
R577 VDDA.n346 VDDA.t248 134.712
R578 VDDA.n346 VDDA.t200 134.712
R579 VDDA.n348 VDDA.t216 134.712
R580 VDDA.n348 VDDA.t189 134.712
R581 VDDA.n349 VDDA.t201 134.712
R582 VDDA.n349 VDDA.t251 134.712
R583 VDDA.n351 VDDA.t247 134.712
R584 VDDA.n351 VDDA.t218 134.712
R585 VDDA.n352 VDDA.t232 134.712
R586 VDDA.n352 VDDA.t194 134.712
R587 VDDA.n361 VDDA.t97 134.712
R588 VDDA.n361 VDDA.t243 134.712
R589 VDDA.n362 VDDA.t192 134.712
R590 VDDA.n362 VDDA.t205 134.712
R591 VDDA.n363 VDDA.t227 134.712
R592 VDDA.n363 VDDA.t198 134.712
R593 VDDA.n364 VDDA.t235 134.712
R594 VDDA.n364 VDDA.t184 134.712
R595 VDDA.n50 VDDA.t175 134.712
R596 VDDA.n50 VDDA.t221 134.712
R597 VDDA.n47 VDDA.t202 134.712
R598 VDDA.n47 VDDA.t213 134.712
R599 VDDA.n165 VDDA.t181 134.712
R600 VDDA.n165 VDDA.t207 134.712
R601 VDDA.n164 VDDA.t214 134.712
R602 VDDA.n164 VDDA.t238 134.712
R603 VDDA.n163 VDDA.t188 134.712
R604 VDDA.n163 VDDA.t228 134.712
R605 VDDA.n162 VDDA.t226 134.712
R606 VDDA.n162 VDDA.t58 134.712
R607 VDDA.t258 VDDA.n112 117.921
R608 VDDA.t15 VDDA.n111 117.921
R609 VDDA.n386 VDDA.t1 84.6474
R610 VDDA.n7 VDDA.t29 84.6474
R611 VDDA.n404 VDDA.t255 84.6474
R612 VDDA.n1 VDDA.t264 84.6474
R613 VDDA.n274 VDDA.n273 74.7248
R614 VDDA.n273 VDDA.n126 74.7248
R615 VDDA.n262 VDDA.n261 74.7248
R616 VDDA.n259 VDDA.n236 74.7248
R617 VDDA.n248 VDDA.n247 74.7248
R618 VDDA.n325 VDDA.n324 74.7248
R619 VDDA.n262 VDDA 73.2546
R620 VDDA.n248 VDDA 73.2546
R621 VDDA.n324 VDDA 73.2546
R622 VDDA.n397 VDDA.t0 71.3334
R623 VDDA.n397 VDDA.t28 71.3334
R624 VDDA.n36 VDDA.t254 64.1959
R625 VDDA VDDA.n260 50.2491
R626 VDDA.n108 VDDA.t16 49.8991
R627 VDDA.n116 VDDA.t262 49.8991
R628 VDDA.n397 VDDA.n10 49.2055
R629 VDDA.n392 VDDA.t259 48.2714
R630 VDDA.n392 VDDA.t266 48.2714
R631 VDDA.n19 VDDA.t267 48.2714
R632 VDDA.n19 VDDA.t263 48.2714
R633 VDDA.n113 VDDA.t258 48.1348
R634 VDDA.n113 VDDA.t15 48.1348
R635 VDDA.n383 VDDA.n382 47.9922
R636 VDDA.n401 VDDA.n4 41.6919
R637 VDDA.n22 VDDA.n2 41.6919
R638 VDDA.n21 VDDA.n4 35.0123
R639 VDDA.t179 VDDA.t171 34.0455
R640 VDDA.t20 VDDA.t8 34.0455
R641 VDDA.t260 VDDA.t56 33.5928
R642 VDDA.t18 VDDA.t24 32.5062
R643 VDDA.n222 VDDA.t25 30.967
R644 VDDA.n244 VDDA.t40 30.6048
R645 VDDA.t153 VDDA.n214 28.9077
R646 VDDA.n215 VDDA.t52 28.2642
R647 VDDA.t6 VDDA.t7 26.3491
R648 VDDA.t31 VDDA.t39 25.987
R649 VDDA.t48 VDDA.n321 23.5422
R650 VDDA.n270 VDDA.t38 23.3612
R651 VDDA.t3 VDDA.t2 23.3612
R652 VDDA.n260 VDDA.n259 23.0059
R653 VDDA.t256 VDDA.t23 22.9084
R654 VDDA.t261 VDDA.t19 21.8219
R655 VDDA.t36 VDDA.t21 21.8219
R656 VDDA.t12 VDDA.n396 21.5134
R657 VDDA.n396 VDDA.t254 21.5134
R658 VDDA.t5 VDDA.t42 21.4597
R659 VDDA.t30 VDDA.t253 18.4717
R660 VDDA.t39 VDDA.n256 17.2041
R661 VDDA.n256 VDDA.t7 16.8419
R662 VDDA.n120 VDDA.n110 16.8187
R663 VDDA.n113 VDDA.n110 16.8187
R664 VDDA.n115 VDDA.n114 16.8187
R665 VDDA.n114 VDDA.n113 16.8187
R666 VDDA.n402 VDDA.n3 16.8187
R667 VDDA.n397 VDDA.n3 16.8187
R668 VDDA.n399 VDDA.n398 16.8187
R669 VDDA.n398 VDDA.n397 16.8187
R670 VDDA.t4 VDDA.t41 15.6648
R671 VDDA.t10 VDDA.t100 15.4837
R672 VDDA.t27 VDDA.t34 15.3026
R673 VDDA.n397 VDDA.t12 14.9909
R674 VDDA.t44 VDDA.t10 14.5783
R675 VDDA.t33 VDDA.t30 14.2161
R676 VDDA.n123 VDDA.n122 13.8332
R677 VDDA.t40 VDDA.t5 12.5863
R678 VDDA.n314 VDDA.t265 12.4052
R679 VDDA.t25 VDDA.t36 12.2241
R680 VDDA.n271 VDDA.t261 11.6808
R681 VDDA.n264 VDDA.t14 11.6808
R682 VDDA.n264 VDDA.t37 11.6808
R683 VDDA.n257 VDDA.t27 11.6808
R684 VDDA.n250 VDDA.t4 11.6808
R685 VDDA.n322 VDDA.t11 11.6808
R686 VDDA.n322 VDDA.t17 11.6808
R687 VDDA.n204 VDDA.n203 11.563
R688 VDDA.n214 VDDA.n204 11.563
R689 VDDA.n213 VDDA.n212 11.563
R690 VDDA.n214 VDDA.n213 11.563
R691 VDDA.n332 VDDA.n55 11.563
R692 VDDA.n333 VDDA.n332 11.563
R693 VDDA.n335 VDDA.n334 11.563
R694 VDDA.n334 VDDA.n333 11.563
R695 VDDA.t32 VDDA.t256 11.1376
R696 VDDA.t24 VDDA.n270 10.6848
R697 VDDA.n146 VDDA.n145 10.2783
R698 VDDA.n147 VDDA.n146 10.2783
R699 VDDA.n129 VDDA.n44 10.2783
R700 VDDA.n147 VDDA.n129 10.2783
R701 VDDA.n83 VDDA.n78 10.2783
R702 VDDA.n321 VDDA.n78 10.2783
R703 VDDA.n320 VDDA.n319 10.2783
R704 VDDA.n321 VDDA.n320 10.2783
R705 VDDA.t56 VDDA.n215 9.59829
R706 VDDA.t14 VDDA.t33 9.14556
R707 VDDA.n87 VDDA.n86 8.96925
R708 VDDA.n131 VDDA.n87 8.96717
R709 VDDA.n139 VDDA.n138 8.84008
R710 VDDA.n138 VDDA.n137 8.83592
R711 VDDA.n21 VDDA.n12 8.81002
R712 VDDA.n396 VDDA.n12 8.81002
R713 VDDA.n30 VDDA.n13 8.81002
R714 VDDA.n396 VDDA.n13 8.81002
R715 VDDA.n395 VDDA.n394 8.81002
R716 VDDA.n396 VDDA.n395 8.81002
R717 VDDA.n40 VDDA.n11 8.81002
R718 VDDA.n396 VDDA.n11 8.81002
R719 VDDA.n315 VDDA.t13 8.78338
R720 VDDA.t17 VDDA.t44 8.78338
R721 VDDA.n400 VDDA.n5 8.40959
R722 VDDA.n9 VDDA.n6 8.40959
R723 VDDA.t34 VDDA.t31 8.05902
R724 VDDA.n205 VDDA.n124 7.70883
R725 VDDA.n214 VDDA.n205 7.70883
R726 VDDA.n71 VDDA.n68 7.70883
R727 VDDA.n333 VDDA.n68 7.70883
R728 VDDA.n331 VDDA.n330 7.70883
R729 VDDA.n333 VDDA.n331 7.70883
R730 VDDA.n241 VDDA.n77 7.70883
R731 VDDA.n322 VDDA.n77 7.70883
R732 VDDA.n252 VDDA.n251 7.70883
R733 VDDA.n251 VDDA.n250 7.70883
R734 VDDA.n240 VDDA.n238 7.70883
R735 VDDA.n257 VDDA.n238 7.70883
R736 VDDA.n266 VDDA.n265 7.70883
R737 VDDA.n265 VDDA.n264 7.70883
R738 VDDA.n218 VDDA.n216 7.70883
R739 VDDA.n271 VDDA.n216 7.70883
R740 VDDA.n324 VDDA.n323 7.70883
R741 VDDA.n323 VDDA.n322 7.70883
R742 VDDA.n249 VDDA.n248 7.70883
R743 VDDA.n250 VDDA.n249 7.70883
R744 VDDA.n259 VDDA.n258 7.70883
R745 VDDA.n258 VDDA.n257 7.70883
R746 VDDA.n263 VDDA.n262 7.70883
R747 VDDA.n264 VDDA.n263 7.70883
R748 VDDA.n273 VDDA.n272 7.70883
R749 VDDA.n272 VDDA.n271 7.70883
R750 VDDA.n210 VDDA.n209 7.70883
R751 VDDA.n214 VDDA.n210 7.70883
R752 VDDA.t41 VDDA.t6 7.69684
R753 VDDA.n257 VDDA.t22 7.06302
R754 VDDA.n224 VDDA.n223 6.85235
R755 VDDA.n223 VDDA.n222 6.85235
R756 VDDA.n255 VDDA.n254 6.85235
R757 VDDA.n256 VDDA.n255 6.85235
R758 VDDA.n269 VDDA.n268 6.85235
R759 VDDA.n270 VDDA.n269 6.85235
R760 VDDA.n246 VDDA.n245 6.85235
R761 VDDA.n245 VDDA.n244 6.85235
R762 VDDA.n76 VDDA.n74 6.85235
R763 VDDA.n76 VDDA.n67 6.85235
R764 VDDA.n127 VDDA.n125 6.85235
R765 VDDA.n215 VDDA.n127 6.85235
R766 VDDA.n46 VDDA 6.4005
R767 VDDA.n235 VDDA.n229 6.33487
R768 VDDA.n235 VDDA.n234 6.33487
R769 VDDA.n287 VDDA.n286 6.33487
R770 VDDA.n296 VDDA.n287 6.33487
R771 VDDA.t171 VDDA.t13 6.06703
R772 VDDA.n329 VDDA.n328 6.02403
R773 VDDA.n336 VDDA.n54 6.02403
R774 VDDA.n389 VDDA.n388 5.93473
R775 VDDA.t9 VDDA.t257 5.70485
R776 VDDA.t8 VDDA.t3 5.70485
R777 VDDA.n112 VDDA.n109 5.60656
R778 VDDA.n119 VDDA.n111 5.60656
R779 VDDA.n16 VDDA.n14 5.28621
R780 VDDA.n14 VDDA.n10 5.28621
R781 VDDA.n17 VDDA.n15 5.28621
R782 VDDA.n36 VDDA.n15 5.28621
R783 VDDA.n214 VDDA.n147 5.17455
R784 VDDA.n330 VDDA.n70 5.04292
R785 VDDA.n327 VDDA.n71 5.04292
R786 VDDA.n376 VDDA.n55 5.04292
R787 VDDA.n335 VDDA.n64 5.04292
R788 VDDA.t2 VDDA.t9 4.98048
R789 VDDA.n381 VDDA.n44 4.89462
R790 VDDA.n319 VDDA.n81 4.89462
R791 VDDA.n83 VDDA.n82 4.89462
R792 VDDA.n145 VDDA.n144 4.89462
R793 VDDA.n209 VDDA.n207 4.89462
R794 VDDA.n275 VDDA.n124 4.89462
R795 VDDA.n203 VDDA.n202 4.89462
R796 VDDA.n212 VDDA.n52 4.89462
R797 VDDA.n35 VDDA.n34 4.6255
R798 VDDA.n36 VDDA.n35 4.6255
R799 VDDA.n28 VDDA.n27 4.6255
R800 VDDA.n27 VDDA.n10 4.6255
R801 VDDA.n25 VDDA.n23 4.6255
R802 VDDA.n25 VDDA.n10 4.6255
R803 VDDA.n38 VDDA.n37 4.6255
R804 VDDA.n37 VDDA.n36 4.6255
R805 VDDA.t22 VDDA.t265 4.6183
R806 VDDA.t63 VDDA.t48 3.89394
R807 VDDA.n244 VDDA.t20 3.44122
R808 VDDA.n222 VDDA.t179 3.07904
R809 VDDA.n118 VDDA.n117 2.44894
R810 VDDA.n315 VDDA.n314 2.17358
R811 VDDA.n118 VDDA.n108 2.04581
R812 VDDA.n116 VDDA.n107 2.04581
R813 VDDA.t42 VDDA.t11 1.90195
R814 VDDA.n234 VDDA.n73 1.86994
R815 VDDA.n122 VDDA.n107 1.78175
R816 VDDA.n135 VDDA.n134 1.74633
R817 VDDA.t19 VDDA.t18 1.53977
R818 VDDA.t21 VDDA.t37 1.53977
R819 VDDA VDDA.n126 1.47077
R820 VDDA.n261 VDDA 1.47077
R821 VDDA VDDA.n236 1.47077
R822 VDDA.n247 VDDA 1.47077
R823 VDDA.n387 VDDA.n386 1.45988
R824 VDDA.n7 VDDA.n0 1.45988
R825 VDDA.n384 VDDA.n41 1.43637
R826 VDDA.n385 VDDA.n384 1.40704
R827 VDDA.n41 VDDA.n18 1.388
R828 VDDA.n380 VDDA.n45 1.3811
R829 VDDA.n315 VDDA.n45 1.3811
R830 VDDA.n130 VDDA.n79 1.3811
R831 VDDA.n315 VDDA.n79 1.3811
R832 VDDA.n260 VDDA.n90 1.3811
R833 VDDA.n314 VDDA.n90 1.3811
R834 VDDA.n313 VDDA.n312 1.3811
R835 VDDA.n314 VDDA.n313 1.3811
R836 VDDA.n377 VDDA.n53 1.3811
R837 VDDA.n314 VDDA.n53 1.3811
R838 VDDA.n89 VDDA.n72 1.37087
R839 VDDA.n314 VDDA.n89 1.37087
R840 VDDA.n337 VDDA.n63 1.37087
R841 VDDA.n314 VDDA.n63 1.37087
R842 VDDA.n317 VDDA.n316 1.36079
R843 VDDA.n316 VDDA.n315 1.36079
R844 VDDA.n326 VDDA 1.34471
R845 VDDA.n374 VDDA.n57 1.32758
R846 VDDA.n389 VDDA.n385 1.32758
R847 VDDA.n300 VDDA.n298 1.30308
R848 VDDA.n298 VDDA.n297 1.30306
R849 VDDA.n297 VDDA.n73 1.30208
R850 VDDA.n200 VDDA.n106 1.29217
R851 VDDA.n277 VDDA.n106 1.29217
R852 VDDA.n277 VDDA.n276 1.29217
R853 VDDA.t26 VDDA.t38 1.26813
R854 VDDA.n134 VDDA.n133 1.24425
R855 VDDA.n143 VDDA.n43 1.24425
R856 VDDA.n382 VDDA.n43 1.24425
R857 VDDA.n133 VDDA.n57 1.24425
R858 VDDA.n405 VDDA.n0 1.19112
R859 VDDA.n276 VDDA.n123 1.15755
R860 VDDA.n391 VDDA 1.02231
R861 VDDA.n391 VDDA.n18 0.998346
R862 VDDA.n157 VDDA.n156 0.947451
R863 VDDA.n306 VDDA.n305 0.947451
R864 VDDA.n156 VDDA.n155 0.91925
R865 VDDA.n155 VDDA.n154 0.91925
R866 VDDA.n154 VDDA.n94 0.91925
R867 VDDA.n310 VDDA.n94 0.91925
R868 VDDA.n310 VDDA.n309 0.91925
R869 VDDA.n309 VDDA.n308 0.91925
R870 VDDA.n308 VDDA.n307 0.91925
R871 VDDA.n307 VDDA.n306 0.91925
R872 VDDA.n187 VDDA.n186 0.91925
R873 VDDA.n186 VDDA.n185 0.91925
R874 VDDA.n185 VDDA.n184 0.91925
R875 VDDA.n184 VDDA.n61 0.91925
R876 VDDA.n344 VDDA.n341 0.91925
R877 VDDA.n347 VDDA.n344 0.91925
R878 VDDA.n350 VDDA.n347 0.91925
R879 VDDA.n353 VDDA.n350 0.91925
R880 VDDA.n375 VDDA.n374 0.919194
R881 VDDA.n250 VDDA.t35 0.905952
R882 VDDA.n375 VDDA.n56 0.847727
R883 VDDA.n299 VDDA.n56 0.846749
R884 VDDA.n300 VDDA.n299 0.846726
R885 VDDA.n201 VDDA.n149 0.837038
R886 VDDA.n201 VDDA.n200 0.837038
R887 VDDA.n148 VDDA.n42 0.837038
R888 VDDA.n149 VDDA.n148 0.837038
R889 VDDA.n117 VDDA.n115 0.7755
R890 VDDA.n121 VDDA.n120 0.7755
R891 VDDA.n403 VDDA.n402 0.7755
R892 VDDA.n399 VDDA.n8 0.7755
R893 VDDA.n142 VDDA.n141 0.7005
R894 VDDA.n122 VDDA.n121 0.667688
R895 VDDA.n143 VDDA.n142 0.658833
R896 VDDA.n85 VDDA.n43 0.63175
R897 VDDA.n133 VDDA.n132 0.63175
R898 VDDA.n390 VDDA.n389 0.623
R899 VDDA.n202 VDDA.n201 0.6205
R900 VDDA.n376 VDDA.n375 0.6205
R901 VDDA.n299 VDDA.n64 0.6205
R902 VDDA.n148 VDDA.n52 0.6205
R903 VDDA VDDA.n390 0.6015
R904 VDDA.n286 VDDA.n277 0.577063
R905 VDDA.n297 VDDA.n296 0.569374
R906 VDDA.t52 VDDA.t122 0.562896
R907 VDDA.n134 VDDA.n81 0.547559
R908 VDDA.n144 VDDA.n143 0.547559
R909 VDDA.n382 VDDA.n381 0.547559
R910 VDDA.n82 VDDA.n57 0.547559
R911 VDDA.n229 VDDA.n123 0.545851
R912 VDDA.n388 VDDA.n387 0.54401
R913 VDDA.n271 VDDA.t32 0.543771
R914 VDDA.n188 VDDA.n187 0.528735
R915 VDDA.n354 VDDA.n353 0.528735
R916 VDDA.n168 VDDA.n167 0.51137
R917 VDDA.n167 VDDA.n166 0.51137
R918 VDDA.n166 VDDA.n48 0.51137
R919 VDDA.n378 VDDA.n51 0.51137
R920 VDDA.n365 VDDA.n51 0.51137
R921 VDDA.n366 VDDA.n365 0.51137
R922 VDDA.n367 VDDA.n366 0.51137
R923 VDDA.n368 VDDA.n367 0.495392
R924 VDDA.n169 VDDA.n168 0.495392
R925 VDDA.n379 VDDA.n48 0.495065
R926 VDDA.n393 VDDA.n392 0.49364
R927 VDDA.n385 VDDA.n19 0.49364
R928 VDDA.n338 VDDA.n61 0.459875
R929 VDDA.n341 VDDA.n338 0.459875
R930 VDDA.t23 VDDA.t260 0.453226
R931 VDDA.n394 VDDA.n393 0.443357
R932 VDDA.n385 VDDA.n40 0.443357
R933 VDDA.n400 VDDA.n0 0.423227
R934 VDDA.n387 VDDA.n6 0.423227
R935 VDDA.n207 VDDA.n106 0.404848
R936 VDDA.n298 VDDA.n70 0.404848
R937 VDDA.n327 VDDA.n73 0.404848
R938 VDDA.n276 VDDA.n275 0.404848
R939 VDDA.n117 VDDA.n116 0.403625
R940 VDDA.n121 VDDA.n108 0.403625
R941 VDDA.n386 VDDA.n8 0.403625
R942 VDDA.n8 VDDA.n7 0.403625
R943 VDDA.n403 VDDA.n1 0.403625
R944 VDDA.n404 VDDA.n403 0.403625
R945 VDDA.n101 VDDA.n58 0.346537
R946 VDDA.n360 VDDA.n359 0.346537
R947 VDDA.n173 VDDA.n172 0.346537
R948 VDDA.n192 VDDA.n191 0.346537
R949 VDDA VDDA.n18 0.299149
R950 VDDA.n119 VDDA.n118 0.291125
R951 VDDA.n109 VDDA.n107 0.291125
R952 VDDA.n196 VDDA.n193 0.288543
R953 VDDA.n196 VDDA.n194 0.288543
R954 VDDA.n105 VDDA.n102 0.288543
R955 VDDA.n105 VDDA.n103 0.288543
R956 VDDA.n233 VDDA.n230 0.288543
R957 VDDA.n233 VDDA.n231 0.288543
R958 VDDA.n228 VDDA.n225 0.288543
R959 VDDA.n228 VDDA.n226 0.288543
R960 VDDA.n285 VDDA.n282 0.288543
R961 VDDA.n285 VDDA.n283 0.288543
R962 VDDA.n281 VDDA.n278 0.288543
R963 VDDA.n281 VDDA.n279 0.288543
R964 VDDA.n295 VDDA.n292 0.288543
R965 VDDA.n295 VDDA.n293 0.288543
R966 VDDA.n291 VDDA.n288 0.288543
R967 VDDA.n291 VDDA.n289 0.288543
R968 VDDA.n383 VDDA.n42 0.285826
R969 VDDA.n390 VDDA.n16 0.274029
R970 VDDA.n41 VDDA.n17 0.274029
R971 VDDA.n384 VDDA.n383 0.273356
R972 VDDA.n405 VDDA.n404 0.26925
R973 VDDA.n142 VDDA 0.261311
R974 VDDA.n156 VDDA.n151 0.255835
R975 VDDA.n155 VDDA.n152 0.255835
R976 VDDA.n154 VDDA.n153 0.255835
R977 VDDA.n94 VDDA.n93 0.255835
R978 VDDA.n310 VDDA.n95 0.255835
R979 VDDA.n309 VDDA.n96 0.255835
R980 VDDA.n308 VDDA.n97 0.255835
R981 VDDA.n307 VDDA.n98 0.255835
R982 VDDA.n306 VDDA.n99 0.255835
R983 VDDA.n187 VDDA.n176 0.255835
R984 VDDA.n187 VDDA.n177 0.255835
R985 VDDA.n186 VDDA.n178 0.255835
R986 VDDA.n186 VDDA.n179 0.255835
R987 VDDA.n185 VDDA.n180 0.255835
R988 VDDA.n185 VDDA.n181 0.255835
R989 VDDA.n184 VDDA.n182 0.255835
R990 VDDA.n184 VDDA.n183 0.255835
R991 VDDA.n61 VDDA.n59 0.255835
R992 VDDA.n61 VDDA.n60 0.255835
R993 VDDA.n341 VDDA.n339 0.255835
R994 VDDA.n341 VDDA.n340 0.255835
R995 VDDA.n344 VDDA.n342 0.255835
R996 VDDA.n344 VDDA.n343 0.255835
R997 VDDA.n347 VDDA.n345 0.255835
R998 VDDA.n347 VDDA.n346 0.255835
R999 VDDA.n350 VDDA.n348 0.255835
R1000 VDDA.n350 VDDA.n349 0.255835
R1001 VDDA.n353 VDDA.n351 0.255835
R1002 VDDA.n353 VDDA.n352 0.255835
R1003 VDDA.n303 VDDA.n105 0.232207
R1004 VDDA.n197 VDDA.n196 0.232207
R1005 VDDA.n157 VDDA.n150 0.227634
R1006 VDDA.n305 VDDA.n100 0.227634
R1007 VDDA.n303 VDDA.n101 0.227634
R1008 VDDA.n197 VDDA.n192 0.227634
R1009 VDDA.n378 VDDA.n49 0.225348
R1010 VDDA.n367 VDDA.n362 0.225348
R1011 VDDA.n366 VDDA.n363 0.225348
R1012 VDDA.n365 VDDA.n364 0.225348
R1013 VDDA.n51 VDDA.n50 0.225348
R1014 VDDA.n48 VDDA.n47 0.225348
R1015 VDDA.n166 VDDA.n165 0.225348
R1016 VDDA.n167 VDDA.n164 0.225348
R1017 VDDA.n168 VDDA.n163 0.225348
R1018 VDDA.n388 VDDA.n1 0.20675
R1019 VDDA.n234 VDDA.n233 0.204006
R1020 VDDA.n229 VDDA.n228 0.204006
R1021 VDDA.n286 VDDA.n281 0.204006
R1022 VDDA.n286 VDDA.n285 0.204006
R1023 VDDA.n296 VDDA.n291 0.204006
R1024 VDDA.n296 VDDA.n295 0.204006
R1025 VDDA.n200 VDDA.n199 0.192606
R1026 VDDA.n174 VDDA.n149 0.186547
R1027 VDDA.n105 VDDA.n104 0.186476
R1028 VDDA.n233 VDDA.n232 0.186476
R1029 VDDA.n228 VDDA.n227 0.186476
R1030 VDDA.n281 VDDA.n280 0.186476
R1031 VDDA.n285 VDDA.n284 0.186476
R1032 VDDA.n291 VDDA.n290 0.186476
R1033 VDDA.n295 VDDA.n294 0.186476
R1034 VDDA.n196 VDDA.n195 0.186476
R1035 VDDA.n301 VDDA.n300 0.184889
R1036 VDDA.n321 VDDA.n67 0.18159
R1037 VDDA.n356 VDDA.n56 0.178804
R1038 VDDA.n358 VDDA.n58 0.168945
R1039 VDDA.n370 VDDA.n360 0.168945
R1040 VDDA.n359 VDDA.n358 0.168945
R1041 VDDA.n368 VDDA.n361 0.168945
R1042 VDDA.n169 VDDA.n162 0.168945
R1043 VDDA.n172 VDDA.n171 0.168945
R1044 VDDA.n190 VDDA.n173 0.168945
R1045 VDDA.n191 VDDA.n190 0.168945
R1046 VDDA.n326 VDDA.n325 0.127387
R1047 VDDA.t122 VDDA.t153 0.112979
R1048 VDDA.n302 VDDA.n301 0.105208
R1049 VDDA.n199 VDDA.n198 0.105208
R1050 VDDA.n358 VDDA.n355 0.10357
R1051 VDDA.n358 VDDA.n357 0.10357
R1052 VDDA.n190 VDDA.n175 0.10357
R1053 VDDA.n190 VDDA.n189 0.10357
R1054 VDDA.n369 VDDA.n368 0.0915853
R1055 VDDA.n370 VDDA.n369 0.0915853
R1056 VDDA.n171 VDDA.n161 0.0915853
R1057 VDDA.n171 VDDA.n170 0.0915853
R1058 VDDA.n170 VDDA.n169 0.0915853
R1059 VDDA.t253 VDDA.t26 0.0910452
R1060 VDDA.t257 VDDA.t35 0.0910452
R1061 VDDA.t100 VDDA.t63 0.0910452
R1062 VDDA.n333 VDDA.n67 0.0910452
R1063 VDDA.n159 VDDA.n42 0.087051
R1064 VDDA.n197 VDDA.n158 0.086539
R1065 VDDA.n158 VDDA.n157 0.086539
R1066 VDDA.n305 VDDA.n304 0.086539
R1067 VDDA.n304 VDDA.n303 0.086539
R1068 VDDA.n303 VDDA.n302 0.086539
R1069 VDDA.n198 VDDA.n197 0.086539
R1070 VDDA.n287 VDDA.n72 0.0731563
R1071 VDDA.n260 VDDA.n235 0.0731563
R1072 VDDA.n312 VDDA.n310 0.0731563
R1073 VDDA.n338 VDDA.n337 0.0731563
R1074 VDDA.n378 VDDA.n377 0.0731563
R1075 VDDA.n138 VDDA.n130 0.072593
R1076 VDDA.n317 VDDA.n87 0.072593
R1077 VDDA.n380 VDDA.n379 0.072593
R1078 VDDA.n355 VDDA.n354 0.0712237
R1079 VDDA.n357 VDDA.n356 0.0712237
R1080 VDDA.n175 VDDA.n174 0.0712237
R1081 VDDA.n189 VDDA.n188 0.0712237
R1082 VDDA.n371 VDDA.n370 0.0707519
R1083 VDDA.n373 VDDA.n372 0.063
R1084 VDDA.n160 VDDA.n159 0.0605775
R1085 VDDA.n137 VDDA.n136 0.0575652
R1086 VDDA.n136 VDDA.n135 0.0575652
R1087 VDDA.n141 VDDA.n140 0.0575652
R1088 VDDA.n140 VDDA.n139 0.0575652
R1089 VDDA VDDA.n405 0.047375
R1090 VDDA.n372 VDDA.n371 0.0213333
R1091 VDDA.n379 VDDA.n378 0.0168043
R1092 VDDA.n374 VDDA.n373 0.0116434
R1093 VDDA.n393 VDDA.n391 0.00812195
R1094 VDDA.n161 VDDA.n160 0.00292248
R1095 VDDA.n86 VDDA.n85 0.00258333
R1096 VDDA.n132 VDDA.n131 0.00258333
R1097 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n62 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t36 214.787
R1098 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n63 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t16 214.787
R1099 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n62 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t66 214.011
R1100 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n63 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t42 214.011
R1101 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n73 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t24 142.488
R1102 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n49 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t37 142.488
R1103 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n42 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t33 142.488
R1104 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n29 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t15 142.488
R1105 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n22 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t86 142.488
R1106 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n10 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t32 142.488
R1107 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n3 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t21 142.488
R1108 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n73 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t46 141.704
R1109 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n74 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t47 141.704
R1110 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n75 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t80 141.704
R1111 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n76 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t83 141.704
R1112 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n77 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t48 141.704
R1113 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n78 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t77 141.704
R1114 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n79 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t57 141.704
R1115 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n80 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t31 141.704
R1116 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n81 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t53 141.704
R1117 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n82 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t75 141.704
R1118 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n83 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t4 141.704
R1119 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n72 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t6 141.704
R1120 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n71 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t52 141.704
R1121 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n70 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t85 141.704
R1122 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n69 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t87 141.704
R1123 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n68 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t34 141.704
R1124 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n67 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t58 141.704
R1125 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n66 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t84 141.704
R1126 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n65 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t10 141.704
R1127 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n49 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t62 141.704
R1128 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n50 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t64 141.704
R1129 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n51 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t20 141.704
R1130 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n52 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t22 141.704
R1131 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n53 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t65 141.704
R1132 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n54 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t19 141.704
R1133 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n55 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t78 141.704
R1134 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n56 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t43 141.704
R1135 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n57 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t72 141.704
R1136 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n58 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t18 141.704
R1137 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n59 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t28 141.704
R1138 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n48 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t29 141.704
R1139 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n47 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t70 141.704
R1140 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n46 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t26 141.704
R1141 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n45 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t27 141.704
R1142 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n44 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t49 141.704
R1143 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n43 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t82 141.704
R1144 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n42 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t25 141.704
R1145 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n29 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t39 141.704
R1146 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n30 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t40 141.704
R1147 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n31 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t69 141.704
R1148 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n32 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t71 141.704
R1149 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n33 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t41 141.704
R1150 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n34 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t68 141.704
R1151 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n35 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t50 141.704
R1152 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n36 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t23 141.704
R1153 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n37 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t45 141.704
R1154 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n38 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t67 141.704
R1155 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n39 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t79 141.704
R1156 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n28 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t81 141.704
R1157 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n27 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t44 141.704
R1158 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n26 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t74 141.704
R1159 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n25 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t76 141.704
R1160 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n24 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t30 141.704
R1161 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n23 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t51 141.704
R1162 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n22 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t73 141.704
R1163 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n10 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t54 141.704
R1164 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n11 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t56 141.704
R1165 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n12 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t8 141.704
R1166 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n13 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t9 141.704
R1167 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n14 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t55 141.704
R1168 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n15 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t7 141.704
R1169 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n16 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t61 141.704
R1170 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n17 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t35 141.704
R1171 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n18 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t60 141.704
R1172 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n19 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t5 141.704
R1173 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n20 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t14 141.704
R1174 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n9 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t17 141.704
R1175 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n8 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t59 141.704
R1176 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n7 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t12 141.704
R1177 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n6 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t13 141.704
R1178 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n5 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t38 141.704
R1179 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n4 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t63 141.704
R1180 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n3 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t11 141.704
R1181 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n87 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n2 119.186
R1182 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n1 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n0 119.186
R1183 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n2 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t1 15.3866
R1184 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n2 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t2 15.3866
R1185 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n0 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t0 15.3866
R1186 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n0 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t3 15.3866
R1187 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n87 10.5297
R1188 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n63 7.95883
R1189 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n64 opa_input_and_self_bias_0/cm_pcell3_0.VB2 6.74425
R1190 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n86 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n85 6.37582
R1191 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n87 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n86 5.23592
R1192 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n86 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n1 5.23592
R1193 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n41 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n21 4.22517
R1194 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n65 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n64 4.13592
R1195 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n41 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n40 3.4105
R1196 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n61 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n60 3.4105
R1197 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n85 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n84 3.4105
R1198 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n64 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n62 0.973417
R1199 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n85 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n61 0.815167
R1200 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n66 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n65 0.783833
R1201 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n67 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n66 0.783833
R1202 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n68 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n67 0.783833
R1203 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n69 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n68 0.783833
R1204 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n70 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n69 0.783833
R1205 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n71 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n70 0.783833
R1206 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n72 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n71 0.783833
R1207 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n83 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n82 0.783833
R1208 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n82 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n81 0.783833
R1209 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n81 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n80 0.783833
R1210 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n80 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n79 0.783833
R1211 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n79 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n78 0.783833
R1212 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n78 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n77 0.783833
R1213 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n77 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n76 0.783833
R1214 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n76 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n75 0.783833
R1215 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n75 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n74 0.783833
R1216 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n74 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n73 0.783833
R1217 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n43 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n42 0.783833
R1218 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n44 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n43 0.783833
R1219 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n45 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n44 0.783833
R1220 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n46 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n45 0.783833
R1221 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n47 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n46 0.783833
R1222 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n48 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n47 0.783833
R1223 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n59 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n58 0.783833
R1224 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n58 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n57 0.783833
R1225 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n57 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n56 0.783833
R1226 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n56 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n55 0.783833
R1227 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n55 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n54 0.783833
R1228 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n54 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n53 0.783833
R1229 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n53 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n52 0.783833
R1230 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n52 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n51 0.783833
R1231 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n51 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n50 0.783833
R1232 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n50 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n49 0.783833
R1233 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n23 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n22 0.783833
R1234 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n24 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n23 0.783833
R1235 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n25 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n24 0.783833
R1236 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n26 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n25 0.783833
R1237 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n27 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n26 0.783833
R1238 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n28 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n27 0.783833
R1239 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n39 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n38 0.783833
R1240 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n38 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n37 0.783833
R1241 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n37 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n36 0.783833
R1242 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n36 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n35 0.783833
R1243 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n35 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n34 0.783833
R1244 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n34 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n33 0.783833
R1245 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n33 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n32 0.783833
R1246 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n32 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n31 0.783833
R1247 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n31 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n30 0.783833
R1248 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n30 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n29 0.783833
R1249 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n4 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n3 0.783833
R1250 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n5 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n4 0.783833
R1251 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n6 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n5 0.783833
R1252 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n7 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n6 0.783833
R1253 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n8 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n7 0.783833
R1254 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n9 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n8 0.783833
R1255 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n20 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n19 0.783833
R1256 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n19 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n18 0.783833
R1257 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n18 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n17 0.783833
R1258 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n17 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n16 0.783833
R1259 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n16 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n15 0.783833
R1260 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n15 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n14 0.783833
R1261 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n14 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n13 0.783833
R1262 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n13 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n12 0.783833
R1263 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n12 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n11 0.783833
R1264 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n11 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n10 0.783833
R1265 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n84 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n72 0.777583
R1266 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n60 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n48 0.777583
R1267 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n40 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n28 0.777583
R1268 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n21 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n9 0.777583
R1269 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n61 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n41 0.39003
R1270 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n1 0.063
R1271 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n84 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n83 0.00675
R1272 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n60 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n59 0.00675
R1273 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n40 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n39 0.00675
R1274 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n21 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n20 0.00675
R1275 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n20 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t1 244.856
R1276 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n21 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t3 222.089
R1277 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n8 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t6 134.738
R1278 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n8 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t8 134.738
R1279 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n10 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t15 134.738
R1280 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n10 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t19 134.738
R1281 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n1 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t20 134.734
R1282 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n1 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t7 134.734
R1283 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n2 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t10 134.734
R1284 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n2 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t22 134.734
R1285 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n4 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t16 134.734
R1286 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n4 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t13 134.734
R1287 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n6 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t11 134.734
R1288 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n6 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t12 134.734
R1289 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n11 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t9 134.734
R1290 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n11 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t4 134.734
R1291 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n13 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t14 134.734
R1292 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n13 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t18 134.734
R1293 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n15 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t5 134.734
R1294 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n15 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t21 134.734
R1295 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n17 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t23 134.734
R1296 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n17 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t17 134.734
R1297 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n23 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t0 15.2609
R1298 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n0 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t24 15.2609
R1299 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n22 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n0 11.485
R1300 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n24 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n23 11.0892
R1301 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n20 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n19 9.71425
R1302 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n3 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n1 7.63383
R1303 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n12 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n10 7.63383
R1304 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n19 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n18 7.15217
R1305 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n19 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n9 6.46995
R1306 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n9 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n8 4.5005
R1307 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n7 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n6 4.5005
R1308 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n5 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n4 4.5005
R1309 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n3 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n2 4.5005
R1310 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n18 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n17 4.5005
R1311 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n16 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n15 4.5005
R1312 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n14 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n13 4.5005
R1313 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n12 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n11 4.5005
R1314 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n23 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t25 4.23377
R1315 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n0 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t2 4.23377
R1316 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n9 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n7 3.13383
R1317 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n7 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n5 3.13383
R1318 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n5 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n3 3.13383
R1319 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n18 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n16 3.13383
R1320 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n16 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n14 3.13383
R1321 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n14 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n12 3.13383
R1322 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n21 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n20 3.05467
R1323 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n22 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n21 0.965083
R1324 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n24 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n22 0.646333
R1325 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n24 0.063
R1326 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n33 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t32 141.215
R1327 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t37 141.215
R1328 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t35 141.215
R1329 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t26 141.215
R1330 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n33 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t23 139.879
R1331 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n34 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t24 139.879
R1332 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n35 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t29 139.879
R1333 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n32 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t25 139.879
R1334 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n31 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t39 139.879
R1335 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n30 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t21 139.879
R1336 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t20 139.879
R1337 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t22 139.879
R1338 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t31 139.879
R1339 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t38 139.879
R1340 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t30 139.879
R1341 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t34 139.879
R1342 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t27 139.879
R1343 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t36 139.879
R1344 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t28 139.879
R1345 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t33 139.879
R1346 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t12 134.738
R1347 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t8 134.738
R1348 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t2 134.738
R1349 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t13 134.738
R1350 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t0 134.738
R1351 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t5 134.738
R1352 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t18 134.738
R1353 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t4 134.738
R1354 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t17 134.738
R1355 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t9 134.738
R1356 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t15 134.738
R1357 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t3 134.738
R1358 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t1 134.738
R1359 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t7 134.738
R1360 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t6 134.738
R1361 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t10 134.738
R1362 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t11 134.738
R1363 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t16 134.738
R1364 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t14 134.738
R1365 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t19 134.738
R1366 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n0 7.63383
R1367 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n5 7.63383
R1368 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n9 7.63383
R1369 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n12 7.63383
R1370 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n37 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n27 5.55541
R1371 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n8 4.52426
R1372 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n1 4.5005
R1373 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n3 4.5005
R1374 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n6 4.5005
R1375 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n15 4.5005
R1376 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n13 4.5005
R1377 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n10 4.5005
R1378 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n37 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n36 3.4105
R1379 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n17 3.4105
R1380 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n2 3.13383
R1381 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n14 3.13383
R1382 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n11 3.00675
R1383 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n28 1.79633
R1384 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n31 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n30 1.79633
R1385 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n34 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n33 1.79633
R1386 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n19 1.79633
R1387 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n21 1.79633
R1388 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n25 1.79633
R1389 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n23 1.79633
R1390 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n7 1.69425
R1391 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n4 1.44008
R1392 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n30 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n29 1.338
R1393 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n32 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n31 1.338
R1394 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n35 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n34 1.338
R1395 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n20 1.338
R1396 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n24 1.338
R1397 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n36 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n35 1.0255
R1398 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n26 0.796333
R1399 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n36 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n32 0.771333
R1400 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n22 0.542167
R1401 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n18 0.265409
R1402 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n16 0.127583
R1403 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n37 0.111591
R1404 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n45 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t5 85.5564
R1405 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n38 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t11 84.4381
R1406 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n35 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t14 84.4381
R1407 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n32 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t21 84.4381
R1408 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n30 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t18 84.4381
R1409 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n33 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t10 84.4381
R1410 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n36 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t26 84.4381
R1411 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n39 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t4 84.4381
R1412 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n43 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t3 84.4381
R1413 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n42 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t1 84.4381
R1414 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n31 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n2 75.1793
R1415 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n34 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n1 75.1793
R1416 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n37 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n0 75.1793
R1417 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n45 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n44 75.1793
R1418 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n41 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n40 75.1793
R1419 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n28 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t16 65.5634
R1420 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n27 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t12 65.0567
R1421 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n25 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n24 59.0738
R1422 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n26 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n22 49.2215
R1423 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n25 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n23 49.0864
R1424 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n29 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n21 24.3828
R1425 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n30 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n29 19.7755
R1426 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n27 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n26 18.5582
R1427 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n33 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n32 10.5047
R1428 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n36 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n35 10.5047
R1429 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n39 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n38 10.5047
R1430 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n43 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n42 10.5047
R1431 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n22 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t15 10.3318
R1432 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n22 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t7 10.3318
R1433 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n24 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t13 10.3318
R1434 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n24 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t19 10.3318
R1435 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t25 10.3318
R1436 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t20 10.3318
R1437 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n31 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 9.74143
R1438 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n34 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 9.74143
R1439 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n37 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 9.74143
R1440 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n41 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 9.74143
R1441 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n45 9.74061
R1442 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t17 9.23217
R1443 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t22 9.23217
R1444 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t6 9.23217
R1445 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t27 9.23217
R1446 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t24 9.23217
R1447 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t9 9.23217
R1448 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n44 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t23 9.23217
R1449 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n44 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t8 9.23217
R1450 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n40 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t2 9.23217
R1451 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n40 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t0 9.23217
R1452 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n28 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 5.863
R1453 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n27 5.72967
R1454 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n29 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n28 5.20675
R1455 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n5 3.90596
R1456 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n8 3.4105
R1457 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n12 3.4105
R1458 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n16 3.4105
R1459 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n20 3.4105
R1460 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n42 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n41 1.08427
R1461 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n26 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n25 1.00227
R1462 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n32 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n31 0.929322
R1463 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n35 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n34 0.929322
R1464 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n38 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n37 0.929322
R1465 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t31 0.523604
R1466 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t33 0.523604
R1467 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t41 0.523604
R1468 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t43 0.523604
R1469 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t34 0.523604
R1470 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t36 0.523604
R1471 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t44 0.523604
R1472 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t47 0.523604
R1473 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t37 0.523604
R1474 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t39 0.523604
R1475 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n17 0.495958
R1476 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n13 0.495958
R1477 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n9 0.495958
R1478 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t46 0.28175
R1479 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t40 0.28175
R1480 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t35 0.28175
R1481 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t29 0.28175
R1482 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t28 0.28175
R1483 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t42 0.28175
R1484 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t38 0.28175
R1485 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t32 0.28175
R1486 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t30 0.28175
R1487 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t45 0.28175
R1488 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n30 0.188
R1489 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n33 0.188
R1490 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n36 0.188
R1491 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n39 0.188
R1492 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n43 0.188
R1493 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n18 0.121427
R1494 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n19 0.121427
R1495 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n14 0.121427
R1496 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n15 0.121427
R1497 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n10 0.121427
R1498 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n11 0.121427
R1499 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n6 0.121427
R1500 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n7 0.121427
R1501 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n3 0.121427
R1502 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n4 0.121427
R1503 VOUT.n2 VOUT.n1 75.2042
R1504 VOUT.n2 VOUT.n0 75.1988
R1505 VOUT.n5 VOUT.n3 66.6872
R1506 VOUT.n5 VOUT.n4 66.6872
R1507 VOUT.n3 VOUT.t2 16.5305
R1508 VOUT.n3 VOUT.t16 16.5305
R1509 VOUT.n4 VOUT.t15 16.5305
R1510 VOUT.n4 VOUT.t42 16.5305
R1511 VOUT.n45 VOUT.n44 13.8209
R1512 VOUT.n0 VOUT.t45 9.23217
R1513 VOUT.n0 VOUT.t12 9.23217
R1514 VOUT.n1 VOUT.t0 9.23217
R1515 VOUT.n1 VOUT.t9 9.23217
R1516 VOUT VOUT.n2 8.64633
R1517 VOUT.n45 VOUT.n5 8.48696
R1518 VOUT.n12 VOUT.n8 3.90596
R1519 VOUT.n12 VOUT.n11 3.4105
R1520 VOUT.n16 VOUT.n15 3.4105
R1521 VOUT.n20 VOUT.n19 3.4105
R1522 VOUT.n24 VOUT.n23 3.4105
R1523 VOUT.n28 VOUT.n27 3.4105
R1524 VOUT.n32 VOUT.n31 3.4105
R1525 VOUT.n36 VOUT.n35 3.4105
R1526 VOUT.n40 VOUT.n39 3.4105
R1527 VOUT.n44 VOUT.n43 3.4105
R1528 VOUT.n41 VOUT.t47 1.082
R1529 VOUT.n37 VOUT.t6 1.082
R1530 VOUT.n33 VOUT.t46 1.082
R1531 VOUT.n29 VOUT.t7 1.082
R1532 VOUT.n25 VOUT.t19 1.082
R1533 VOUT.n21 VOUT.t37 1.082
R1534 VOUT.n17 VOUT.t27 1.082
R1535 VOUT.n13 VOUT.t34 1.082
R1536 VOUT.n9 VOUT.t24 1.082
R1537 VOUT.n6 VOUT.t31 1.082
R1538 VOUT.n28 VOUT.n24 0.991417
R1539 VOUT.n43 VOUT.t14 0.90575
R1540 VOUT.n39 VOUT.t41 0.90575
R1541 VOUT.n35 VOUT.t17 0.90575
R1542 VOUT.n31 VOUT.t5 0.90575
R1543 VOUT.n27 VOUT.t10 0.90575
R1544 VOUT.n23 VOUT.t35 0.90575
R1545 VOUT.n19 VOUT.t25 0.90575
R1546 VOUT.n15 VOUT.t32 0.90575
R1547 VOUT.n11 VOUT.t21 0.90575
R1548 VOUT.n8 VOUT.t29 0.90575
R1549 VOUT.n41 VOUT.t3 0.7295
R1550 VOUT.n42 VOUT.t44 0.7295
R1551 VOUT.n37 VOUT.t11 0.7295
R1552 VOUT.n38 VOUT.t8 0.7295
R1553 VOUT.n33 VOUT.t1 0.7295
R1554 VOUT.n34 VOUT.t43 0.7295
R1555 VOUT.n29 VOUT.t4 0.7295
R1556 VOUT.n30 VOUT.t18 0.7295
R1557 VOUT.n25 VOUT.t13 0.7295
R1558 VOUT.n26 VOUT.t20 0.7295
R1559 VOUT.n21 VOUT.t22 0.7295
R1560 VOUT.n22 VOUT.t28 0.7295
R1561 VOUT.n17 VOUT.t33 0.7295
R1562 VOUT.n18 VOUT.t39 0.7295
R1563 VOUT.n13 VOUT.t40 0.7295
R1564 VOUT.n14 VOUT.t26 0.7295
R1565 VOUT.n9 VOUT.t30 0.7295
R1566 VOUT.n10 VOUT.t36 0.7295
R1567 VOUT.n6 VOUT.t38 0.7295
R1568 VOUT.n7 VOUT.t23 0.7295
R1569 VOUT.n44 VOUT.n40 0.495958
R1570 VOUT.n40 VOUT.n36 0.495958
R1571 VOUT.n36 VOUT.n32 0.495958
R1572 VOUT.n32 VOUT.n28 0.495958
R1573 VOUT.n24 VOUT.n20 0.495958
R1574 VOUT.n20 VOUT.n16 0.495958
R1575 VOUT.n16 VOUT.n12 0.495958
R1576 VOUT.n42 VOUT.n41 0.353
R1577 VOUT.n38 VOUT.n37 0.353
R1578 VOUT.n34 VOUT.n33 0.353
R1579 VOUT.n30 VOUT.n29 0.353
R1580 VOUT.n26 VOUT.n25 0.353
R1581 VOUT.n22 VOUT.n21 0.353
R1582 VOUT.n18 VOUT.n17 0.353
R1583 VOUT.n14 VOUT.n13 0.353
R1584 VOUT.n10 VOUT.n9 0.353
R1585 VOUT.n7 VOUT.n6 0.353
R1586 VOUT.n43 VOUT.n42 0.17675
R1587 VOUT.n39 VOUT.n38 0.17675
R1588 VOUT.n35 VOUT.n34 0.17675
R1589 VOUT.n31 VOUT.n30 0.17675
R1590 VOUT.n27 VOUT.n26 0.17675
R1591 VOUT.n23 VOUT.n22 0.17675
R1592 VOUT.n19 VOUT.n18 0.17675
R1593 VOUT.n15 VOUT.n14 0.17675
R1594 VOUT.n11 VOUT.n10 0.17675
R1595 VOUT.n8 VOUT.n7 0.17675
R1596 VOUT VOUT.n45 0.0838333
R1597 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n32 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t30 141.399
R1598 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t22 141.399
R1599 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t23 141.399
R1600 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t31 141.399
R1601 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n32 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t27 140.061
R1602 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n33 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t20 140.061
R1603 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n34 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t26 140.061
R1604 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n35 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t29 140.061
R1605 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n31 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t24 140.061
R1606 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n30 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t38 140.061
R1607 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t25 140.061
R1608 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t28 140.061
R1609 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t36 140.061
R1610 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t37 140.061
R1611 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t21 140.061
R1612 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t39 140.061
R1613 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t32 140.061
R1614 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t34 140.061
R1615 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t33 140.061
R1616 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t35 140.061
R1617 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t9 134.738
R1618 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t17 134.738
R1619 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t3 134.738
R1620 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t4 134.738
R1621 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t15 134.738
R1622 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t6 134.738
R1623 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t1 134.738
R1624 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t16 134.738
R1625 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t2 134.738
R1626 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t0 134.738
R1627 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t12 134.738
R1628 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t13 134.738
R1629 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t18 134.738
R1630 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t14 134.738
R1631 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t7 134.738
R1632 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t10 134.738
R1633 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t8 134.738
R1634 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t11 134.738
R1635 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t5 134.738
R1636 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t19 134.738
R1637 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n9 7.63383
R1638 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n14 7.63383
R1639 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n0 7.63383
R1640 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n3 7.63383
R1641 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n37 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n27 5.68074
R1642 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n8 4.64959
R1643 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n10 4.5005
R1644 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n12 4.5005
R1645 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n15 4.5005
R1646 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n1 4.5005
R1647 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n4 4.5005
R1648 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n6 4.5005
R1649 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n37 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n36 3.4105
R1650 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n17 3.4105
R1651 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n11 3.13383
R1652 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n5 3.13383
R1653 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n2 2.74425
R1654 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n16 1.95675
R1655 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n28 1.79633
R1656 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n31 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n30 1.79633
R1657 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n35 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n34 1.79633
R1658 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n33 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n32 1.79633
R1659 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n19 1.79633
R1660 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n21 1.79633
R1661 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n24 1.79633
R1662 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n30 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n29 1.338
R1663 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n34 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n33 1.338
R1664 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n20 1.338
R1665 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n22 1.338
R1666 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n25 1.338
R1667 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n26 1.288
R1668 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n13 1.17758
R1669 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n36 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n35 1.05883
R1670 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n23 0.508833
R1671 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n7 0.390083
R1672 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n36 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n31 0.279667
R1673 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n18 0.202742
R1674 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n37 0.0489242
R1675 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n68 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n67 194.3
R1676 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n0 194.3
R1677 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n19 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t9 135.499
R1678 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n20 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t15 135.499
R1679 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n19 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t8 134.715
R1680 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n20 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t41 134.715
R1681 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n8 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t24 111.398
R1682 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n4 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t4 111.398
R1683 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n26 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t60 111.398
R1684 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n40 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t20 111.398
R1685 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n37 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t63 111.398
R1686 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n55 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t12 111.398
R1687 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n51 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t5 111.398
R1688 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n8 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t46 110.615
R1689 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n9 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t6 110.615
R1690 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n10 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t47 110.615
R1691 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n11 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t26 110.615
R1692 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n12 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t58 110.615
R1693 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n13 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t25 110.615
R1694 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n14 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t45 110.615
R1695 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n15 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t39 110.615
R1696 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n16 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t62 110.615
R1697 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n17 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t29 110.615
R1698 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n7 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t66 110.615
R1699 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n6 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t40 110.615
R1700 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n5 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t19 110.615
R1701 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n4 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t43 110.615
R1702 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n26 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t23 110.615
R1703 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n27 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t61 110.615
R1704 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n28 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t36 110.615
R1705 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n29 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t11 110.615
R1706 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n30 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t35 110.615
R1707 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n31 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t57 110.615
R1708 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n32 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t48 110.615
R1709 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n33 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t13 110.615
R1710 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n34 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t38 110.615
R1711 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n25 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t16 110.615
R1712 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n24 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t51 110.615
R1713 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n23 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t34 110.615
R1714 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n22 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t52 110.615
R1715 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n40 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t53 110.615
R1716 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n41 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t54 110.615
R1717 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n42 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t18 110.615
R1718 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n43 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t22 110.615
R1719 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n44 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t44 110.615
R1720 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n45 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t17 110.615
R1721 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n46 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t67 110.615
R1722 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n47 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t42 110.615
R1723 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n48 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t64 110.615
R1724 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n39 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t65 110.615
R1725 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n38 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t28 110.615
R1726 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n37 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t30 110.615
R1727 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n55 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t50 110.615
R1728 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n56 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t21 110.615
R1729 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n57 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t7 110.615
R1730 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n58 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t49 110.615
R1731 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n59 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t14 110.615
R1732 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n60 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t56 110.615
R1733 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n61 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t27 110.615
R1734 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n62 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t33 110.615
R1735 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n63 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t55 110.615
R1736 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n64 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t37 110.615
R1737 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n54 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t32 110.615
R1738 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n53 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t10 110.615
R1739 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n52 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t59 110.615
R1740 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n51 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t31 110.615
R1741 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n67 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t3 27.5505
R1742 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n67 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t1 27.5505
R1743 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n0 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t0 27.5505
R1744 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n0 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t2 27.5505
R1745 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n22 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n21 13.3067
R1746 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n20 6.23592
R1747 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n21 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n19 5.8755
R1748 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n69 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n68 5.04842
R1749 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n3 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n1 5.04842
R1750 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n68 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n2 5.04633
R1751 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n73 4.98383
R1752 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n36 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n18 3.84917
R1753 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n72 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n71 3.62129
R1754 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n71 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n70 3.4105
R1755 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n66 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n65 3.4105
R1756 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n50 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n49 3.4105
R1757 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n36 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n35 3.4105
R1758 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n71 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n66 1.97948
R1759 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n21 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.860917
R1760 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n5 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n4 0.783833
R1761 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n6 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n5 0.783833
R1762 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n7 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n6 0.783833
R1763 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n17 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n16 0.783833
R1764 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n16 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n15 0.783833
R1765 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n15 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n14 0.783833
R1766 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n14 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n13 0.783833
R1767 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n13 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n12 0.783833
R1768 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n12 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n11 0.783833
R1769 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n11 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n10 0.783833
R1770 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n10 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n9 0.783833
R1771 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n9 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n8 0.783833
R1772 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n23 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n22 0.783833
R1773 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n24 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n23 0.783833
R1774 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n25 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n24 0.783833
R1775 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n34 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n33 0.783833
R1776 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n33 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n32 0.783833
R1777 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n32 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n31 0.783833
R1778 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n31 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n30 0.783833
R1779 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n30 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n29 0.783833
R1780 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n29 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n28 0.783833
R1781 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n28 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n27 0.783833
R1782 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n27 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n26 0.783833
R1783 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n38 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n37 0.783833
R1784 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n39 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n38 0.783833
R1785 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n48 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n47 0.783833
R1786 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n47 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n46 0.783833
R1787 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n46 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n45 0.783833
R1788 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n45 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n44 0.783833
R1789 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n44 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n43 0.783833
R1790 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n43 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n42 0.783833
R1791 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n42 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n41 0.783833
R1792 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n41 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n40 0.783833
R1793 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n52 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n51 0.783833
R1794 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n53 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n52 0.783833
R1795 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n54 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n53 0.783833
R1796 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n64 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n63 0.783833
R1797 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n63 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n62 0.783833
R1798 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n62 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n61 0.783833
R1799 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n61 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n60 0.783833
R1800 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n60 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n59 0.783833
R1801 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n59 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n58 0.783833
R1802 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n58 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n57 0.783833
R1803 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n57 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n56 0.783833
R1804 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n56 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n55 0.783833
R1805 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n50 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n36 0.642121
R1806 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n70 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n69 0.548417
R1807 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n72 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n3 0.548417
R1808 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n70 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n2 0.546333
R1809 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n73 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n72 0.546333
R1810 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n69 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n3 0.492167
R1811 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n73 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n2 0.492167
R1812 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n66 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n50 0.439167
R1813 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n18 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n17 0.413
R1814 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n35 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n34 0.413
R1815 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n49 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n48 0.413
R1816 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n65 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n64 0.413
R1817 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n18 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n7 0.371333
R1818 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n35 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n25 0.371333
R1819 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n49 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n39 0.371333
R1820 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n65 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n54 0.371333
R1821 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n1 0.063
R1822 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n36 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t20 238.911
R1823 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n36 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t21 222.089
R1824 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t13 221.974
R1825 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t2 221.974
R1826 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t6 221.913
R1827 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t5 221.913
R1828 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t8 221.913
R1829 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t9 221.913
R1830 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t7 221.911
R1831 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t1 221.911
R1832 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t19 221.851
R1833 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t11 221.851
R1834 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t18 221.851
R1835 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t3 221.851
R1836 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t12 221.851
R1837 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t17 221.851
R1838 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t14 221.851
R1839 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t16 221.851
R1840 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t4 221.851
R1841 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t15 221.851
R1842 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t10 221.851
R1843 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t0 221.851
R1844 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n45 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t74 111.398
R1845 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t72 111.398
R1846 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n70 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t53 111.398
R1847 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n38 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t69 111.398
R1848 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n53 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t81 110.615
R1849 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n54 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t59 110.615
R1850 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n55 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t27 110.615
R1851 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n56 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t76 110.615
R1852 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n57 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t58 110.615
R1853 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n58 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t23 110.615
R1854 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n59 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t65 110.615
R1855 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n52 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t31 110.615
R1856 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n51 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t40 110.615
R1857 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n50 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t64 110.615
R1858 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n49 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t47 110.615
R1859 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n48 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t36 110.615
R1860 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n47 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t78 110.615
R1861 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n46 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t68 110.615
R1862 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n45 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t35 110.615
R1863 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n85 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t79 110.615
R1864 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n86 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t57 110.615
R1865 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n87 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t26 110.615
R1866 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n88 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t75 110.615
R1867 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n89 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t56 110.615
R1868 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n90 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t22 110.615
R1869 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n91 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t63 110.615
R1870 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n35 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t30 110.615
R1871 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n34 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t39 110.615
R1872 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n33 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t62 110.615
R1873 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n32 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t46 110.615
R1874 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n31 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t34 110.615
R1875 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n30 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t77 110.615
R1876 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t67 110.615
R1877 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t33 110.615
R1878 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n83 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t25 110.615
R1879 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n82 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t50 110.615
R1880 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n81 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t43 110.615
R1881 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n80 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t24 110.615
R1882 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n79 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t48 110.615
R1883 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n78 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t29 110.615
R1884 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n76 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t52 110.615
R1885 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n75 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t61 110.615
R1886 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n74 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t28 110.615
R1887 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n73 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t71 110.615
R1888 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n72 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t54 110.615
R1889 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n71 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t45 110.615
R1890 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n70 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t32 110.615
R1891 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n68 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t38 110.615
R1892 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n67 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t60 110.615
R1893 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n66 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t49 110.615
R1894 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n65 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t37 110.615
R1895 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n64 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t55 110.615
R1896 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n63 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t42 110.615
R1897 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n44 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t66 110.615
R1898 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n43 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t73 110.615
R1899 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n42 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t41 110.615
R1900 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n41 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t80 110.615
R1901 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n40 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t70 110.615
R1902 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n39 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t51 110.615
R1903 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n38 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t44 110.615
R1904 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n37 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 8.31322
R1905 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n2 5.697
R1906 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n13 5.697
R1907 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n20 5.697
R1908 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n11 5.6845
R1909 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n21 5.55802
R1910 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n14 5.55802
R1911 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n16 5.55802
R1912 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n9 5.55802
R1913 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n7 5.55802
R1914 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n5 5.55802
R1915 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n3 5.55802
R1916 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n23 5.55802
R1917 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n12 5.43008
R1918 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n84 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n83 5.35189
R1919 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n69 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n68 5.35189
R1920 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n85 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n84 4.88189
R1921 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n53 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n37 4.56856
R1922 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n61 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n60 3.72383
R1923 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n62 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n61 3.4105
R1924 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n77 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n27 3.4105
R1925 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n93 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n92 3.4105
R1926 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n25 3.4105
R1927 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n6 2.888
R1928 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n17 1.57967
R1929 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n36 1.30883
R1930 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n24 1.30883
R1931 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n18 1.07342
R1932 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n0 1.07342
R1933 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n28 0.783833
R1934 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n30 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n29 0.783833
R1935 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n31 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n30 0.783833
R1936 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n32 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n31 0.783833
R1937 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n33 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n32 0.783833
R1938 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n34 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n33 0.783833
R1939 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n35 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n34 0.783833
R1940 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n91 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n90 0.783833
R1941 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n90 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n89 0.783833
R1942 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n89 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n88 0.783833
R1943 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n88 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n87 0.783833
R1944 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n87 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n86 0.783833
R1945 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n86 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n85 0.783833
R1946 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n71 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n70 0.783833
R1947 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n72 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n71 0.783833
R1948 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n73 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n72 0.783833
R1949 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n74 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n73 0.783833
R1950 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n75 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n74 0.783833
R1951 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n76 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n75 0.783833
R1952 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n79 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n78 0.783833
R1953 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n80 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n79 0.783833
R1954 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n81 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n80 0.783833
R1955 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n82 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n81 0.783833
R1956 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n83 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n82 0.783833
R1957 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n39 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n38 0.783833
R1958 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n40 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n39 0.783833
R1959 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n41 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n40 0.783833
R1960 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n42 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n41 0.783833
R1961 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n43 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n42 0.783833
R1962 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n44 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n43 0.783833
R1963 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n64 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n63 0.783833
R1964 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n65 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n64 0.783833
R1965 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n66 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n65 0.783833
R1966 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n67 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n66 0.783833
R1967 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n68 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n67 0.783833
R1968 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n46 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n45 0.783833
R1969 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n47 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n46 0.783833
R1970 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n48 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n47 0.783833
R1971 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n49 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n48 0.783833
R1972 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n50 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n49 0.783833
R1973 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n51 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n50 0.783833
R1974 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n52 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n51 0.783833
R1975 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n59 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n58 0.783833
R1976 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n58 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n57 0.783833
R1977 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n57 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n56 0.783833
R1978 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n56 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n55 0.783833
R1979 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n55 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n54 0.783833
R1980 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n54 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n53 0.783833
R1981 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n92 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n35 0.527583
R1982 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n77 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n76 0.527583
R1983 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n62 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n44 0.527583
R1984 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n60 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n52 0.527583
R1985 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n84 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n69 0.390742
R1986 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n61 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n27 0.390742
R1987 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n69 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n37 0.313833
R1988 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n93 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n27 0.313833
R1989 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n92 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n91 0.25675
R1990 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n78 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n77 0.25675
R1991 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n63 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n62 0.25675
R1992 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n60 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n59 0.25675
R1993 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n3 0.246333
R1994 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n7 0.246333
R1995 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n14 0.246333
R1996 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n21 0.246333
R1997 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n93 0.174258
R1998 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n15 0.123417
R1999 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n8 0.123417
R2000 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n4 0.123417
R2001 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n22 0.123417
R2002 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n26 0.0916515
R2003 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n19 0.0604849
R2004 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n1 0.0604849
R2005 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n10 0.013
R2006 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t18 228.413
R2007 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t16 228.413
R2008 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t1 228.413
R2009 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t19 228.413
R2010 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t7 227.093
R2011 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t13 227.093
R2012 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t8 227.093
R2013 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t12 227.093
R2014 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t0 227.093
R2015 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t6 227.093
R2016 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t15 227.093
R2017 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t11 227.093
R2018 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t2 227.093
R2019 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t17 227.093
R2020 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t4 224.073
R2021 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t14 224.073
R2022 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t28 221.974
R2023 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t21 221.974
R2024 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n33 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t35 221.911
R2025 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n33 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t34 221.911
R2026 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n34 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t38 221.911
R2027 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n34 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t30 221.911
R2028 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n31 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t29 221.911
R2029 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n31 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t26 221.911
R2030 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n30 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t33 221.911
R2031 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t36 221.911
R2032 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t23 221.911
R2033 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t37 221.911
R2034 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t24 221.911
R2035 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t39 221.911
R2036 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t32 221.911
R2037 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t31 221.911
R2038 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t9 221.851
R2039 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t10 221.851
R2040 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t5 221.851
R2041 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t3 221.851
R2042 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t27 221.851
R2043 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t20 221.851
R2044 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t22 221.851
R2045 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t25 221.851
R2046 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n35 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n33 7.90675
R2047 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n32 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n30 7.90675
R2048 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n24 7.90675
R2049 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n19 7.90675
R2050 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n1 5.2428
R2051 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n13 5.2428
R2052 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n8 5.17941
R2053 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n35 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n34 4.77342
R2054 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n32 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n31 4.77342
R2055 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n25 4.77342
R2056 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n20 4.77342
R2057 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n37 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n27 4.55274
R2058 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n37 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n36 3.4105
R2059 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n17 3.4105
R2060 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n36 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n32 3.00675
R2061 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n9 1.813
R2062 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n14 1.813
R2063 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n2 1.813
R2064 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n4 1.813
R2065 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n6 1.813
R2066 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n0 1.70775
R2067 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n12 1.70775
R2068 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n26 1.69425
R2069 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n28 1.65556
R2070 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n22 1.65556
R2071 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n21 1.44008
R2072 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n10 1.32133
R2073 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n15 1.32133
R2074 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n3 1.32133
R2075 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n16 1.03383
R2076 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n7 0.788
R2077 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n11 0.779667
R2078 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n5 0.533833
R2079 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n18 0.216985
R2080 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n36 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n35 0.127583
R2081 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n37 0.111591
R2082 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n30 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n29 0.0619583
R2083 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n23 0.0619583
R2084 GNDA.t82 GNDA.n215 229046
R2085 GNDA.n441 GNDA.n7 15808.4
R2086 GNDA.n441 GNDA.n8 15808.4
R2087 GNDA.n147 GNDA.n7 15805.2
R2088 GNDA.n147 GNDA.n8 15805.2
R2089 GNDA.n367 GNDA.n172 13405
R2090 GNDA.n367 GNDA.n146 13405
R2091 GNDA.n149 GNDA.n95 12564.6
R2092 GNDA.n196 GNDA.n95 12564.6
R2093 GNDA.n193 GNDA.n168 11046.2
R2094 GNDA.n168 GNDA.n144 11046.2
R2095 GNDA.n299 GNDA.n171 11046.2
R2096 GNDA.n171 GNDA.n145 11046.2
R2097 GNDA.n300 GNDA.n137 11046.2
R2098 GNDA.n148 GNDA.n137 11046.2
R2099 GNDA.n276 GNDA.n203 5956.02
R2100 GNDA.n219 GNDA.n203 5956.02
R2101 GNDA.n227 GNDA.n223 4724.07
R2102 GNDA.n223 GNDA.n214 4724.07
R2103 GNDA.n281 GNDA.n280 4431.2
R2104 GNDA.n280 GNDA.n201 4431.2
R2105 GNDA.n383 GNDA.n150 4431.2
R2106 GNDA.n383 GNDA.n151 4431.2
R2107 GNDA.n276 GNDA.n202 3513.17
R2108 GNDA.n220 GNDA.n219 3513.17
R2109 GNDA.n336 GNDA.n191 2982.78
R2110 GNDA.n338 GNDA.n191 2982.78
R2111 GNDA.n338 GNDA.n190 2982.78
R2112 GNDA.n336 GNDA.n190 2982.78
R2113 GNDA.n281 GNDA.n197 2750.4
R2114 GNDA.n291 GNDA.n197 2750.4
R2115 GNDA.n291 GNDA.n166 2750.4
R2116 GNDA.n370 GNDA.n166 2750.4
R2117 GNDA.n370 GNDA.n159 2750.4
R2118 GNDA.n375 GNDA.n159 2750.4
R2119 GNDA.n375 GNDA.n163 2750.4
R2120 GNDA.n163 GNDA.n150 2750.4
R2121 GNDA.n201 GNDA.n198 2750.4
R2122 GNDA.n293 GNDA.n198 2750.4
R2123 GNDA.n293 GNDA.n285 2750.4
R2124 GNDA.n285 GNDA.n167 2750.4
R2125 GNDA.n167 GNDA.n157 2750.4
R2126 GNDA.n377 GNDA.n157 2750.4
R2127 GNDA.n377 GNDA.n158 2750.4
R2128 GNDA.n158 GNDA.n151 2750.4
R2129 GNDA.t116 GNDA.n215 2601.35
R2130 GNDA.n445 GNDA.n4 2533.93
R2131 GNDA.n445 GNDA.n5 2533.93
R2132 GNDA.n252 GNDA.n5 2533.93
R2133 GNDA.n252 GNDA.n4 2533.93
R2134 GNDA.n232 GNDA.n218 2384.32
R2135 GNDA.n232 GNDA.n231 2384.32
R2136 GNDA.n250 GNDA.n218 2339.75
R2137 GNDA.n250 GNDA.n220 2339.75
R2138 GNDA.n231 GNDA.n227 2339.75
R2139 GNDA.n231 GNDA.n230 2339.75
R2140 GNDA.n230 GNDA.n202 2339.75
R2141 GNDA.n218 GNDA.n214 2339.75
R2142 GNDA.n385 GNDA.n144 2317.47
R2143 GNDA.n385 GNDA.n145 2317.47
R2144 GNDA.n194 GNDA.n193 2317.47
R2145 GNDA.n299 GNDA.n194 2317.47
R2146 GNDA.n193 GNDA.n172 2276.08
R2147 GNDA.n146 GNDA.n144 2276.08
R2148 GNDA.t82 GNDA.n216 1917.57
R2149 GNDA.t116 GNDA.n216 1917.57
R2150 GNDA.n440 GNDA.n9 1874.45
R2151 GNDA.n11 GNDA.n9 1874.07
R2152 GNDA.n439 GNDA.n11 1874.07
R2153 GNDA GNDA.n439 1728.75
R2154 GNDA.n163 GNDA.n162 1680.8
R2155 GNDA.n162 GNDA.n158 1680.8
R2156 GNDA.n169 GNDA.n159 1680.8
R2157 GNDA.n169 GNDA.n157 1680.8
R2158 GNDA.n288 GNDA.n166 1680.8
R2159 GNDA.n288 GNDA.n285 1680.8
R2160 GNDA.n297 GNDA.n197 1680.8
R2161 GNDA.n297 GNDA.n198 1680.8
R2162 GNDA.n431 GNDA.n430 1485.93
R2163 GNDA.n430 GNDA.n94 1485.93
R2164 GNDA.n329 GNDA.n299 1477.07
R2165 GNDA.n329 GNDA.n300 1477.07
R2166 GNDA.n145 GNDA.n139 1477.07
R2167 GNDA.n148 GNDA.n139 1477.07
R2168 GNDA.n149 GNDA.n148 1435.68
R2169 GNDA.n300 GNDA.n196 1435.68
R2170 GNDA.n392 GNDA.n136 1306.35
R2171 GNDA.n392 GNDA.n391 1306.35
R2172 GNDA.n355 GNDA.n354 1306.35
R2173 GNDA.n354 GNDA.n143 1306.35
R2174 GNDA.n327 GNDA.n326 1306.35
R2175 GNDA.n326 GNDA.n138 1306.35
R2176 GNDA.n331 GNDA.t198 1215.45
R2177 GNDA.n443 GNDA.n442 1003.15
R2178 GNDA.n235 GNDA.n220 922.962
R2179 GNDA.n235 GNDA.n202 922.962
R2180 GNDA.n275 GNDA.n274 709.271
R2181 GNDA.n274 GNDA.n206 709.271
R2182 GNDA.n279 GNDA.n277 655.385
R2183 GNDA.n200 GNDA.n199 528.942
R2184 GNDA.n282 GNDA.n199 528.942
R2185 GNDA.n382 GNDA.n152 528.942
R2186 GNDA.n226 GNDA.n225 521.788
R2187 GNDA.n331 GNDA.t118 445.034
R2188 GNDA.n275 GNDA.n204 422.582
R2189 GNDA.n248 GNDA.n206 422.582
R2190 GNDA.n279 GNDA.n278 399.562
R2191 GNDA.t110 GNDA.t100 363.033
R2192 GNDA.t94 GNDA.t98 358.81
R2193 GNDA.n335 GNDA.n189 357.647
R2194 GNDA.n339 GNDA.n189 357.647
R2195 GNDA.n339 GNDA.n188 357.647
R2196 GNDA.n335 GNDA.n188 357.647
R2197 GNDA.n219 GNDA.t285 353.01
R2198 GNDA.n283 GNDA.n282 325.272
R2199 GNDA.n290 GNDA.n283 325.272
R2200 GNDA.n290 GNDA.n165 325.272
R2201 GNDA.n371 GNDA.n165 325.272
R2202 GNDA.n372 GNDA.n371 325.272
R2203 GNDA.n374 GNDA.n372 325.272
R2204 GNDA.n374 GNDA.n373 325.272
R2205 GNDA.n373 GNDA.n152 325.272
R2206 GNDA.n277 GNDA.t234 316.447
R2207 GNDA.n200 GNDA.n176 309.8
R2208 GNDA.n446 GNDA.n2 304.565
R2209 GNDA.n253 GNDA.n2 304.565
R2210 GNDA.n224 GNDA.n213 281.976
R2211 GNDA.n234 GNDA.n233 281.976
R2212 GNDA.n233 GNDA.n222 281.976
R2213 GNDA.n226 GNDA.n222 281.601
R2214 GNDA.n221 GNDA.n213 281.601
R2215 GNDA.n234 GNDA.n221 281.601
R2216 GNDA.n249 GNDA.n234 281.601
R2217 GNDA.n249 GNDA.n248 281.601
R2218 GNDA.n228 GNDA.n222 281.601
R2219 GNDA.n228 GNDA.n204 281.601
R2220 GNDA.n381 GNDA.n154 278.966
R2221 GNDA.n357 GNDA.n176 278.966
R2222 GNDA.n355 GNDA.n177 278.966
R2223 GNDA.n327 GNDA.n177 278.966
R2224 GNDA.n386 GNDA.n143 278.966
R2225 GNDA.n386 GNDA.n138 278.966
R2226 GNDA.n153 GNDA.n143 274.072
R2227 GNDA.n356 GNDA.n355 274.072
R2228 GNDA.n126 GNDA.t226 222.456
R2229 GNDA.n404 GNDA.t260 222.456
R2230 GNDA.n348 GNDA.t283 222.456
R2231 GNDA.n344 GNDA.t189 222.456
R2232 GNDA.n183 GNDA.t238 222.456
R2233 GNDA.n179 GNDA.t146 222.456
R2234 GNDA.n401 GNDA.t290 222.456
R2235 GNDA.n121 GNDA.t252 222.456
R2236 GNDA.n100 GNDA.t180 222.452
R2237 GNDA.n422 GNDA.t157 222.452
R2238 GNDA.n304 GNDA.t167 222.452
R2239 GNDA.n349 GNDA.t130 222.452
R2240 GNDA.n345 GNDA.t202 222.452
R2241 GNDA.n182 GNDA.t246 222.452
R2242 GNDA.n178 GNDA.t258 222.452
R2243 GNDA.n315 GNDA.t183 222.452
R2244 GNDA.n90 GNDA.t150 222.379
R2245 GNDA.n103 GNDA.t200 222.379
R2246 GNDA.n91 GNDA.t151 222.355
R2247 GNDA.n104 GNDA.t199 222.355
R2248 GNDA.n89 GNDA.t276 222.297
R2249 GNDA.n437 GNDA.t207 222.297
R2250 GNDA.n87 GNDA.t275 222.263
R2251 GNDA.n435 GNDA.t208 222.263
R2252 GNDA.n140 GNDA.t296 222.228
R2253 GNDA.n140 GNDA.t295 222.228
R2254 GNDA.n360 GNDA.t172 222.228
R2255 GNDA.n360 GNDA.t171 222.228
R2256 GNDA.n362 GNDA.t229 222.228
R2257 GNDA.n362 GNDA.t228 222.228
R2258 GNDA.n318 GNDA.t160 222.228
R2259 GNDA.n318 GNDA.t159 222.228
R2260 GNDA.n96 GNDA.t68 221.851
R2261 GNDA.n96 GNDA.t59 221.851
R2262 GNDA.n101 GNDA.t25 221.851
R2263 GNDA.n101 GNDA.t181 221.851
R2264 GNDA.n99 GNDA.t31 221.851
R2265 GNDA.n99 GNDA.t64 221.851
R2266 GNDA.n98 GNDA.t63 221.851
R2267 GNDA.n98 GNDA.t21 221.851
R2268 GNDA.n97 GNDA.t36 221.851
R2269 GNDA.n97 GNDA.t52 221.851
R2270 GNDA.n419 GNDA.t76 221.851
R2271 GNDA.n419 GNDA.t35 221.851
R2272 GNDA.n420 GNDA.t23 221.851
R2273 GNDA.n420 GNDA.t41 221.851
R2274 GNDA.n421 GNDA.t40 221.851
R2275 GNDA.n421 GNDA.t73 221.851
R2276 GNDA.n423 GNDA.t156 221.851
R2277 GNDA.n423 GNDA.t18 221.851
R2278 GNDA.n122 GNDA.t251 221.851
R2279 GNDA.n122 GNDA.t232 221.851
R2280 GNDA.n127 GNDA.t225 221.851
R2281 GNDA.n127 GNDA.t192 221.851
R2282 GNDA.n120 GNDA.t231 221.851
R2283 GNDA.n120 GNDA.t70 221.851
R2284 GNDA.n130 GNDA.t191 221.851
R2285 GNDA.n130 GNDA.t61 221.851
R2286 GNDA.n398 GNDA.t46 221.851
R2287 GNDA.n398 GNDA.t249 221.851
R2288 GNDA.n406 GNDA.t30 221.851
R2289 GNDA.n406 GNDA.t215 221.851
R2290 GNDA.n402 GNDA.t248 221.851
R2291 GNDA.n402 GNDA.t291 221.851
R2292 GNDA.n405 GNDA.t214 221.851
R2293 GNDA.n405 GNDA.t261 221.851
R2294 GNDA.n301 GNDA.t77 221.851
R2295 GNDA.n301 GNDA.t38 221.851
R2296 GNDA.n302 GNDA.t24 221.851
R2297 GNDA.n302 GNDA.t43 221.851
R2298 GNDA.n303 GNDA.t42 221.851
R2299 GNDA.n303 GNDA.t74 221.851
R2300 GNDA.n305 GNDA.t166 221.851
R2301 GNDA.n305 GNDA.t20 221.851
R2302 GNDA.n346 GNDA.t188 221.851
R2303 GNDA.n346 GNDA.t203 221.851
R2304 GNDA.n350 GNDA.t282 221.851
R2305 GNDA.n350 GNDA.t131 221.851
R2306 GNDA.n180 GNDA.t257 221.851
R2307 GNDA.n180 GNDA.t147 221.851
R2308 GNDA.n184 GNDA.t245 221.851
R2309 GNDA.n184 GNDA.t239 221.851
R2310 GNDA.n311 GNDA.t69 221.851
R2311 GNDA.n311 GNDA.t60 221.851
R2312 GNDA.n312 GNDA.t37 221.851
R2313 GNDA.n312 GNDA.t53 221.851
R2314 GNDA.n313 GNDA.t65 221.851
R2315 GNDA.n313 GNDA.t22 221.851
R2316 GNDA.n314 GNDA.t32 221.851
R2317 GNDA.n314 GNDA.t66 221.851
R2318 GNDA.n316 GNDA.t27 221.851
R2319 GNDA.n316 GNDA.t184 221.851
R2320 GNDA.n107 GNDA.t54 221.851
R2321 GNDA.n107 GNDA.t67 221.851
R2322 GNDA.n108 GNDA.t48 221.851
R2323 GNDA.n108 GNDA.t55 221.851
R2324 GNDA.n109 GNDA.t28 221.851
R2325 GNDA.n109 GNDA.t45 221.851
R2326 GNDA.n110 GNDA.t19 221.851
R2327 GNDA.n110 GNDA.t29 221.851
R2328 GNDA.n111 GNDA.t33 221.851
R2329 GNDA.n111 GNDA.t72 221.851
R2330 GNDA.n112 GNDA.t26 221.851
R2331 GNDA.n112 GNDA.t58 221.851
R2332 GNDA.n113 GNDA.t71 221.851
R2333 GNDA.n113 GNDA.t47 221.851
R2334 GNDA.n114 GNDA.t57 221.851
R2335 GNDA.n114 GNDA.t34 221.851
R2336 GNDA.n115 GNDA.t75 221.851
R2337 GNDA.n115 GNDA.t51 221.851
R2338 GNDA.n116 GNDA.t62 221.851
R2339 GNDA.n116 GNDA.t44 221.851
R2340 GNDA.n117 GNDA.t49 221.851
R2341 GNDA.n117 GNDA.t56 221.851
R2342 GNDA.n118 GNDA.t39 221.851
R2343 GNDA.n118 GNDA.t50 221.851
R2344 GNDA.n442 GNDA.t198 221.787
R2345 GNDA.n373 GNDA.n155 203.672
R2346 GNDA.n379 GNDA.n155 203.672
R2347 GNDA.n372 GNDA.n164 203.672
R2348 GNDA.n164 GNDA.n156 203.672
R2349 GNDA.n287 GNDA.n165 203.672
R2350 GNDA.n287 GNDA.n284 203.672
R2351 GNDA.n296 GNDA.n283 203.672
R2352 GNDA.n296 GNDA.n295 203.672
R2353 GNDA.n382 GNDA.n381 203.672
R2354 GNDA.t89 GNDA.t102 200.107
R2355 GNDA.n328 GNDA.n327 179.577
R2356 GNDA.n328 GNDA.n136 179.577
R2357 GNDA.n390 GNDA.n138 179.577
R2358 GNDA.n391 GNDA.n390 179.577
R2359 GNDA.t96 GNDA.n192 177.296
R2360 GNDA.n337 GNDA.t81 177.296
R2361 GNDA.n391 GNDA.n93 174.683
R2362 GNDA.n195 GNDA.n136 174.683
R2363 GNDA.n255 GNDA.n254 161.882
R2364 GNDA.n255 GNDA.n3 161.882
R2365 GNDA.t106 GNDA.t82 152.794
R2366 GNDA.n440 GNDA 145.695
R2367 GNDA.n446 GNDA.n3 142.683
R2368 GNDA.n254 GNDA.n253 142.683
R2369 GNDA.n443 GNDA.t102 141.935
R2370 GNDA.t12 GNDA.t1 141.353
R2371 GNDA.t5 GNDA.t13 141.353
R2372 GNDA.n332 GNDA.n331 135.083
R2373 GNDA.t7 GNDA.n289 133.083
R2374 GNDA.n209 GNDA.t287 132.465
R2375 GNDA.n263 GNDA.t284 132.465
R2376 GNDA.n270 GNDA.t233 132.465
R2377 GNDA.n243 GNDA.t253 132.465
R2378 GNDA.n161 GNDA.t11 122.556
R2379 GNDA.n251 GNDA.t285 119.444
R2380 GNDA.n229 GNDA.t234 119.444
R2381 GNDA.n331 GNDA.n330 115.415
R2382 GNDA.t9 GNDA.t78 113.91
R2383 GNDA.n88 GNDA.t274 108.365
R2384 GNDA.n436 GNDA.t206 108.365
R2385 GNDA.n100 GNDA.t179 108.365
R2386 GNDA.n422 GNDA.t154 108.365
R2387 GNDA.n126 GNDA.t224 108.365
R2388 GNDA.n124 GNDA.t230 108.365
R2389 GNDA.n129 GNDA.t190 108.365
R2390 GNDA.n408 GNDA.t213 108.365
R2391 GNDA.n404 GNDA.t259 108.365
R2392 GNDA.n304 GNDA.t165 108.365
R2393 GNDA.n140 GNDA.t294 108.365
R2394 GNDA.n360 GNDA.t170 108.365
R2395 GNDA.n362 GNDA.t227 108.365
R2396 GNDA.n349 GNDA.t129 108.365
R2397 GNDA.n348 GNDA.t281 108.365
R2398 GNDA.n345 GNDA.t201 108.365
R2399 GNDA.n344 GNDA.t187 108.365
R2400 GNDA.n183 GNDA.t237 108.365
R2401 GNDA.n182 GNDA.t244 108.365
R2402 GNDA.n179 GNDA.t144 108.365
R2403 GNDA.n178 GNDA.t256 108.365
R2404 GNDA.n315 GNDA.t182 108.365
R2405 GNDA.n318 GNDA.t158 108.365
R2406 GNDA.n401 GNDA.t289 108.365
R2407 GNDA.n400 GNDA.t247 108.365
R2408 GNDA.n121 GNDA.t250 108.365
R2409 GNDA.n90 GNDA.t148 108.365
R2410 GNDA.n103 GNDA.t197 108.365
R2411 GNDA.t99 GNDA.t0 103.383
R2412 GNDA.n384 GNDA.t155 103.008
R2413 GNDA.n217 GNDA.t116 100.053
R2414 GNDA.t80 GNDA.t113 96.993
R2415 GNDA.t3 GNDA.t101 95.1133
R2416 GNDA.n298 GNDA.t145 92.4817
R2417 GNDA.t92 GNDA.n215 88.4193
R2418 GNDA.n444 GNDA.n6 86.0925
R2419 GNDA.t87 GNDA.t6 84.587
R2420 GNDA.n1 GNDA.t117 83.4151
R2421 GNDA.n211 GNDA.t83 83.4151
R2422 GNDA.n257 GNDA.t115 83.4151
R2423 GNDA.n0 GNDA.t299 83.4151
R2424 GNDA.n251 GNDA.t106 80.6633
R2425 GNDA.n229 GNDA.t89 80.6633
R2426 GNDA.t114 GNDA.t118 75.9403
R2427 GNDA.n295 GNDA.n294 74.7248
R2428 GNDA.n294 GNDA.n284 74.7248
R2429 GNDA.n284 GNDA.n173 74.7248
R2430 GNDA.n378 GNDA.n156 74.7248
R2431 GNDA.n379 GNDA.n378 74.7248
R2432 GNDA.n380 GNDA.n379 74.7248
R2433 GNDA.n381 GNDA.n380 74.7248
R2434 GNDA.n248 GNDA.n247 74.3199
R2435 GNDA.n247 GNDA.n204 74.3199
R2436 GNDA.n366 GNDA.n173 73.514
R2437 GNDA.t0 GNDA.n368 70.6772
R2438 GNDA.t10 GNDA.t79 69.5494
R2439 GNDA.n170 GNDA.t9 65.414
R2440 GNDA.t108 GNDA.t149 65.414
R2441 GNDA.t15 GNDA.t108 65.0381
R2442 GNDA.t98 GNDA.n332 64.7271
R2443 GNDA.n286 GNDA.t91 59.7749
R2444 GNDA.n174 GNDA.t95 59.6649
R2445 GNDA.n187 GNDA.t97 59.6649
R2446 GNDA.n242 GNDA.t255 59.4285
R2447 GNDA.n269 GNDA.t236 59.4285
R2448 GNDA.n262 GNDA.t286 59.4285
R2449 GNDA.n260 GNDA.t288 59.4285
R2450 GNDA.t112 GNDA.t4 59.0231
R2451 GNDA.n253 GNDA.n252 58.5005
R2452 GNDA.n252 GNDA.n251 58.5005
R2453 GNDA.n446 GNDA.n445 58.5005
R2454 GNDA.n445 GNDA.n444 58.5005
R2455 GNDA.n441 GNDA.n440 58.5005
R2456 GNDA.n442 GNDA.n441 58.5005
R2457 GNDA.n147 GNDA.n11 58.5005
R2458 GNDA.n384 GNDA.n147 58.5005
R2459 GNDA.t11 GNDA.t87 56.7674
R2460 GNDA.n278 GNDA.t110 56.2845
R2461 GNDA.t17 GNDA.t114 54.5118
R2462 GNDA.n4 GNDA.n2 53.1823
R2463 GNDA.n216 GNDA.n4 53.1823
R2464 GNDA.n255 GNDA.n5 53.1823
R2465 GNDA.n217 GNDA.n5 53.1823
R2466 GNDA.n336 GNDA.n335 53.1823
R2467 GNDA.n337 GNDA.n336 53.1823
R2468 GNDA.n339 GNDA.n338 53.1823
R2469 GNDA.n338 GNDA.n337 53.1823
R2470 GNDA.t297 GNDA.n217 52.7416
R2471 GNDA.n245 GNDA.n240 49.3146
R2472 GNDA.n239 GNDA.n236 49.3146
R2473 GNDA.n265 GNDA.n207 49.3146
R2474 GNDA.n272 GNDA.n266 49.3146
R2475 GNDA.n238 GNDA.n237 49.1993
R2476 GNDA.n244 GNDA.n241 49.0972
R2477 GNDA.n271 GNDA.n267 49.0972
R2478 GNDA.n264 GNDA.n208 49.0972
R2479 GNDA.n292 GNDA.t85 48.4967
R2480 GNDA.n292 GNDA.t84 48.4967
R2481 GNDA.n369 GNDA.t112 48.4967
R2482 GNDA.n376 GNDA.t79 48.4967
R2483 GNDA.t88 GNDA.n160 48.4967
R2484 GNDA.n160 GNDA.t120 48.4967
R2485 GNDA.t82 GNDA.t297 47.3123
R2486 GNDA.t101 GNDA.t7 46.2411
R2487 GNDA.t16 GNDA.t92 45.7611
R2488 GNDA.t104 GNDA.t14 45.7611
R2489 GNDA.t85 GNDA.t17 42.4817
R2490 GNDA.n225 GNDA.n224 41.7887
R2491 GNDA.n196 GNDA.n195 41.7862
R2492 GNDA.n330 GNDA.n196 41.7862
R2493 GNDA.n329 GNDA.n328 41.7862
R2494 GNDA.n330 GNDA.n329 41.7862
R2495 GNDA.n149 GNDA.n93 41.7862
R2496 GNDA.n384 GNDA.n149 41.7862
R2497 GNDA.n390 GNDA.n139 41.7862
R2498 GNDA.n384 GNDA.n139 41.7862
R2499 GNDA.n190 GNDA.n188 39.0005
R2500 GNDA.n278 GNDA.n190 39.0005
R2501 GNDA.n191 GNDA.n189 39.0005
R2502 GNDA.n332 GNDA.n191 39.0005
R2503 GNDA.n288 GNDA.n287 39.0005
R2504 GNDA.n289 GNDA.n288 39.0005
R2505 GNDA.n169 GNDA.n164 39.0005
R2506 GNDA.n170 GNDA.n169 39.0005
R2507 GNDA.n162 GNDA.n155 39.0005
R2508 GNDA.n162 GNDA.n161 39.0005
R2509 GNDA.n297 GNDA.n296 39.0005
R2510 GNDA.n298 GNDA.n297 39.0005
R2511 GNDA.n280 GNDA.n199 39.0005
R2512 GNDA.n280 GNDA.n279 39.0005
R2513 GNDA.n383 GNDA.n382 39.0005
R2514 GNDA.n384 GNDA.n383 39.0005
R2515 GNDA.t4 GNDA.t99 37.9704
R2516 GNDA.t86 GNDA.n286 37.2185
R2517 GNDA.n219 GNDA.n206 36.563
R2518 GNDA.n276 GNDA.n275 36.563
R2519 GNDA.n277 GNDA.n276 36.563
R2520 GNDA.n369 GNDA.t2 33.8351
R2521 GNDA.t120 GNDA.t15 31.9554
R2522 GNDA.n254 GNDA.n213 30.1181
R2523 GNDA.n225 GNDA.n3 30.1181
R2524 GNDA.t1 GNDA.t86 29.6997
R2525 GNDA.n224 GNDA.n223 27.8576
R2526 GNDA.n223 GNDA.n6 27.8576
R2527 GNDA.n221 GNDA.n214 27.8576
R2528 GNDA.n251 GNDA.n214 27.8576
R2529 GNDA.n227 GNDA.n226 27.8576
R2530 GNDA.n229 GNDA.n227 27.8576
R2531 GNDA.n233 GNDA.n232 27.8576
R2532 GNDA.n232 GNDA.n6 27.8576
R2533 GNDA.n250 GNDA.n249 27.8576
R2534 GNDA.n251 GNDA.n250 27.8576
R2535 GNDA.n230 GNDA.n228 27.8576
R2536 GNDA.n230 GNDA.n229 27.8576
R2537 GNDA.n153 GNDA.n146 27.8576
R2538 GNDA.n384 GNDA.n146 27.8576
R2539 GNDA.n356 GNDA.n172 27.8576
R2540 GNDA.n330 GNDA.n172 27.8576
R2541 GNDA.t78 GNDA.t10 27.4441
R2542 GNDA.n194 GNDA.n177 26.5914
R2543 GNDA.n330 GNDA.n194 26.5914
R2544 GNDA.n386 GNDA.n385 26.5914
R2545 GNDA.n385 GNDA.n384 26.5914
R2546 GNDA.t113 GNDA.t8 25.1885
R2547 GNDA.n201 GNDA.n200 24.3755
R2548 GNDA.n201 GNDA.n192 24.3755
R2549 GNDA.n152 GNDA.n150 24.3755
R2550 GNDA.n160 GNDA.n150 24.3755
R2551 GNDA.n375 GNDA.n374 24.3755
R2552 GNDA.n376 GNDA.n375 24.3755
R2553 GNDA.n371 GNDA.n370 24.3755
R2554 GNDA.n370 GNDA.n369 24.3755
R2555 GNDA.n291 GNDA.n290 24.3755
R2556 GNDA.n292 GNDA.n291 24.3755
R2557 GNDA.n282 GNDA.n281 24.3755
R2558 GNDA.n281 GNDA.n192 24.3755
R2559 GNDA.n380 GNDA.n151 24.3755
R2560 GNDA.n160 GNDA.n151 24.3755
R2561 GNDA.n378 GNDA.n377 24.3755
R2562 GNDA.n377 GNDA.n376 24.3755
R2563 GNDA.n173 GNDA.n167 24.3755
R2564 GNDA.n369 GNDA.n167 24.3755
R2565 GNDA.n294 GNDA.n293 24.3755
R2566 GNDA.n293 GNDA.n292 24.3755
R2567 GNDA.t13 GNDA.t80 19.1734
R2568 GNDA.n161 GNDA.t5 18.7975
R2569 GNDA.t8 GNDA.t119 18.4216
R2570 GNDA.n274 GNDA.n203 15.8113
R2571 GNDA.n203 GNDA.n6 15.8113
R2572 GNDA.t91 GNDA.t2 14.6622
R2573 GNDA.n444 GNDA.t104 13.9614
R2574 GNDA.t14 GNDA.n443 12.4102
R2575 GNDA.t6 GNDA.t88 12.4065
R2576 GNDA.n215 GNDA.n6 11.6346
R2577 GNDA.t145 GNDA.t118 10.9028
R2578 GNDA.t149 GNDA.t155 10.9028
R2579 GNDA.n330 GNDA.n298 10.5268
R2580 GNDA.n237 GNDA.t288 10.3318
R2581 GNDA.n237 GNDA.t107 10.3318
R2582 GNDA.n240 GNDA.t105 10.3318
R2583 GNDA.n240 GNDA.t111 10.3318
R2584 GNDA.n236 GNDA.t300 10.3318
R2585 GNDA.n236 GNDA.t93 10.3318
R2586 GNDA.n241 GNDA.t90 10.3318
R2587 GNDA.n241 GNDA.t254 10.3318
R2588 GNDA.n267 GNDA.t109 10.3318
R2589 GNDA.n267 GNDA.t235 10.3318
R2590 GNDA.n207 GNDA.t298 10.3318
R2591 GNDA.n207 GNDA.t302 10.3318
R2592 GNDA.n266 GNDA.t301 10.3318
R2593 GNDA.n266 GNDA.t103 10.3318
R2594 GNDA.t286 GNDA.n208 10.3318
R2595 GNDA.n208 GNDA.t303 10.3318
R2596 GNDA.n235 GNDA.n6 10.0867
R2597 GNDA.n247 GNDA.n235 10.0867
R2598 GNDA.n438 GNDA.n89 8.8505
R2599 GNDA.n438 GNDA.n437 8.8505
R2600 GNDA.n289 GNDA.t12 8.27118
R2601 GNDA.n430 GNDA.n95 5.79258
R2602 GNDA.n368 GNDA.n95 5.79258
R2603 GNDA.n367 GNDA.n366 5.79258
R2604 GNDA.n368 GNDA.n367 5.79258
R2605 GNDA.n86 GNDA.t263 5.6933
R2606 GNDA.n392 GNDA.n137 5.68011
R2607 GNDA.n368 GNDA.n137 5.68011
R2608 GNDA.n354 GNDA.n168 5.68011
R2609 GNDA.n368 GNDA.n168 5.68011
R2610 GNDA.n326 GNDA.n171 5.68011
R2611 GNDA.n368 GNDA.n171 5.68011
R2612 GNDA.n368 GNDA.n170 5.26366
R2613 GNDA.n431 GNDA.n93 4.89462
R2614 GNDA.n195 GNDA.n94 4.89462
R2615 GNDA.n154 GNDA.n153 4.89462
R2616 GNDA.n357 GNDA.n356 4.89462
R2617 GNDA.n376 GNDA.t119 4.88772
R2618 GNDA.n365 GNDA.n361 4.86612
R2619 GNDA.n365 GNDA.n364 4.86612
R2620 GNDA.n353 GNDA.n343 4.57238
R2621 GNDA.n353 GNDA.n352 4.57238
R2622 GNDA.n9 GNDA.n7 4.36617
R2623 GNDA.n286 GNDA.n7 4.36617
R2624 GNDA.n439 GNDA.n8 4.36617
R2625 GNDA.n286 GNDA.n8 4.36617
R2626 GNDA.t100 GNDA.t96 4.2218
R2627 GNDA.n337 GNDA.n192 4.2218
R2628 GNDA.t81 GNDA.t94 4.2218
R2629 GNDA.n413 GNDA.n105 3.91726
R2630 GNDA GNDA.n258 3.2614
R2631 GNDA.n295 GNDA.n176 2.42212
R2632 GNDA.t84 GNDA.t3 1.8802
R2633 GNDA.t116 GNDA.t16 1.55171
R2634 GNDA.n334 GNDA.n333 1.44894
R2635 GNDA.n364 GNDA.n363 1.42278
R2636 GNDA.n242 GNDA.n205 1.27784
R2637 GNDA.n435 GNDA.n434 1.23175
R2638 GNDA.n366 GNDA.n156 1.21131
R2639 GNDA.n388 GNDA.n387 1.13129
R2640 GNDA.n363 GNDA.n142 1.13126
R2641 GNDA.n387 GNDA.n142 1.13028
R2642 GNDA.n342 GNDA.n186 1.12238
R2643 GNDA.n319 GNDA.n186 1.12238
R2644 GNDA.n25 GNDA.t210 1.082
R2645 GNDA.n333 GNDA.n187 1.04581
R2646 GNDA.n434 GNDA.n11 0.9305
R2647 GNDA.n440 GNDA.n10 0.9305
R2648 GNDA.n310 GNDA.n309 0.91925
R2649 GNDA.n309 GNDA.n308 0.91925
R2650 GNDA.n308 GNDA.n307 0.91925
R2651 GNDA.n325 GNDA.n324 0.91925
R2652 GNDA.n324 GNDA.n323 0.91925
R2653 GNDA.n323 GNDA.n322 0.91925
R2654 GNDA.n322 GNDA.n321 0.91925
R2655 GNDA.n397 GNDA.n396 0.91925
R2656 GNDA.n396 GNDA.n395 0.91925
R2657 GNDA.n395 GNDA.n394 0.91925
R2658 GNDA.n135 GNDA.n134 0.91925
R2659 GNDA.n134 GNDA.n133 0.91925
R2660 GNDA.n133 GNDA.n132 0.91925
R2661 GNDA.n32 GNDA.t219 0.909177
R2662 GNDA.n262 GNDA.n261 0.908052
R2663 GNDA.n325 GNDA 0.883312
R2664 GNDA.n86 GNDA.n10 0.873417
R2665 GNDA.n447 GNDA.n446 0.845955
R2666 GNDA.n253 GNDA.n212 0.845955
R2667 GNDA.n261 GNDA.n260 0.833625
R2668 GNDA.n212 GNDA.n211 0.8255
R2669 GNDA.n447 GNDA.n1 0.8255
R2670 GNDA.n239 GNDA.n238 0.821833
R2671 GNDA.n245 GNDA.n244 0.788781
R2672 GNDA.n272 GNDA.n271 0.788781
R2673 GNDA.n265 GNDA.n264 0.788781
R2674 GNDA.n340 GNDA.n339 0.7755
R2675 GNDA.n335 GNDA.n334 0.7755
R2676 GNDA.n256 GNDA.n255 0.7755
R2677 GNDA.n210 GNDA.n2 0.7755
R2678 GNDA.n434 GNDA.n433 0.747767
R2679 GNDA.n104 GNDA.n10 0.74425
R2680 GNDA.n29 GNDA.t174 0.7295
R2681 GNDA.n31 GNDA.t124 0.7295
R2682 GNDA.n38 GNDA.t241 0.7295
R2683 GNDA.n40 GNDA.t128 0.7295
R2684 GNDA.n42 GNDA.t196 0.7295
R2685 GNDA.n44 GNDA.t267 0.7295
R2686 GNDA.n46 GNDA.t269 0.7295
R2687 GNDA.n48 GNDA.t164 0.7295
R2688 GNDA.n50 GNDA.t217 0.7295
R2689 GNDA.n52 GNDA.t133 0.7295
R2690 GNDA.n54 GNDA.t205 0.7295
R2691 GNDA.n56 GNDA.t293 0.7295
R2692 GNDA.n58 GNDA.t141 0.7295
R2693 GNDA.n60 GNDA.t243 0.7295
R2694 GNDA.n67 GNDA.t122 0.7295
R2695 GNDA.n15 GNDA.t271 0.7295
R2696 GNDA.n16 GNDA.t162 0.7295
R2697 GNDA.n17 GNDA.t212 0.7295
R2698 GNDA.n18 GNDA.t280 0.7295
R2699 GNDA.n69 GNDA.t221 0.7295
R2700 GNDA.n71 GNDA.t137 0.7295
R2701 GNDA.n73 GNDA.t265 0.7295
R2702 GNDA.n75 GNDA.t176 0.7295
R2703 GNDA.n77 GNDA.t273 0.7295
R2704 GNDA.n79 GNDA.t143 0.7295
R2705 GNDA.n13 GNDA.t178 0.7295
R2706 GNDA.n22 GNDA.t223 0.7295
R2707 GNDA.n23 GNDA.t126 0.7295
R2708 GNDA.n24 GNDA.t186 0.7295
R2709 GNDA.n81 GNDA.t169 0.7295
R2710 GNDA.n83 GNDA.t153 0.7295
R2711 GNDA.n28 GNDA.t139 0.7295
R2712 GNDA.n25 GNDA.t278 0.7295
R2713 GNDA.n26 GNDA.t135 0.7295
R2714 GNDA.n27 GNDA.t194 0.7295
R2715 GNDA.t263 GNDA.n85 0.7295
R2716 GNDA.n433 GNDA.n432 0.721109
R2717 GNDA.n389 GNDA.n92 0.71857
R2718 GNDA.n432 GNDA.n92 0.717584
R2719 GNDA.n389 GNDA.n388 0.717564
R2720 GNDA.n390 GNDA.n389 0.715885
R2721 GNDA.n328 GNDA.n106 0.715885
R2722 GNDA.n412 GNDA.n94 0.715885
R2723 GNDA.n432 GNDA.n431 0.715885
R2724 GNDA.n319 GNDA.n106 0.709875
R2725 GNDA.n411 GNDA.n106 0.709875
R2726 GNDA.n412 GNDA.n411 0.709875
R2727 GNDA.n413 GNDA.n412 0.709875
R2728 GNDA.n189 GNDA.n175 0.664786
R2729 GNDA.n333 GNDA.n188 0.664786
R2730 GNDA.n361 GNDA.n359 0.615539
R2731 GNDA.n341 GNDA.n340 0.609875
R2732 GNDA.n343 GNDA.n342 0.59425
R2733 GNDA.n411 GNDA.n410 0.59425
R2734 GNDA.n352 GNDA.n142 0.587766
R2735 GNDA.n119 GNDA.n92 0.58772
R2736 GNDA.n275 GNDA.n205 0.58175
R2737 GNDA.n261 GNDA.n206 0.58175
R2738 GNDA.n448 GNDA.n447 0.55675
R2739 GNDA.n415 GNDA.n414 0.51137
R2740 GNDA.n416 GNDA.n415 0.51137
R2741 GNDA.n429 GNDA.n418 0.51137
R2742 GNDA.n429 GNDA.n428 0.51137
R2743 GNDA.n428 GNDA.n427 0.51137
R2744 GNDA.n427 GNDA.n426 0.51137
R2745 GNDA.n426 GNDA.n425 0.51137
R2746 GNDA.n394 GNDA.n393 0.459875
R2747 GNDA.n393 GNDA.n135 0.459875
R2748 GNDA.n363 GNDA.n154 0.443357
R2749 GNDA.n358 GNDA.n357 0.443357
R2750 GNDA.n186 GNDA.n177 0.443357
R2751 GNDA.n387 GNDA.n386 0.443357
R2752 GNDA.n334 GNDA.n174 0.403625
R2753 GNDA.n340 GNDA.n187 0.403625
R2754 GNDA.n211 GNDA.n210 0.403625
R2755 GNDA.n210 GNDA.n1 0.403625
R2756 GNDA.n246 GNDA.n239 0.403625
R2757 GNDA.n246 GNDA.n245 0.403625
R2758 GNDA.n273 GNDA.n265 0.403625
R2759 GNDA.n273 GNDA.n272 0.403625
R2760 GNDA.n257 GNDA.n256 0.403625
R2761 GNDA.n256 GNDA.n0 0.403625
R2762 GNDA.n268 GNDA 0.392688
R2763 GNDA.n269 GNDA.n268 0.368469
R2764 GNDA.n87 GNDA.n86 0.360917
R2765 GNDA.n268 GNDA.n205 0.359875
R2766 GNDA.n16 GNDA.n15 0.353
R2767 GNDA.n17 GNDA.n16 0.353
R2768 GNDA.n18 GNDA.n17 0.353
R2769 GNDA.n22 GNDA.n13 0.353
R2770 GNDA.n23 GNDA.n22 0.353
R2771 GNDA.n24 GNDA.n23 0.353
R2772 GNDA.n26 GNDA.n25 0.353
R2773 GNDA.n27 GNDA.n26 0.353
R2774 GNDA.n141 GNDA.n140 0.338152
R2775 GNDA.n361 GNDA.n360 0.338152
R2776 GNDA.n364 GNDA.n362 0.338152
R2777 GNDA.n352 GNDA.n347 0.338152
R2778 GNDA.n352 GNDA.n351 0.338152
R2779 GNDA.n343 GNDA.n181 0.338152
R2780 GNDA.n343 GNDA.n185 0.338152
R2781 GNDA.n320 GNDA.n318 0.338152
R2782 GNDA.n258 GNDA.n212 0.332591
R2783 GNDA.n410 GNDA.n397 0.33175
R2784 GNDA.n132 GNDA.n119 0.33175
R2785 GNDA.n67 GNDA.n15 0.3295
R2786 GNDA.n60 GNDA.n18 0.3295
R2787 GNDA.n79 GNDA.n13 0.3295
R2788 GNDA.n48 GNDA.n24 0.3295
R2789 GNDA.n28 GNDA.n27 0.3295
R2790 GNDA.n414 GNDA.n413 0.314359
R2791 GNDA.n320 GNDA.n319 0.3005
R2792 GNDA.n388 GNDA.n141 0.293992
R2793 GNDA.n310 GNDA.n301 0.291659
R2794 GNDA.n309 GNDA.n302 0.291659
R2795 GNDA.n308 GNDA.n303 0.291659
R2796 GNDA.n325 GNDA.n311 0.291659
R2797 GNDA.n324 GNDA.n312 0.291659
R2798 GNDA.n323 GNDA.n313 0.291659
R2799 GNDA.n322 GNDA.n314 0.291659
R2800 GNDA.n396 GNDA.n107 0.291659
R2801 GNDA.n396 GNDA.n108 0.291659
R2802 GNDA.n395 GNDA.n109 0.291659
R2803 GNDA.n395 GNDA.n110 0.291659
R2804 GNDA.n394 GNDA.n111 0.291659
R2805 GNDA.n394 GNDA.n112 0.291659
R2806 GNDA.n135 GNDA.n113 0.291659
R2807 GNDA.n135 GNDA.n114 0.291659
R2808 GNDA.n134 GNDA.n115 0.291659
R2809 GNDA.n134 GNDA.n116 0.291659
R2810 GNDA.n133 GNDA.n117 0.291659
R2811 GNDA.n133 GNDA.n118 0.291659
R2812 GNDA.n102 GNDA.n100 0.288543
R2813 GNDA.n424 GNDA.n422 0.288543
R2814 GNDA.n128 GNDA.n126 0.288543
R2815 GNDA.n131 GNDA.n129 0.288543
R2816 GNDA.n129 GNDA.n128 0.288543
R2817 GNDA.n409 GNDA.n404 0.288543
R2818 GNDA.n306 GNDA.n304 0.288543
R2819 GNDA.n351 GNDA.n348 0.288543
R2820 GNDA.n351 GNDA.n349 0.288543
R2821 GNDA.n347 GNDA.n344 0.288543
R2822 GNDA.n347 GNDA.n345 0.288543
R2823 GNDA.n185 GNDA.n182 0.288543
R2824 GNDA.n185 GNDA.n183 0.288543
R2825 GNDA.n181 GNDA.n178 0.288543
R2826 GNDA.n181 GNDA.n179 0.288543
R2827 GNDA.n317 GNDA.n315 0.288543
R2828 GNDA.n403 GNDA.n400 0.288543
R2829 GNDA.n400 GNDA.n399 0.288543
R2830 GNDA.n403 GNDA.n401 0.288543
R2831 GNDA.n409 GNDA.n408 0.288543
R2832 GNDA.n408 GNDA.n407 0.288543
R2833 GNDA.n123 GNDA.n121 0.288543
R2834 GNDA.n125 GNDA.n124 0.288543
R2835 GNDA.n124 GNDA.n123 0.288543
R2836 GNDA.n21 GNDA.t185 0.28175
R2837 GNDA.n20 GNDA.t125 0.28175
R2838 GNDA.n19 GNDA.t222 0.28175
R2839 GNDA.n14 GNDA.t177 0.28175
R2840 GNDA.n84 GNDA.t262 0.28175
R2841 GNDA.n82 GNDA.t152 0.28175
R2842 GNDA.n80 GNDA.t168 0.28175
R2843 GNDA.n78 GNDA.t142 0.28175
R2844 GNDA.n76 GNDA.t272 0.28175
R2845 GNDA.n74 GNDA.t175 0.28175
R2846 GNDA.n72 GNDA.t264 0.28175
R2847 GNDA.n70 GNDA.t136 0.28175
R2848 GNDA.n68 GNDA.t220 0.28175
R2849 GNDA.n66 GNDA.t121 0.28175
R2850 GNDA.n65 GNDA.t270 0.28175
R2851 GNDA.n64 GNDA.t161 0.28175
R2852 GNDA.n63 GNDA.t211 0.28175
R2853 GNDA.n62 GNDA.t279 0.28175
R2854 GNDA.n61 GNDA.t242 0.28175
R2855 GNDA.n59 GNDA.t140 0.28175
R2856 GNDA.n57 GNDA.t292 0.28175
R2857 GNDA.n55 GNDA.t204 0.28175
R2858 GNDA.n53 GNDA.t132 0.28175
R2859 GNDA.n51 GNDA.t216 0.28175
R2860 GNDA.n49 GNDA.t163 0.28175
R2861 GNDA.n47 GNDA.t268 0.28175
R2862 GNDA.n45 GNDA.t266 0.28175
R2863 GNDA.n43 GNDA.t195 0.28175
R2864 GNDA.n41 GNDA.t127 0.28175
R2865 GNDA.n39 GNDA.t240 0.28175
R2866 GNDA.n37 GNDA.t138 0.28175
R2867 GNDA.n36 GNDA.t193 0.28175
R2868 GNDA.n35 GNDA.t134 0.28175
R2869 GNDA.n34 GNDA.t277 0.28175
R2870 GNDA.n33 GNDA.t209 0.28175
R2871 GNDA.n32 GNDA.t218 0.28175
R2872 GNDA.n30 GNDA.t123 0.28175
R2873 GNDA.n12 GNDA.t173 0.28175
R2874 GNDA GNDA.n105 0.271125
R2875 GNDA.n448 GNDA.n0 0.26925
R2876 GNDA.n418 GNDA.n417 0.262728
R2877 GNDA.n429 GNDA.n96 0.261171
R2878 GNDA.n415 GNDA.n99 0.261171
R2879 GNDA.n416 GNDA.n98 0.261171
R2880 GNDA.n418 GNDA.n97 0.261171
R2881 GNDA.n428 GNDA.n419 0.261171
R2882 GNDA.n427 GNDA.n420 0.261171
R2883 GNDA.n426 GNDA.n421 0.261171
R2884 GNDA.n247 GNDA.n246 0.251851
R2885 GNDA.n274 GNDA.n273 0.251851
R2886 GNDA.n417 GNDA.n416 0.249141
R2887 GNDA.n21 GNDA.n20 0.242354
R2888 GNDA.n20 GNDA.n19 0.242354
R2889 GNDA.n19 GNDA.n14 0.242354
R2890 GNDA.n65 GNDA.n64 0.242354
R2891 GNDA.n64 GNDA.n63 0.242354
R2892 GNDA.n63 GNDA.n62 0.242354
R2893 GNDA.n36 GNDA.n35 0.242354
R2894 GNDA.n35 GNDA.n34 0.242354
R2895 GNDA.n34 GNDA.n33 0.242354
R2896 GNDA.n49 GNDA.n21 0.218854
R2897 GNDA.n78 GNDA.n14 0.218854
R2898 GNDA.n66 GNDA.n65 0.218854
R2899 GNDA.n62 GNDA.n61 0.218854
R2900 GNDA.n37 GNDA.n36 0.218854
R2901 GNDA.n33 GNDA.n32 0.218854
R2902 GNDA.n359 GNDA.n174 0.20675
R2903 GNDA.n258 GNDA.n257 0.20675
R2904 GNDA.n84 GNDA.n83 0.205635
R2905 GNDA.n82 GNDA.n81 0.205635
R2906 GNDA.n80 GNDA.n79 0.205635
R2907 GNDA.n78 GNDA.n77 0.205635
R2908 GNDA.n76 GNDA.n75 0.205635
R2909 GNDA.n74 GNDA.n73 0.205635
R2910 GNDA.n72 GNDA.n71 0.205635
R2911 GNDA.n70 GNDA.n69 0.205635
R2912 GNDA.n68 GNDA.n67 0.205635
R2913 GNDA.n60 GNDA.n59 0.205635
R2914 GNDA.n58 GNDA.n57 0.205635
R2915 GNDA.n56 GNDA.n55 0.205635
R2916 GNDA.n54 GNDA.n53 0.205635
R2917 GNDA.n52 GNDA.n51 0.205635
R2918 GNDA.n50 GNDA.n49 0.205635
R2919 GNDA.n48 GNDA.n47 0.205635
R2920 GNDA.n46 GNDA.n45 0.205635
R2921 GNDA.n44 GNDA.n43 0.205635
R2922 GNDA.n42 GNDA.n41 0.205635
R2923 GNDA.n40 GNDA.n39 0.205635
R2924 GNDA.n38 GNDA.n37 0.205635
R2925 GNDA.n32 GNDA.n31 0.205635
R2926 GNDA.n30 GNDA.n29 0.205635
R2927 GNDA.n85 GNDA.n12 0.205635
R2928 GNDA.n307 GNDA.n306 0.204006
R2929 GNDA.n321 GNDA.n317 0.204006
R2930 GNDA.n410 GNDA.n403 0.204006
R2931 GNDA.n410 GNDA.n409 0.204006
R2932 GNDA.n399 GNDA.n397 0.204006
R2933 GNDA.n407 GNDA.n397 0.204006
R2934 GNDA.n132 GNDA.n125 0.204006
R2935 GNDA.n132 GNDA.n131 0.204006
R2936 GNDA.n123 GNDA.n119 0.204006
R2937 GNDA.n128 GNDA.n119 0.204006
R2938 GNDA.n433 GNDA.n91 0.199748
R2939 GNDA.n85 GNDA.n84 0.180177
R2940 GNDA.n83 GNDA.n82 0.180177
R2941 GNDA.n81 GNDA.n80 0.180177
R2942 GNDA.n79 GNDA.n78 0.180177
R2943 GNDA.n77 GNDA.n76 0.180177
R2944 GNDA.n75 GNDA.n74 0.180177
R2945 GNDA.n73 GNDA.n72 0.180177
R2946 GNDA.n71 GNDA.n70 0.180177
R2947 GNDA.n69 GNDA.n68 0.180177
R2948 GNDA.n67 GNDA.n66 0.180177
R2949 GNDA.n61 GNDA.n60 0.180177
R2950 GNDA.n59 GNDA.n58 0.180177
R2951 GNDA.n57 GNDA.n56 0.180177
R2952 GNDA.n55 GNDA.n54 0.180177
R2953 GNDA.n53 GNDA.n52 0.180177
R2954 GNDA.n51 GNDA.n50 0.180177
R2955 GNDA.n49 GNDA.n48 0.180177
R2956 GNDA.n47 GNDA.n46 0.180177
R2957 GNDA.n45 GNDA.n44 0.180177
R2958 GNDA.n43 GNDA.n42 0.180177
R2959 GNDA.n41 GNDA.n40 0.180177
R2960 GNDA.n39 GNDA.n38 0.180177
R2961 GNDA.n37 GNDA.n28 0.180177
R2962 GNDA.n31 GNDA.n30 0.180177
R2963 GNDA.n29 GNDA.n12 0.180177
R2964 GNDA.n414 GNDA.n102 0.173518
R2965 GNDA.n425 GNDA.n424 0.173518
R2966 GNDA.n342 GNDA.n341 0.146789
R2967 GNDA.n341 GNDA.n175 0.139475
R2968 GNDA.n359 GNDA.n358 0.1255
R2969 GNDA.n425 GNDA.n91 0.112592
R2970 GNDA.n244 GNDA.n243 0.101281
R2971 GNDA.n243 GNDA.n242 0.101281
R2972 GNDA.n271 GNDA.n270 0.101281
R2973 GNDA.n270 GNDA.n269 0.101281
R2974 GNDA.n263 GNDA.n262 0.101281
R2975 GNDA.n264 GNDA.n263 0.101281
R2976 GNDA.n366 GNDA.n365 0.0963763
R2977 GNDA.n354 GNDA.n353 0.0963763
R2978 GNDA.n326 GNDA.n325 0.0963763
R2979 GNDA.n393 GNDA.n392 0.0963763
R2980 GNDA.n430 GNDA.n429 0.0963763
R2981 GNDA.n102 GNDA.n101 0.0881524
R2982 GNDA.n424 GNDA.n423 0.0881524
R2983 GNDA.n306 GNDA.n305 0.0881524
R2984 GNDA.n347 GNDA.n346 0.0881524
R2985 GNDA.n351 GNDA.n350 0.0881524
R2986 GNDA.n181 GNDA.n180 0.0881524
R2987 GNDA.n185 GNDA.n184 0.0881524
R2988 GNDA.n317 GNDA.n316 0.0881524
R2989 GNDA.n403 GNDA.n402 0.0881524
R2990 GNDA.n409 GNDA.n405 0.0881524
R2991 GNDA.n399 GNDA.n398 0.0881524
R2992 GNDA.n407 GNDA.n406 0.0881524
R2993 GNDA.n125 GNDA.n120 0.0881524
R2994 GNDA.n131 GNDA.n130 0.0881524
R2995 GNDA.n123 GNDA.n122 0.0881524
R2996 GNDA.n128 GNDA.n127 0.0881524
R2997 GNDA.n260 GNDA.n259 0.077375
R2998 GNDA.n417 GNDA.n9 0.072593
R2999 GNDA.n439 GNDA.n438 0.072593
R3000 GNDA.n436 GNDA.n435 0.0591735
R3001 GNDA.n88 GNDA.n87 0.0591735
R3002 GNDA.n437 GNDA.n436 0.0489694
R3003 GNDA.n89 GNDA.n88 0.0489694
R3004 GNDA GNDA.n448 0.047375
R3005 GNDA.n259 GNDA 0.0390417
R3006 GNDA.n307 GNDA.n141 0.038
R3007 GNDA.n321 GNDA.n320 0.038
R3008 GNDA GNDA.n310 0.0364375
R3009 GNDA.n238 GNDA.n209 0.03425
R3010 GNDA.n358 GNDA.n175 0.0144752
R3011 GNDA.n105 GNDA.n104 0.009875
R3012 GNDA.n91 GNDA.n90 0.00912069
R3013 GNDA.n104 GNDA.n103 0.00912069
R3014 GNDA.n259 GNDA.n209 0.00425
R3015 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t8 142.458
R3016 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t0 142.458
R3017 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t23 141.674
R3018 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t26 141.674
R3019 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t10 140.891
R3020 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t13 140.891
R3021 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t30 139.879
R3022 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t21 139.879
R3023 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t22 139.879
R3024 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t18 139.879
R3025 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t27 139.879
R3026 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t16 139.879
R3027 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t31 139.879
R3028 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t17 139.879
R3029 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t19 139.879
R3030 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t29 139.879
R3031 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t24 135.441
R3032 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t25 135.441
R3033 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t28 135.435
R3034 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t20 135.435
R3035 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t14 134.732
R3036 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t2 134.732
R3037 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t12 134.732
R3038 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t7 134.732
R3039 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t6 134.732
R3040 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t1 134.732
R3041 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t9 134.732
R3042 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t15 134.732
R3043 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t4 134.712
R3044 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t11 134.712
R3045 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t5 134.712
R3046 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t3 134.712
R3047 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n12 5.61925
R3048 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n20 4.9505
R3049 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n9 4.57291
R3050 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n4 4.57291
R3051 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n0 4.5005
R3052 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n2 4.5005
R3053 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n7 4.5005
R3054 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n11 4.5005
R3055 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n5 4.05258
R3056 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n6 4.02292
R3057 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n1 3.78175
R3058 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n21 3.67541
R3059 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n24 3.5885
R3060 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n15 3.5885
R3061 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n28 3.4105
R3062 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n13 3.4105
R3063 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n27 3.38383
R3064 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n3 3.13383
R3065 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n8 3.13383
R3066 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n23 3.113
R3067 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n10 2.21508
R3068 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n25 1.79633
R3069 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n16 1.79633
R3070 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n18 1.54633
R3071 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n22 1.338
R3072 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n26 1.338
R3073 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n17 1.338
R3074 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n19 1.338
R3075 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n29 1.05159
R3076 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n14 0.516076
R3077 opa_folded_cascode_0.monticelli_top_0.B.n4 opa_folded_cascode_0.monticelli_top_0.B.t6 118.626
R3078 opa_folded_cascode_0.monticelli_top_0.B.n5 opa_folded_cascode_0.monticelli_top_0.B.t8 118.626
R3079 opa_folded_cascode_0.monticelli_top_0.B.n4 opa_folded_cascode_0.monticelli_top_0.B.t9 118.005
R3080 opa_folded_cascode_0.monticelli_top_0.B.n5 opa_folded_cascode_0.monticelli_top_0.B.t7 118.005
R3081 opa_folded_cascode_0.monticelli_top_0.B.n2 opa_folded_cascode_0.monticelli_top_0.B.t4 70.0103
R3082 opa_folded_cascode_0.monticelli_top_0.B.n3 opa_folded_cascode_0.monticelli_top_0.B.t5 69.7645
R3083 opa_folded_cascode_0.monticelli_top_0.B.n1 opa_folded_cascode_0.monticelli_top_0.B.t0 69.622
R3084 opa_folded_cascode_0.monticelli_top_0.B.n1 opa_folded_cascode_0.monticelli_top_0.B.t1 59.4447
R3085 opa_folded_cascode_0.monticelli_top_0.B.n0 opa_folded_cascode_0.monticelli_top_0.B.t3 50.8746
R3086 opa_folded_cascode_0.monticelli_top_0.B.n0 opa_folded_cascode_0.monticelli_top_0.B.t2 49.6789
R3087 opa_folded_cascode_0.monticelli_top_0.B opa_folded_cascode_0.monticelli_top_0.B.n0 16.5734
R3088 opa_folded_cascode_0.monticelli_top_0.B.n2 opa_folded_cascode_0.monticelli_top_0.B.n1 11.3963
R3089 opa_folded_cascode_0.monticelli_top_0.B.n7 opa_folded_cascode_0.monticelli_top_0.B.n6 9.83175
R3090 opa_folded_cascode_0.monticelli_top_0.B.n7 opa_folded_cascode_0.monticelli_top_0.B.n3 2.93383
R3091 opa_folded_cascode_0.monticelli_top_0.B.n3 opa_folded_cascode_0.monticelli_top_0.B.n2 2.42967
R3092 opa_folded_cascode_0.monticelli_top_0.B opa_folded_cascode_0.monticelli_top_0.B.n7 2.11508
R3093 opa_folded_cascode_0.monticelli_top_0.B.n6 opa_folded_cascode_0.monticelli_top_0.B.n4 0.629667
R3094 opa_folded_cascode_0.monticelli_top_0.B.n6 opa_folded_cascode_0.monticelli_top_0.B.n5 0.629667
R3095 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t10 228.174
R3096 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t15 228.174
R3097 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t5 228.174
R3098 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t11 228.174
R3099 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t14 226.853
R3100 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t7 226.853
R3101 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t8 226.853
R3102 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t9 226.853
R3103 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t6 226.853
R3104 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t1 226.853
R3105 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t4 226.853
R3106 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t13 226.853
R3107 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t3 226.853
R3108 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t12 226.853
R3109 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t2 226.853
R3110 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t0 226.853
R3111 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t16 221.911
R3112 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n23 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t23 221.911
R3113 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t24 221.911
R3114 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n24 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t31 221.911
R3115 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t26 221.911
R3116 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n26 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t22 221.911
R3117 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t17 221.911
R3118 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n22 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t20 221.911
R3119 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t30 221.911
R3120 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n18 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t18 221.911
R3121 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t21 221.911
R3122 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n19 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t29 221.911
R3123 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t25 221.911
R3124 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n16 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t27 221.911
R3125 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t28 221.911
R3126 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n15 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t19 221.911
R3127 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n23 7.63383
R3128 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n15 7.63383
R3129 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n18 7.63383
R3130 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n22 7.49842
R3131 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n6 5.05408
R3132 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n26 4.5005
R3133 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n25 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n24 4.5005
R3134 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n17 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n16 4.5005
R3135 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n20 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n19 4.5005
R3136 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n21 4.30208
R3137 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n29 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n28 3.4105
R3138 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n14 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n13 3.4105
R3139 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n27 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n25 3.13383
R3140 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n0 1.813
R3141 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n4 1.813
R3142 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n2 1.813
R3143 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n7 1.813
R3144 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n10 1.813
R3145 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n20 1.70258
R3146 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n21 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n17 1.43175
R3147 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n3 1.32133
R3148 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n8 1.32133
R3149 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n11 1.32133
R3150 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n12 1.04217
R3151 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n5 0.796333
R3152 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n9 0.771333
R3153 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n1 0.5255
R3154 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n14 0.279652
R3155 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n29 0.236924
R3156 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n28 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n27 0.135917
R3157 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n44 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t7 84.3405
R3158 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n38 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t8 83.2221
R3159 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n34 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t10 83.2221
R3160 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n30 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t6 83.2221
R3161 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n28 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t23 83.2221
R3162 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n32 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t11 83.2221
R3163 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n36 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t17 83.2221
R3164 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n45 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t22 83.2221
R3165 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n42 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t2 83.2221
R3166 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n40 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t0 83.2221
R3167 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n29 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n3 66.665
R3168 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n33 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n2 66.665
R3169 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n37 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n1 66.665
R3170 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n44 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n43 66.665
R3171 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n41 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n0 66.665
R3172 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t20 59.8851
R3173 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t14 55.7878
R3174 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t15 55.5545
R3175 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t21 49.6518
R3176 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n26 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n6 18.1401
R3177 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n26 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n25 16.8247
R3178 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t16 16.5305
R3179 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t3 16.5305
R3180 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t18 16.5305
R3181 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t12 16.5305
R3182 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t5 16.5305
R3183 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t13 16.5305
R3184 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n43 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t4 16.5305
R3185 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n43 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t19 16.5305
R3186 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t1 16.5305
R3187 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t9 16.5305
R3188 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n29 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n28 9.92893
R3189 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n33 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n32 9.92893
R3190 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n37 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n36 9.92893
R3191 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n45 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n44 9.92811
R3192 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n41 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n40 9.92811
R3193 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n27 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n26 7.49008
R3194 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n5 7.44425
R3195 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n4 7.39008
R3196 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 7.00883
R3197 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n31 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n30 6.00467
R3198 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n35 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n34 6.00467
R3199 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n39 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n38 6.00467
R3200 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n46 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n42 6.00467
R3201 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n28 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n27 4.5005
R3202 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n32 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n31 4.5005
R3203 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n36 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n35 4.5005
R3204 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n46 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n45 4.5005
R3205 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n40 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n39 4.5005
R3206 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n16 3.90596
R3207 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n9 3.90547
R3208 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n19 3.4105
R3209 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n24 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n23 3.4105
R3210 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n12 3.4105
R3211 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n42 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n41 1.08427
R3212 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n30 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n29 0.929322
R3213 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n34 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n33 0.929322
R3214 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n38 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n37 0.929322
R3215 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t28 0.523604
R3216 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t40 0.523604
R3217 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t33 0.523604
R3218 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t25 0.523604
R3219 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t43 0.523604
R3220 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n24 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n20 0.495958
R3221 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t26 0.402677
R3222 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t37 0.402677
R3223 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t30 0.402677
R3224 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t42 0.402677
R3225 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t41 0.402677
R3226 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n25 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n24 0.319708
R3227 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t34 0.28175
R3228 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t39 0.28175
R3229 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t27 0.28175
R3230 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t32 0.28175
R3231 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t38 0.28175
R3232 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n22 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t24 0.28175
R3233 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t31 0.28175
R3234 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t36 0.28175
R3235 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t29 0.28175
R3236 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t35 0.28175
R3237 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n7 0.242354
R3238 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n10 0.242354
R3239 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n22 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n21 0.242354
R3240 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n17 0.242354
R3241 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n14 0.242354
R3242 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n25 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n13 0.17724
R3243 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n8 0.121427
R3244 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n11 0.121427
R3245 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n22 0.121427
R3246 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n18 0.121427
R3247 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n15 0.121427
R3248 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n27 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.04425
R3249 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n31 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.04425
R3250 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n35 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.04425
R3251 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n39 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.04425
R3252 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n46 0.04425
R3253 N_IN.n43 N_IN.t2 170.625
R3254 N_IN.n44 N_IN.t4 170.625
R3255 N_IN.n41 N_IN.t16 170.625
R3256 N_IN.n38 N_IN.t36 170.625
R3257 N_IN.n51 N_IN.t21 170.625
R3258 N_IN.n52 N_IN.t8 170.625
R3259 N_IN.n37 N_IN.t12 170.625
R3260 N_IN.n36 N_IN.t14 170.625
R3261 N_IN.n1 N_IN.t1 170.625
R3262 N_IN.n2 N_IN.t19 170.625
R3263 N_IN.n42 N_IN.t20 170.625
R3264 N_IN.n40 N_IN.t11 170.625
R3265 N_IN.n47 N_IN.t30 170.625
R3266 N_IN.n48 N_IN.t18 170.625
R3267 N_IN.n39 N_IN.t27 170.625
R3268 N_IN.n35 N_IN.t6 170.625
R3269 N_IN.n55 N_IN.t24 170.625
R3270 N_IN.n56 N_IN.t26 170.625
R3271 N_IN.n34 N_IN.t33 170.625
R3272 N_IN.n33 N_IN.t23 170.625
R3273 N_IN.n13 N_IN.t37 120.255
R3274 N_IN.n14 N_IN.t38 120.255
R3275 N_IN.n11 N_IN.t9 120.255
R3276 N_IN.n8 N_IN.t31 120.255
R3277 N_IN.n21 N_IN.t17 120.255
R3278 N_IN.n22 N_IN.t0 120.255
R3279 N_IN.n7 N_IN.t5 120.255
R3280 N_IN.n4 N_IN.t7 120.255
R3281 N_IN.n29 N_IN.t34 120.255
R3282 N_IN.n30 N_IN.t13 120.255
R3283 N_IN.n12 N_IN.t35 120.255
R3284 N_IN.n10 N_IN.t29 120.255
R3285 N_IN.n17 N_IN.t22 120.255
R3286 N_IN.n18 N_IN.t32 120.255
R3287 N_IN.n9 N_IN.t15 120.255
R3288 N_IN.n6 N_IN.t28 120.255
R3289 N_IN.n25 N_IN.t3 120.255
R3290 N_IN.n26 N_IN.t10 120.255
R3291 N_IN.n5 N_IN.t25 120.255
R3292 N_IN.n3 N_IN.t39 120.255
R3293 N_IN.n13 N_IN.n12 12.4588
R3294 N_IN.n16 N_IN.n15 10.7088
R3295 N_IN.n20 N_IN.n19 10.7088
R3296 N_IN.n24 N_IN.n23 10.7088
R3297 N_IN.n28 N_IN.n27 10.7088
R3298 N_IN.n32 N_IN.n2 9.62342
R3299 N_IN.n31 N_IN.n3 7.38592
R3300 N_IN.n43 N_IN 7.30883
R3301 N_IN N_IN.n42 6.8505
R3302 N_IN.n46 N_IN 6.24425
R3303 N_IN N_IN.n49 6.24425
R3304 N_IN.n54 N_IN 6.24425
R3305 N_IN N_IN.n57 6.24425
R3306 N_IN.n31 N_IN.n30 6.21508
R3307 N_IN N_IN.n45 6.16508
R3308 N_IN.n50 N_IN 6.16508
R3309 N_IN N_IN.n53 6.16508
R3310 N_IN N_IN.n0 6.16508
R3311 N_IN.n33 N_IN.n32 5.67758
R3312 N_IN.n36 N_IN.n0 1.91925
R3313 N_IN.n53 N_IN.n52 1.91925
R3314 N_IN.n50 N_IN.n38 1.91925
R3315 N_IN.n45 N_IN.n44 1.91925
R3316 N_IN.n28 N_IN.n4 1.91925
R3317 N_IN.n23 N_IN.n22 1.91925
R3318 N_IN.n20 N_IN.n8 1.91925
R3319 N_IN.n15 N_IN.n14 1.91925
R3320 N_IN.n34 N_IN.n33 1.613
R3321 N_IN.n56 N_IN.n55 1.613
R3322 N_IN.n39 N_IN.n35 1.613
R3323 N_IN.n48 N_IN.n47 1.613
R3324 N_IN.n42 N_IN.n40 1.613
R3325 N_IN.n5 N_IN.n3 1.613
R3326 N_IN.n26 N_IN.n25 1.613
R3327 N_IN.n9 N_IN.n6 1.613
R3328 N_IN.n18 N_IN.n17 1.613
R3329 N_IN.n12 N_IN.n10 1.613
R3330 N_IN.n57 N_IN.n56 1.38175
R3331 N_IN.n54 N_IN.n35 1.38175
R3332 N_IN.n49 N_IN.n48 1.38175
R3333 N_IN.n46 N_IN.n40 1.38175
R3334 N_IN.n27 N_IN.n26 1.38175
R3335 N_IN.n24 N_IN.n6 1.38175
R3336 N_IN.n19 N_IN.n18 1.38175
R3337 N_IN.n16 N_IN.n10 1.38175
R3338 N_IN.n1 N_IN.n0 1.14425
R3339 N_IN.n53 N_IN.n37 1.14425
R3340 N_IN.n51 N_IN.n50 1.14425
R3341 N_IN.n45 N_IN.n41 1.14425
R3342 N_IN.n29 N_IN.n28 1.14425
R3343 N_IN.n23 N_IN.n7 1.14425
R3344 N_IN.n21 N_IN.n20 1.14425
R3345 N_IN.n15 N_IN.n11 1.14425
R3346 N_IN.n32 N_IN 0.871333
R3347 N_IN N_IN.n31 0.846333
R3348 N_IN.n57 N_IN.n34 0.60675
R3349 N_IN.n55 N_IN.n54 0.60675
R3350 N_IN.n49 N_IN.n39 0.60675
R3351 N_IN.n47 N_IN.n46 0.60675
R3352 N_IN.n27 N_IN.n5 0.60675
R3353 N_IN.n25 N_IN.n24 0.60675
R3354 N_IN.n19 N_IN.n9 0.60675
R3355 N_IN.n17 N_IN.n16 0.60675
R3356 N_IN.n2 N_IN.n1 0.538
R3357 N_IN.n37 N_IN.n36 0.538
R3358 N_IN.n52 N_IN.n51 0.538
R3359 N_IN.n41 N_IN.n38 0.538
R3360 N_IN.n44 N_IN.n43 0.538
R3361 N_IN.n30 N_IN.n29 0.538
R3362 N_IN.n7 N_IN.n4 0.538
R3363 N_IN.n22 N_IN.n21 0.538
R3364 N_IN.n11 N_IN.n8 0.538
R3365 N_IN.n14 N_IN.n13 0.538
R3366 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t12 93.1806
R3367 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t13 83.2221
R3368 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t8 83.2221
R3369 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t9 83.2221
R3370 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t6 83.2221
R3371 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t4 83.2221
R3372 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t18 83.2221
R3373 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t17 83.2221
R3374 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n25 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t2 83.2221
R3375 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t0 83.2221
R3376 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n19 66.665
R3377 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n24 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n18 66.665
R3378 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n0 66.665
R3379 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n1 66.665
R3380 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n2 66.665
R3381 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t21 55.7445
R3382 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t22 55.4987
R3383 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t23 50.8944
R3384 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t20 49.6614
R3385 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n5 25.8797
R3386 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t14 16.5305
R3387 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t11 16.5305
R3388 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t1 16.5305
R3389 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t3 16.5305
R3390 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t15 16.5305
R3391 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t16 16.5305
R3392 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t10 16.5305
R3393 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t7 16.5305
R3394 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t19 16.5305
R3395 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t5 16.5305
R3396 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n8 9.92893
R3397 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n12 9.92893
R3398 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n16 9.92893
R3399 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n24 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n23 9.92893
R3400 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n3 8.70614
R3401 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n4 7.27133
R3402 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 6.8255
R3403 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n22 6.00467
R3404 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n9 6.00467
R3405 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n13 6.00467
R3406 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n26 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n17 6.00467
R3407 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n22 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n21 4.5005
R3408 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n6 4.5005
R3409 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n10 4.5005
R3410 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n14 4.5005
R3411 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n26 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n25 4.5005
R3412 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n20 1.08427
R3413 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n7 0.929322
R3414 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n11 0.929322
R3415 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n15 0.929322
R3416 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n25 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n24 0.929322
R3417 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n22 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.04425
R3418 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.04425
R3419 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.04425
R3420 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.04425
R3421 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n26 0.04425
R3422 a_n9736_226.n9 a_n9736_226.t1 221.916
R3423 a_n9736_226.n7 a_n9736_226.t2 221.913
R3424 a_n9736_226.n7 a_n9736_226.t3 221.91
R3425 a_n9736_226.t0 a_n9736_226.n9 221.909
R3426 a_n9736_226.n2 a_n9736_226.n1 71.3963
R3427 a_n9736_226.n2 a_n9736_226.n0 71.3963
R3428 a_n9736_226.n5 a_n9736_226.n4 71.3963
R3429 a_n9736_226.n5 a_n9736_226.n3 71.3963
R3430 a_n9736_226.n1 a_n9736_226.t6 16.5305
R3431 a_n9736_226.n1 a_n9736_226.t9 16.5305
R3432 a_n9736_226.n0 a_n9736_226.t11 16.5305
R3433 a_n9736_226.n0 a_n9736_226.t8 16.5305
R3434 a_n9736_226.n4 a_n9736_226.t10 16.5305
R3435 a_n9736_226.n4 a_n9736_226.t7 16.5305
R3436 a_n9736_226.n3 a_n9736_226.t5 16.5305
R3437 a_n9736_226.n3 a_n9736_226.t4 16.5305
R3438 a_n9736_226.n9 a_n9736_226.n8 9.24407
R3439 a_n9736_226.n8 a_n9736_226.n7 7.48275
R3440 a_n9736_226.n8 a_n9736_226.n6 4.33483
R3441 a_n9736_226.n6 a_n9736_226.n2 0.3505
R3442 a_n9736_226.n6 a_n9736_226.n5 0.3505
R3443 opa_folded_cascode_0.VB2.n7 opa_folded_cascode_0.VB2.t12 135.499
R3444 opa_folded_cascode_0.VB2.n8 opa_folded_cascode_0.VB2.t13 135.499
R3445 opa_folded_cascode_0.VB2.n0 opa_folded_cascode_0.VB2.t4 134.734
R3446 opa_folded_cascode_0.VB2.n4 opa_folded_cascode_0.VB2.t6 134.734
R3447 opa_folded_cascode_0.VB2.n4 opa_folded_cascode_0.VB2.t3 134.734
R3448 opa_folded_cascode_0.VB2.n0 opa_folded_cascode_0.VB2.t0 134.734
R3449 opa_folded_cascode_0.VB2.n1 opa_folded_cascode_0.VB2.t1 134.734
R3450 opa_folded_cascode_0.VB2.n1 opa_folded_cascode_0.VB2.t5 134.734
R3451 opa_folded_cascode_0.VB2.n3 opa_folded_cascode_0.VB2.t2 134.734
R3452 opa_folded_cascode_0.VB2.n3 opa_folded_cascode_0.VB2.t7 134.734
R3453 opa_folded_cascode_0.VB2.n7 opa_folded_cascode_0.VB2.t14 134.715
R3454 opa_folded_cascode_0.VB2.n8 opa_folded_cascode_0.VB2.t15 134.715
R3455 opa_folded_cascode_0.VB2.n11 opa_folded_cascode_0.VB2.t8 133.338
R3456 opa_folded_cascode_0.VB2.n10 opa_folded_cascode_0.VB2.t10 132.731
R3457 opa_folded_cascode_0.VB2.n12 opa_folded_cascode_0.VB2.t11 58.9067
R3458 opa_folded_cascode_0.VB2.n11 opa_folded_cascode_0.VB2.t9 58.9067
R3459 opa_folded_cascode_0.VB2.n5 opa_folded_cascode_0.VB2.n3 15.4672
R3460 opa_folded_cascode_0.VB2.n2 opa_folded_cascode_0.VB2.n0 15.4672
R3461 opa_folded_cascode_0.VB2.n9 opa_folded_cascode_0.VB2 9.85842
R3462 opa_folded_cascode_0.VB2.n10 opa_folded_cascode_0.VB2.n9 8.58003
R3463 opa_folded_cascode_0.VB2.n6 opa_folded_cascode_0.VB2.n5 8.3355
R3464 opa_folded_cascode_0.VB2.n6 opa_folded_cascode_0.VB2.n2 7.15195
R3465 opa_folded_cascode_0.VB2 opa_folded_cascode_0.VB2.n7 6.49842
R3466 opa_folded_cascode_0.VB2 opa_folded_cascode_0.VB2.n8 6.33383
R3467 opa_folded_cascode_0.VB2.n5 opa_folded_cascode_0.VB2.n4 4.5005
R3468 opa_folded_cascode_0.VB2.n2 opa_folded_cascode_0.VB2.n1 4.5005
R3469 opa_folded_cascode_0.VB2.n12 opa_folded_cascode_0.VB2.n11 2.09724
R3470 opa_folded_cascode_0.VB2.n9 opa_folded_cascode_0.VB2.n6 1.70389
R3471 opa_folded_cascode_0.VB2 opa_folded_cascode_0.VB2.n12 0.508501
R3472 opa_folded_cascode_0.VB2 opa_folded_cascode_0.VB2.n10 0.0282778
R3473 opa_folded_cascode_0.monticelli_top_0.A.n3 opa_folded_cascode_0.monticelli_top_0.A.t7 168.994
R3474 opa_folded_cascode_0.monticelli_top_0.A.n4 opa_folded_cascode_0.monticelli_top_0.A.t9 168.994
R3475 opa_folded_cascode_0.monticelli_top_0.A.n3 opa_folded_cascode_0.monticelli_top_0.A.t6 168.375
R3476 opa_folded_cascode_0.monticelli_top_0.A.n4 opa_folded_cascode_0.monticelli_top_0.A.t8 168.375
R3477 opa_folded_cascode_0.monticelli_top_0.A.n7 opa_folded_cascode_0.monticelli_top_0.A.t4 69.6491
R3478 opa_folded_cascode_0.monticelli_top_0.A.n1 opa_folded_cascode_0.monticelli_top_0.A.t3 60.3003
R3479 opa_folded_cascode_0.monticelli_top_0.A.n0 opa_folded_cascode_0.monticelli_top_0.A.t1 59.8253
R3480 opa_folded_cascode_0.monticelli_top_0.A.n7 opa_folded_cascode_0.monticelli_top_0.A.t5 59.4176
R3481 opa_folded_cascode_0.monticelli_top_0.A.n2 opa_folded_cascode_0.monticelli_top_0.A.t0 49.8882
R3482 opa_folded_cascode_0.monticelli_top_0.A.n0 opa_folded_cascode_0.monticelli_top_0.A.t2 49.6789
R3483 opa_folded_cascode_0.monticelli_top_0.A.n1 opa_folded_cascode_0.monticelli_top_0.A.n0 12.9172
R3484 opa_folded_cascode_0.monticelli_top_0.A.n6 opa_folded_cascode_0.monticelli_top_0.A.n5 10.0151
R3485 opa_folded_cascode_0.monticelli_top_0.A opa_folded_cascode_0.monticelli_top_0.A.n7 6.413
R3486 opa_folded_cascode_0.monticelli_top_0.A.n2 opa_folded_cascode_0.monticelli_top_0.A.n1 5.5094
R3487 opa_folded_cascode_0.monticelli_top_0.A.n6 opa_folded_cascode_0.monticelli_top_0.A.n2 2.75326
R3488 opa_folded_cascode_0.monticelli_top_0.A.n5 opa_folded_cascode_0.monticelli_top_0.A.n4 1.48383
R3489 opa_folded_cascode_0.monticelli_top_0.A.n5 opa_folded_cascode_0.monticelli_top_0.A.n3 1.47967
R3490 opa_folded_cascode_0.monticelli_top_0.A opa_folded_cascode_0.monticelli_top_0.A.n6 0.8255
R3491 a_n11789_1598.n7 a_n11789_1598.t13 221.913
R3492 a_n11789_1598.t15 a_n11789_1598.n33 221.913
R3493 a_n11789_1598.n33 a_n11789_1598.t8 221.911
R3494 a_n11789_1598.n7 a_n11789_1598.t4 221.911
R3495 a_n11789_1598.n22 a_n11789_1598.t12 221.851
R3496 a_n11789_1598.n23 a_n11789_1598.t14 221.851
R3497 a_n11789_1598.n26 a_n11789_1598.t2 221.851
R3498 a_n11789_1598.n27 a_n11789_1598.t9 221.851
R3499 a_n11789_1598.n30 a_n11789_1598.t6 221.851
R3500 a_n11789_1598.n31 a_n11789_1598.t7 221.851
R3501 a_n11789_1598.n18 a_n11789_1598.t11 221.851
R3502 a_n11789_1598.n17 a_n11789_1598.t3 221.851
R3503 a_n11789_1598.n14 a_n11789_1598.t10 221.851
R3504 a_n11789_1598.n13 a_n11789_1598.t1 221.851
R3505 a_n11789_1598.n10 a_n11789_1598.t5 221.851
R3506 a_n11789_1598.n9 a_n11789_1598.t0 221.851
R3507 a_n11789_1598.n2 a_n11789_1598.n1 71.3963
R3508 a_n11789_1598.n2 a_n11789_1598.n0 71.3963
R3509 a_n11789_1598.n5 a_n11789_1598.n4 71.3963
R3510 a_n11789_1598.n5 a_n11789_1598.n3 71.3963
R3511 a_n11789_1598.n1 a_n11789_1598.t18 16.5305
R3512 a_n11789_1598.n1 a_n11789_1598.t21 16.5305
R3513 a_n11789_1598.n0 a_n11789_1598.t23 16.5305
R3514 a_n11789_1598.n0 a_n11789_1598.t17 16.5305
R3515 a_n11789_1598.n4 a_n11789_1598.t22 16.5305
R3516 a_n11789_1598.n4 a_n11789_1598.t19 16.5305
R3517 a_n11789_1598.n3 a_n11789_1598.t20 16.5305
R3518 a_n11789_1598.n3 a_n11789_1598.t16 16.5305
R3519 a_n11789_1598.n21 a_n11789_1598.n20 6.69433
R3520 a_n11789_1598.n33 a_n11789_1598.n32 5.57739
R3521 a_n11789_1598.n8 a_n11789_1598.n7 5.57739
R3522 a_n11789_1598.n19 a_n11789_1598.n18 5.49597
R3523 a_n11789_1598.n24 a_n11789_1598.n23 5.31889
R3524 a_n11789_1598.n22 a_n11789_1598.n21 5.31889
R3525 a_n11789_1598.n28 a_n11789_1598.n27 5.31889
R3526 a_n11789_1598.n26 a_n11789_1598.n25 5.31889
R3527 a_n11789_1598.n32 a_n11789_1598.n31 5.31889
R3528 a_n11789_1598.n30 a_n11789_1598.n29 5.31889
R3529 a_n11789_1598.n17 a_n11789_1598.n16 5.31889
R3530 a_n11789_1598.n15 a_n11789_1598.n14 5.31889
R3531 a_n11789_1598.n13 a_n11789_1598.n12 5.31889
R3532 a_n11789_1598.n11 a_n11789_1598.n10 5.31889
R3533 a_n11789_1598.n9 a_n11789_1598.n8 5.31889
R3534 a_n11789_1598.n20 a_n11789_1598.n6 4.0215
R3535 a_n11789_1598.n20 a_n11789_1598.n19 3.4105
R3536 a_n11789_1598.n12 a_n11789_1598.n11 2.888
R3537 a_n11789_1598.n16 a_n11789_1598.n15 2.888
R3538 a_n11789_1598.n29 a_n11789_1598.n28 2.888
R3539 a_n11789_1598.n25 a_n11789_1598.n24 2.888
R3540 a_n11789_1598.n6 a_n11789_1598.n2 0.3505
R3541 a_n11789_1598.n6 a_n11789_1598.n5 0.3505
R3542 a_n11789_1598.n11 a_n11789_1598.n8 0.246333
R3543 a_n11789_1598.n15 a_n11789_1598.n12 0.246333
R3544 a_n11789_1598.n32 a_n11789_1598.n29 0.246333
R3545 a_n11789_1598.n28 a_n11789_1598.n25 0.246333
R3546 a_n11789_1598.n24 a_n11789_1598.n21 0.246333
R3547 a_n11789_1598.n23 a_n11789_1598.n22 0.123417
R3548 a_n11789_1598.n27 a_n11789_1598.n26 0.123417
R3549 a_n11789_1598.n31 a_n11789_1598.n30 0.123417
R3550 a_n11789_1598.n18 a_n11789_1598.n17 0.123417
R3551 a_n11789_1598.n14 a_n11789_1598.n13 0.123417
R3552 a_n11789_1598.n10 a_n11789_1598.n9 0.123417
R3553 a_n11789_1598.n19 a_n11789_1598.n16 0.06925
R3554 P_IN[2].n0 P_IN[2].t7 172.237
R3555 P_IN[2].n5 P_IN[2].t4 171.161
R3556 P_IN[2].n0 P_IN[2].t3 170.625
R3557 P_IN[2].n5 P_IN[2].t5 170.625
R3558 P_IN[2].n2 P_IN[2].t6 121.868
R3559 P_IN[2].n1 P_IN[2].t0 120.793
R3560 P_IN[2].n2 P_IN[2].t1 120.255
R3561 P_IN[2].n1 P_IN[2].t2 120.255
R3562 P_IN[2].n4 P_IN[2] 11.763
R3563 P_IN[2].n3 P_IN[2].n1 7.53592
R3564 P_IN[2] P_IN[2].n0 7.138
R3565 P_IN[2].n6 P_IN[2].n5 5.82758
R3566 P_IN[2].n3 P_IN[2].n2 5.29008
R3567 P_IN[2] P_IN[2].n6 1.56092
R3568 P_IN[2].n6 P_IN[2].n4 0.9505
R3569 P_IN[2].n4 P_IN[2].n3 0.767167
R3570 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t6 151.438
R3571 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t7 149.923
R3572 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n2 79.7972
R3573 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n0 79.7972
R3574 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n1 79.7972
R3575 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n7 79.6389
R3576 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t9 9.23217
R3577 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t1 9.23217
R3578 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t3 9.23217
R3579 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t8 9.23217
R3580 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t5 9.23217
R3581 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t2 9.23217
R3582 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t0 9.23217
R3583 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t4 9.23217
R3584 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n4 4.75071
R3585 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n5 0.429667
R3586 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n3 0.429667
R3587 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n6 0.158833
R3588 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t22 94.3966
R3589 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t19 84.4381
R3590 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t15 84.4381
R3591 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t18 84.4381
R3592 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t7 84.4381
R3593 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t13 84.4381
R3594 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t4 84.4381
R3595 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t6 84.4381
R3596 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t9 84.4381
R3597 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t10 84.4381
R3598 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n4 75.1793
R3599 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n3 75.1793
R3600 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n2 75.1793
R3601 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n1 75.1793
R3602 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n0 75.1793
R3603 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n25 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t0 65.725
R3604 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t1 65.2617
R3605 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n22 50.0985
R3606 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n21 49.0864
R3607 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n24 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n20 49.0864
R3608 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n18 24.7318
R3609 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n25 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n24 17.6109
R3610 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n6 10.5047
R3611 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n9 10.5047
R3612 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n12 10.5047
R3613 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n15 10.5047
R3614 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t2 10.3318
R3615 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t24 10.3318
R3616 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n22 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t27 10.3318
R3617 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n22 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t26 10.3318
R3618 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t23 10.3318
R3619 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t25 10.3318
R3620 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n24 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n23 10.2127
R3621 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n7 9.92811
R3622 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n10 9.92811
R3623 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n13 9.92811
R3624 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n16 9.92811
R3625 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t20 9.23217
R3626 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t21 9.23217
R3627 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t17 9.23217
R3628 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t8 9.23217
R3629 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t16 9.23217
R3630 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t14 9.23217
R3631 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t3 9.23217
R3632 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t5 9.23217
R3633 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t11 9.23217
R3634 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t12 9.23217
R3635 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n25 5.913
R3636 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n19 5.67967
R3637 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n5 0.896768
R3638 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n8 0.896768
R3639 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n11 0.896768
R3640 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n14 0.896768
R3641 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n17 0.896768
R3642 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.188
R3643 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.188
R3644 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.188
R3645 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.188
R3646 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.188
R3647 P_IN[4].n0 P_IN[4].t4 172.237
R3648 P_IN[4].n5 P_IN[4].t2 171.161
R3649 P_IN[4].n0 P_IN[4].t0 170.625
R3650 P_IN[4].n5 P_IN[4].t1 170.625
R3651 P_IN[4].n2 P_IN[4].t3 121.868
R3652 P_IN[4].n1 P_IN[4].t7 120.793
R3653 P_IN[4].n2 P_IN[4].t5 120.255
R3654 P_IN[4].n1 P_IN[4].t6 120.255
R3655 P_IN[4].n3 P_IN[4].n1 7.53592
R3656 P_IN[4] P_IN[4].n0 7.138
R3657 P_IN[4].n6 P_IN[4].n5 5.82758
R3658 P_IN[4].n3 P_IN[4].n2 5.29008
R3659 P_IN[4].n4 P_IN[4] 4.563
R3660 P_IN[4] P_IN[4].n6 1.56092
R3661 P_IN[4].n6 P_IN[4].n4 1.31717
R3662 P_IN[4].n4 P_IN[4].n3 0.4005
R3663 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t20 142.597
R3664 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t8 141.03
R3665 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t19 139.588
R3666 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t23 139.588
R3667 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t15 134.712
R3668 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t14 134.712
R3669 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t13 134.712
R3670 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t22 134.712
R3671 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t21 134.712
R3672 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t17 134.712
R3673 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t18 134.712
R3674 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t9 134.712
R3675 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t12 134.712
R3676 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n14 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t11 134.712
R3677 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t16 134.712
R3678 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t10 134.712
R3679 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n19 79.7972
R3680 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n1 79.7972
R3681 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n0 79.7972
R3682 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n21 79.6389
R3683 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t0 9.23217
R3684 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n19 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t6 9.23217
R3685 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t2 9.23217
R3686 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t4 9.23217
R3687 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t5 9.23217
R3688 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t1 9.23217
R3689 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t7 9.23217
R3690 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n21 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t3 9.23217
R3691 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n4 7.83383
R3692 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n13 7.83383
R3693 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n17 5.12671
R3694 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n7 4.61407
R3695 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n5 4.61407
R3696 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n3 4.61407
R3697 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n12 4.61407
R3698 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n15 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n14 4.61407
R3699 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n10 4.61407
R3700 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n9 3.97054
R3701 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n16 3.45425
R3702 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n6 3.13383
R3703 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n11 3.13383
R3704 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n16 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n15 3.01092
R3705 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n8 1.44425
R3706 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n18 0.429667
R3707 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n18 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n2 0.429667
R3708 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n20 0.158833
R3709 a_n4822_n1462.n1 a_n4822_n1462.t0 213.52
R3710 a_n4822_n1462.n2 a_n4822_n1462.t2 213.52
R3711 a_n4822_n1462.n1 a_n4822_n1462.n0 42.5016
R3712 a_n4822_n1462.n3 a_n4822_n1462.n2 42.5016
R3713 a_n4822_n1462.n2 a_n4822_n1462.n1 11.7539
R3714 a_n4822_n1462.n0 a_n4822_n1462.t4 5.77029
R3715 a_n4822_n1462.n0 a_n4822_n1462.t1 5.77029
R3716 a_n4822_n1462.t3 a_n4822_n1462.n3 5.77029
R3717 a_n4822_n1462.n3 a_n4822_n1462.t5 5.77029
R3718 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t5 227.827
R3719 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t4 227.827
R3720 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t3 227.827
R3721 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t0 227.827
R3722 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t7 226.506
R3723 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t2 226.506
R3724 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t6 226.506
R3725 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t1 226.506
R3726 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t12 221.911
R3727 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t15 221.911
R3728 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t14 221.911
R3729 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t8 221.911
R3730 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t10 221.911
R3731 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t13 221.911
R3732 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t9 221.911
R3733 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t11 221.911
R3734 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n11 8.30397
R3735 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n7 6.99147
R3736 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n8 6.73731
R3737 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n10 5.4248
R3738 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n2 4.30208
R3739 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n9 4.05141
R3740 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n12 3.4105
R3741 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n5 3.4105
R3742 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n1 3.12967
R3743 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n3 1.81717
R3744 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n4 1.563
R3745 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n6 0.655651
R3746 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n13 0.362258
R3747 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n0 0.2505
R3748 opa_folded_cascode_0.monticelli_top_0.Bx.n3 opa_folded_cascode_0.monticelli_top_0.Bx.t10 135.254
R3749 opa_folded_cascode_0.monticelli_top_0.Bx.n1 opa_folded_cascode_0.monticelli_top_0.Bx.t12 135.254
R3750 opa_folded_cascode_0.monticelli_top_0.Bx.n8 opa_folded_cascode_0.monticelli_top_0.Bx.t7 135.254
R3751 opa_folded_cascode_0.monticelli_top_0.Bx.n6 opa_folded_cascode_0.monticelli_top_0.Bx.t9 135.254
R3752 opa_folded_cascode_0.monticelli_top_0.Bx.n3 opa_folded_cascode_0.monticelli_top_0.Bx.t6 134.715
R3753 opa_folded_cascode_0.monticelli_top_0.Bx.n4 opa_folded_cascode_0.monticelli_top_0.Bx.t16 134.715
R3754 opa_folded_cascode_0.monticelli_top_0.Bx.n2 opa_folded_cascode_0.monticelli_top_0.Bx.t14 134.715
R3755 opa_folded_cascode_0.monticelli_top_0.Bx.n1 opa_folded_cascode_0.monticelli_top_0.Bx.t11 134.715
R3756 opa_folded_cascode_0.monticelli_top_0.Bx.n8 opa_folded_cascode_0.monticelli_top_0.Bx.t17 134.715
R3757 opa_folded_cascode_0.monticelli_top_0.Bx.n9 opa_folded_cascode_0.monticelli_top_0.Bx.t15 134.715
R3758 opa_folded_cascode_0.monticelli_top_0.Bx.n7 opa_folded_cascode_0.monticelli_top_0.Bx.t13 134.715
R3759 opa_folded_cascode_0.monticelli_top_0.Bx.n6 opa_folded_cascode_0.monticelli_top_0.Bx.t8 134.715
R3760 opa_folded_cascode_0.monticelli_top_0.Bx.n14 opa_folded_cascode_0.monticelli_top_0.Bx.t4 69.7645
R3761 opa_folded_cascode_0.monticelli_top_0.Bx.n11 opa_folded_cascode_0.monticelli_top_0.Bx.t1 60.5923
R3762 opa_folded_cascode_0.monticelli_top_0.Bx.n13 opa_folded_cascode_0.monticelli_top_0.Bx.t5 59.8932
R3763 opa_folded_cascode_0.monticelli_top_0.Bx.n0 opa_folded_cascode_0.monticelli_top_0.Bx.t2 59.8572
R3764 opa_folded_cascode_0.monticelli_top_0.Bx.n11 opa_folded_cascode_0.monticelli_top_0.Bx.t0 59.4447
R3765 opa_folded_cascode_0.monticelli_top_0.Bx.n0 opa_folded_cascode_0.monticelli_top_0.Bx.t3 49.6789
R3766 opa_folded_cascode_0.monticelli_top_0.Bx opa_folded_cascode_0.monticelli_top_0.Bx.n0 15.0818
R3767 opa_folded_cascode_0.monticelli_top_0.Bx.n14 opa_folded_cascode_0.monticelli_top_0.Bx.n13 12.9172
R3768 opa_folded_cascode_0.monticelli_top_0.Bx.n12 opa_folded_cascode_0.monticelli_top_0.Bx.n11 9.36508
R3769 opa_folded_cascode_0.monticelli_top_0.Bx.n12 opa_folded_cascode_0.monticelli_top_0.Bx.n10 7.19425
R3770 opa_folded_cascode_0.monticelli_top_0.Bx opa_folded_cascode_0.monticelli_top_0.Bx.n14 3.55675
R3771 opa_folded_cascode_0.monticelli_top_0.Bx.n13 opa_folded_cascode_0.monticelli_top_0.Bx.n12 2.72758
R3772 opa_folded_cascode_0.monticelli_top_0.Bx.n10 opa_folded_cascode_0.monticelli_top_0.Bx.n5 1.9005
R3773 opa_folded_cascode_0.monticelli_top_0.Bx.n2 opa_folded_cascode_0.monticelli_top_0.Bx.n1 0.538
R3774 opa_folded_cascode_0.monticelli_top_0.Bx.n4 opa_folded_cascode_0.monticelli_top_0.Bx.n3 0.538
R3775 opa_folded_cascode_0.monticelli_top_0.Bx.n7 opa_folded_cascode_0.monticelli_top_0.Bx.n6 0.538
R3776 opa_folded_cascode_0.monticelli_top_0.Bx.n9 opa_folded_cascode_0.monticelli_top_0.Bx.n8 0.538
R3777 opa_folded_cascode_0.monticelli_top_0.Bx.n5 opa_folded_cascode_0.monticelli_top_0.Bx.n2 0.26925
R3778 opa_folded_cascode_0.monticelli_top_0.Bx.n5 opa_folded_cascode_0.monticelli_top_0.Bx.n4 0.26925
R3779 opa_folded_cascode_0.monticelli_top_0.Bx.n10 opa_folded_cascode_0.monticelli_top_0.Bx.n7 0.26925
R3780 opa_folded_cascode_0.monticelli_top_0.Bx.n10 opa_folded_cascode_0.monticelli_top_0.Bx.n9 0.26925
R3781 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t4 227.707
R3782 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t7 227.707
R3783 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t2 227.707
R3784 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t0 227.707
R3785 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t3 226.386
R3786 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t6 226.386
R3787 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t5 226.386
R3788 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t1 226.386
R3789 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t15 221.911
R3790 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t10 221.911
R3791 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t9 221.911
R3792 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t12 221.911
R3793 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t11 221.911
R3794 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t14 221.911
R3795 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t13 221.911
R3796 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t8 221.911
R3797 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n7 9.59425
R3798 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n11 8.80675
R3799 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n10 8.02758
R3800 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n8 7.24008
R3801 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n3 4.43383
R3802 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n2 4.17674
R3803 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n9 3.92608
R3804 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n1 3.64633
R3805 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n12 3.4105
R3806 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n5 3.4105
R3807 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n0 2.86717
R3808 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n4 2.07967
R3809 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n6 0.718318
R3810 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n13 0.424924
R3811 P_IN[1].n0 P_IN[1].t5 172.237
R3812 P_IN[1].n5 P_IN[1].t7 171.161
R3813 P_IN[1].n0 P_IN[1].t4 170.625
R3814 P_IN[1].n5 P_IN[1].t6 170.625
R3815 P_IN[1].n2 P_IN[1].t3 121.868
R3816 P_IN[1].n1 P_IN[1].t2 120.793
R3817 P_IN[1].n2 P_IN[1].t0 120.255
R3818 P_IN[1].n1 P_IN[1].t1 120.255
R3819 P_IN[1].n4 P_IN[1] 15.363
R3820 P_IN[1].n3 P_IN[1].n1 7.53592
R3821 P_IN[1] P_IN[1].n0 7.138
R3822 P_IN[1].n6 P_IN[1].n5 5.82758
R3823 P_IN[1].n3 P_IN[1].n2 5.29008
R3824 P_IN[1] P_IN[1].n6 1.56092
R3825 P_IN[1].n4 P_IN[1].n3 0.9505
R3826 P_IN[1].n6 P_IN[1].n4 0.767167
R3827 a_n9242_n890.n7 a_n9242_n890.t1 236.924
R3828 a_n9242_n890.t0 a_n9242_n890.n7 235.214
R3829 a_n9242_n890.n2 a_n9242_n890.n1 71.3963
R3830 a_n9242_n890.n2 a_n9242_n890.n0 71.3963
R3831 a_n9242_n890.n5 a_n9242_n890.n4 71.3963
R3832 a_n9242_n890.n5 a_n9242_n890.n3 71.3963
R3833 a_n9242_n890.n1 a_n9242_n890.t8 16.5305
R3834 a_n9242_n890.n1 a_n9242_n890.t5 16.5305
R3835 a_n9242_n890.n0 a_n9242_n890.t2 16.5305
R3836 a_n9242_n890.n0 a_n9242_n890.t7 16.5305
R3837 a_n9242_n890.n4 a_n9242_n890.t4 16.5305
R3838 a_n9242_n890.n4 a_n9242_n890.t9 16.5305
R3839 a_n9242_n890.n3 a_n9242_n890.t6 16.5305
R3840 a_n9242_n890.n3 a_n9242_n890.t3 16.5305
R3841 a_n9242_n890.n7 a_n9242_n890.n6 4.7735
R3842 a_n9242_n890.n6 a_n9242_n890.n2 0.3505
R3843 a_n9242_n890.n6 a_n9242_n890.n5 0.3505
R3844 P_IN[0].n0 P_IN[0].t0 172.237
R3845 P_IN[0].n5 P_IN[0].t5 171.161
R3846 P_IN[0].n0 P_IN[0].t4 170.625
R3847 P_IN[0].n5 P_IN[0].t2 170.625
R3848 P_IN[0].n2 P_IN[0].t7 121.868
R3849 P_IN[0].n1 P_IN[0].t1 120.793
R3850 P_IN[0].n2 P_IN[0].t3 120.255
R3851 P_IN[0].n1 P_IN[0].t6 120.255
R3852 P_IN[0].n4 P_IN[0] 18.963
R3853 P_IN[0].n3 P_IN[0].n1 7.53592
R3854 P_IN[0] P_IN[0].n0 7.138
R3855 P_IN[0].n6 P_IN[0].n5 5.82758
R3856 P_IN[0].n3 P_IN[0].n2 5.29008
R3857 P_IN[0] P_IN[0].n6 1.56092
R3858 P_IN[0].n4 P_IN[0].n3 1.13383
R3859 P_IN[0].n6 P_IN[0].n4 0.583833
R3860 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t15 140.945
R3861 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t13 140.945
R3862 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t11 140.945
R3863 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t12 140.945
R3864 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n11 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t14 139.635
R3865 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t9 139.635
R3866 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n10 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t8 139.625
R3867 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n8 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t10 139.625
R3868 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t6 134.712
R3869 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t4 134.712
R3870 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t3 134.712
R3871 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t2 134.712
R3872 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t1 134.712
R3873 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t5 134.712
R3874 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t0 134.712
R3875 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t7 134.712
R3876 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n0 11.8254
R3877 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n3 10.2587
R3878 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n4 9.9879
R3879 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n1 8.42123
R3880 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n10 6.5255
R3881 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n7 4.95883
R3882 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n9 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n8 4.688
R3883 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n9 4.42741
R3884 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n2 4.14826
R3885 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n13 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n12 3.4105
R3886 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n6 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n5 3.4105
R3887 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n12 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n11 3.12133
R3888 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n13 0.675591
R3889 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n6 0.453409
R3890 opa_folded_cascode_0.monticelli_top_0.Ax.n1 opa_folded_cascode_0.monticelli_top_0.Ax.t9 217.037
R3891 opa_folded_cascode_0.monticelli_top_0.Ax.n0 opa_folded_cascode_0.monticelli_top_0.Ax.t8 217.037
R3892 opa_folded_cascode_0.monticelli_top_0.Ax.n1 opa_folded_cascode_0.monticelli_top_0.Ax.t7 211.755
R3893 opa_folded_cascode_0.monticelli_top_0.Ax.n0 opa_folded_cascode_0.monticelli_top_0.Ax.t6 211.755
R3894 opa_folded_cascode_0.monticelli_top_0.Ax.n7 opa_folded_cascode_0.monticelli_top_0.Ax.t5 60.6506
R3895 opa_folded_cascode_0.monticelli_top_0.Ax.n5 opa_folded_cascode_0.monticelli_top_0.Ax.t0 60.0612
R3896 opa_folded_cascode_0.monticelli_top_0.Ax.n7 opa_folded_cascode_0.monticelli_top_0.Ax.t4 59.4176
R3897 opa_folded_cascode_0.monticelli_top_0.Ax.n3 opa_folded_cascode_0.monticelli_top_0.Ax.t2 51.0085
R3898 opa_folded_cascode_0.monticelli_top_0.Ax.n6 opa_folded_cascode_0.monticelli_top_0.Ax.t1 50.7632
R3899 opa_folded_cascode_0.monticelli_top_0.Ax.n3 opa_folded_cascode_0.monticelli_top_0.Ax.t3 49.6518
R3900 opa_folded_cascode_0.monticelli_top_0.Ax.n4 opa_folded_cascode_0.monticelli_top_0.Ax.n2 12.2317
R3901 opa_folded_cascode_0.monticelli_top_0.Ax.n2 opa_folded_cascode_0.monticelli_top_0.Ax.n0 5.26748
R3902 opa_folded_cascode_0.monticelli_top_0.Ax.n6 opa_folded_cascode_0.monticelli_top_0.Ax.n5 5.03383
R3903 opa_folded_cascode_0.monticelli_top_0.Ax.n5 opa_folded_cascode_0.monticelli_top_0.Ax.n4 4.99626
R3904 opa_folded_cascode_0.monticelli_top_0.Ax opa_folded_cascode_0.monticelli_top_0.Ax.n7 4.92133
R3905 opa_folded_cascode_0.monticelli_top_0.Ax opa_folded_cascode_0.monticelli_top_0.Ax.n6 3.04842
R3906 opa_folded_cascode_0.monticelli_top_0.Ax.n2 opa_folded_cascode_0.monticelli_top_0.Ax.n1 0.565401
R3907 opa_folded_cascode_0.monticelli_top_0.Ax.n4 opa_folded_cascode_0.monticelli_top_0.Ax.n3 0.338
R3908 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t6 134.734
R3909 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t5 134.734
R3910 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t7 134.734
R3911 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t4 134.734
R3912 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n2 79.7972
R3913 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n0 79.7972
R3914 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n1 79.7972
R3915 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n9 79.6389
R3916 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n4 11.8125
R3917 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t9 9.23217
R3918 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t0 9.23217
R3919 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t1 9.23217
R3920 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t11 9.23217
R3921 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t8 9.23217
R3922 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t2 9.23217
R3923 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t3 9.23217
R3924 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.t10 9.23217
R3925 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n5 8.03342
R3926 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n6 5.19579
R3927 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n7 0.429667
R3928 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n3 0.429667
R3929 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD.n8 0.158833
R3930 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t0 228.496
R3931 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t3 228.496
R3932 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t2 227.538
R3933 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t1 227.538
R3934 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t5 221.974
R3935 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t4 221.974
R3936 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t7 221.851
R3937 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t6 221.851
R3938 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n4 9.92404
R3939 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n3 9.90278
R3940 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n0 6.28466
R3941 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n1 4.10425
R3942 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n2 0.404985
R3943 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n5 0.299591
R3944 a_n10488_226.n15 a_n10488_226.t3 221.913
R3945 a_n10488_226.n0 a_n10488_226.t1 221.913
R3946 a_n10488_226.n8 a_n10488_226.t5 221.913
R3947 a_n10488_226.n0 a_n10488_226.t4 221.911
R3948 a_n10488_226.n8 a_n10488_226.t0 221.911
R3949 a_n10488_226.t7 a_n10488_226.n15 221.911
R3950 a_n10488_226.n11 a_n10488_226.t6 221.851
R3951 a_n10488_226.n10 a_n10488_226.t2 221.851
R3952 a_n10488_226.n3 a_n10488_226.n2 71.3963
R3953 a_n10488_226.n3 a_n10488_226.n1 71.3963
R3954 a_n10488_226.n6 a_n10488_226.n5 71.3963
R3955 a_n10488_226.n6 a_n10488_226.n4 71.3963
R3956 a_n10488_226.n2 a_n10488_226.t14 16.5305
R3957 a_n10488_226.n2 a_n10488_226.t10 16.5305
R3958 a_n10488_226.n1 a_n10488_226.t8 16.5305
R3959 a_n10488_226.n1 a_n10488_226.t12 16.5305
R3960 a_n10488_226.n5 a_n10488_226.t15 16.5305
R3961 a_n10488_226.n5 a_n10488_226.t13 16.5305
R3962 a_n10488_226.n4 a_n10488_226.t11 16.5305
R3963 a_n10488_226.n4 a_n10488_226.t9 16.5305
R3964 a_n10488_226.n9 a_n10488_226.n8 6.97216
R3965 a_n10488_226.n15 a_n10488_226.n14 5.78883
R3966 a_n10488_226.n10 a_n10488_226.n9 4.97106
R3967 a_n10488_226.n12 a_n10488_226.n11 4.97106
R3968 a_n10488_226.n13 a_n10488_226.n12 4.69233
R3969 a_n10488_226.n13 a_n10488_226.n7 4.3975
R3970 a_n10488_226.n14 a_n10488_226.n0 3.69924
R3971 a_n10488_226.n14 a_n10488_226.n13 3.4105
R3972 a_n10488_226.n7 a_n10488_226.n3 0.3505
R3973 a_n10488_226.n7 a_n10488_226.n6 0.3505
R3974 a_n10488_226.n12 a_n10488_226.n9 0.246333
R3975 a_n10488_226.n11 a_n10488_226.n10 0.123417
R3976 opa_folded_cascode_0.VB1.n5 opa_folded_cascode_0.VB1.t1 221.913
R3977 opa_folded_cascode_0.VB1.n10 opa_folded_cascode_0.VB1.t2 221.913
R3978 opa_folded_cascode_0.VB1.n5 opa_folded_cascode_0.VB1.t5 221.911
R3979 opa_folded_cascode_0.VB1.n10 opa_folded_cascode_0.VB1.t6 221.911
R3980 opa_folded_cascode_0.VB1.n8 opa_folded_cascode_0.VB1.t3 221.851
R3981 opa_folded_cascode_0.VB1.n12 opa_folded_cascode_0.VB1.t4 221.851
R3982 opa_folded_cascode_0.VB1.n13 opa_folded_cascode_0.VB1.t0 221.851
R3983 opa_folded_cascode_0.VB1.n7 opa_folded_cascode_0.VB1.t7 221.851
R3984 opa_folded_cascode_0.VB1.n0 opa_folded_cascode_0.VB1.t15 214.787
R3985 opa_folded_cascode_0.VB1.n1 opa_folded_cascode_0.VB1.t12 214.787
R3986 opa_folded_cascode_0.VB1.n0 opa_folded_cascode_0.VB1.t13 214.005
R3987 opa_folded_cascode_0.VB1.n1 opa_folded_cascode_0.VB1.t14 214.005
R3988 opa_folded_cascode_0.VB1.n3 opa_folded_cascode_0.VB1.t10 212.323
R3989 opa_folded_cascode_0.VB1.n18 opa_folded_cascode_0.VB1.t8 212.106
R3990 opa_folded_cascode_0.VB1.n4 opa_folded_cascode_0.VB1.t11 48.2714
R3991 opa_folded_cascode_0.VB1.n17 opa_folded_cascode_0.VB1.t9 48.2714
R3992 opa_folded_cascode_0.VB1.n3 opa_folded_cascode_0.VB1.n2 17.7367
R3993 opa_folded_cascode_0.VB1.n11 opa_folded_cascode_0.VB1.n10 9.98379
R3994 opa_folded_cascode_0.VB1.n6 opa_folded_cascode_0.VB1.n5 9.98379
R3995 opa_folded_cascode_0.VB1.n16 opa_folded_cascode_0.VB1.n15 9.65976
R3996 opa_folded_cascode_0.VB1.n15 opa_folded_cascode_0.VB1.n9 8.23783
R3997 opa_folded_cascode_0.VB1.n2 opa_folded_cascode_0.VB1.n0 7.77967
R3998 opa_folded_cascode_0.VB1 opa_folded_cascode_0.VB1.n1 7.65675
R3999 opa_folded_cascode_0.VB1.n15 opa_folded_cascode_0.VB1.n14 5.65425
R4000 opa_folded_cascode_0.VB1.n7 opa_folded_cascode_0.VB1.n6 4.73193
R4001 opa_folded_cascode_0.VB1.n14 opa_folded_cascode_0.VB1.n13 4.73193
R4002 opa_folded_cascode_0.VB1.n12 opa_folded_cascode_0.VB1.n11 4.73193
R4003 opa_folded_cascode_0.VB1.n9 opa_folded_cascode_0.VB1.n8 4.73193
R4004 opa_folded_cascode_0.VB1.n16 opa_folded_cascode_0.VB1.n4 2.42885
R4005 opa_folded_cascode_0.VB1.n18 opa_folded_cascode_0.VB1.n17 1.41626
R4006 opa_folded_cascode_0.VB1.n17 opa_folded_cascode_0.VB1.n16 1.40802
R4007 opa_folded_cascode_0.VB1.n4 opa_folded_cascode_0.VB1.n3 1.09089
R4008 opa_folded_cascode_0.VB1.n14 opa_folded_cascode_0.VB1.n11 0.246333
R4009 opa_folded_cascode_0.VB1.n9 opa_folded_cascode_0.VB1.n6 0.246333
R4010 opa_folded_cascode_0.VB1.n13 opa_folded_cascode_0.VB1.n12 0.123417
R4011 opa_folded_cascode_0.VB1.n8 opa_folded_cascode_0.VB1.n7 0.123417
R4012 opa_folded_cascode_0.VB1.n2 opa_folded_cascode_0.VB1 0.0734167
R4013 opa_folded_cascode_0.VB1 opa_folded_cascode_0.VB1.n18 0.063
R4014 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t9 147.899
R4015 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t8 146.752
R4016 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n5 79.7972
R4017 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n1 79.7972
R4018 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n0 79.7972
R4019 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n7 79.6389
R4020 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t2 9.23217
R4021 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t6 9.23217
R4022 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t1 9.23217
R4023 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t5 9.23217
R4024 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t4 9.23217
R4025 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t0 9.23217
R4026 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t7 9.23217
R4027 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t3 9.23217
R4028 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n3 4.68805
R4029 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n4 0.429667
R4030 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n2 0.429667
R4031 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n6 0.158833
R4032 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t2 146.321
R4033 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t3 144.415
R4034 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t1 143.702
R4035 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t0 143.431
R4036 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n0 0.390742
R4037 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n1 0.362258
R4038 P_IN[3].n0 P_IN[3].t7 172.237
R4039 P_IN[3].n5 P_IN[3].t1 171.161
R4040 P_IN[3].n0 P_IN[3].t3 170.625
R4041 P_IN[3].n5 P_IN[3].t4 170.625
R4042 P_IN[3].n2 P_IN[3].t6 121.868
R4043 P_IN[3].n1 P_IN[3].t5 120.793
R4044 P_IN[3].n2 P_IN[3].t2 120.255
R4045 P_IN[3].n1 P_IN[3].t0 120.255
R4046 P_IN[3].n4 P_IN[3] 8.163
R4047 P_IN[3].n3 P_IN[3].n1 7.53592
R4048 P_IN[3] P_IN[3].n0 7.138
R4049 P_IN[3].n6 P_IN[3].n5 5.82758
R4050 P_IN[3].n3 P_IN[3].n2 5.29008
R4051 P_IN[3] P_IN[3].n6 1.56092
R4052 P_IN[3].n6 P_IN[3].n4 1.13383
R4053 P_IN[3].n4 P_IN[3].n3 0.583833
R4054 a_n4822_464.n2 a_n4822_464.t2 133.338
R4055 a_n4822_464.n1 a_n4822_464.t0 133.338
R4056 a_n4822_464.n1 a_n4822_464.n0 48.5755
R4057 a_n4822_464.n3 a_n4822_464.n2 48.5755
R4058 a_n4822_464.n0 a_n4822_464.t1 10.3318
R4059 a_n4822_464.n0 a_n4822_464.t5 10.3318
R4060 a_n4822_464.n3 a_n4822_464.t4 10.3318
R4061 a_n4822_464.t3 a_n4822_464.n3 10.3318
R4062 a_n4822_464.n2 a_n4822_464.n1 10.0148
R4063 ROUT.n1 ROUT.t1 160.632
R4064 ROUT.n1 ROUT.t3 134.811
R4065 ROUT.n2 ROUT.t0 16.8154
R4066 ROUT.n0 ROUT.t4 16.8154
R4067 ROUT.n4 ROUT.n0 12.0038
R4068 ROUT.n3 ROUT.n2 6.5267
R4069 ROUT.n2 ROUT.t5 5.78822
R4070 ROUT.n0 ROUT.t2 5.78822
R4071 ROUT.n4 ROUT.n3 5.72758
R4072 ROUT.n3 ROUT 3.44682
R4073 ROUT.n4 ROUT.n1 0.965083
R4074 ROUT ROUT.n4 0.063
R4075 a_n7784_12197.n1 a_n7784_12197.n0 243.671
R4076 a_n7784_12197.n0 a_n7784_12197.t2 15.3866
R4077 a_n7784_12197.n0 a_n7784_12197.t1 15.3866
R4078 a_n7784_12197.t0 a_n7784_12197.n1 15.3866
R4079 a_n7784_12197.n1 a_n7784_12197.t3 15.3866
R4080 a_n11843_11539.n5 a_n11843_11539.t1 160.791
R4081 a_n11843_11539.n0 a_n11843_11539.t4 154.608
R4082 a_n11843_11539.n0 a_n11843_11539.t5 134.811
R4083 a_n11843_11539.t3 a_n11843_11539.n5 134.811
R4084 a_n11843_11539.n3 a_n11843_11539.t6 16.8154
R4085 a_n11843_11539.n1 a_n11843_11539.t0 16.8154
R4086 a_n11843_11539.n4 a_n11843_11539.n3 12.0038
R4087 a_n11843_11539.n2 a_n11843_11539.n0 6.72342
R4088 a_n11843_11539.n2 a_n11843_11539.n1 6.5892
R4089 a_n11843_11539.n3 a_n11843_11539.t2 5.78822
R4090 a_n11843_11539.n1 a_n11843_11539.t7 5.78822
R4091 a_n11843_11539.n4 a_n11843_11539.n2 5.66508
R4092 a_n11843_11539.n5 a_n11843_11539.n4 0.965083
R4093 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t5 141.129
R4094 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t4 141.129
R4095 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t6 139.808
R4096 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t7 139.808
R4097 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t2 134.732
R4098 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t1 134.732
R4099 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t0 134.732
R4100 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t3 134.732
R4101 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n1 9.87092
R4102 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n0 9.44517
R4103 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n3 5.85274
R4104 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n5 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n4 3.923
R4105 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n2 0.641409
R4106 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n5 0.612924
R4107 a_n9242_226.t0 a_n9242_226.n7 238.363
R4108 a_n9242_226.n7 a_n9242_226.t1 237.559
R4109 a_n9242_226.n2 a_n9242_226.n1 71.3963
R4110 a_n9242_226.n2 a_n9242_226.n0 71.3963
R4111 a_n9242_226.n5 a_n9242_226.n4 71.3963
R4112 a_n9242_226.n5 a_n9242_226.n3 71.3963
R4113 a_n9242_226.n1 a_n9242_226.t7 16.5305
R4114 a_n9242_226.n1 a_n9242_226.t4 16.5305
R4115 a_n9242_226.n0 a_n9242_226.t2 16.5305
R4116 a_n9242_226.n0 a_n9242_226.t9 16.5305
R4117 a_n9242_226.n4 a_n9242_226.t3 16.5305
R4118 a_n9242_226.n4 a_n9242_226.t8 16.5305
R4119 a_n9242_226.n3 a_n9242_226.t6 16.5305
R4120 a_n9242_226.n3 a_n9242_226.t5 16.5305
R4121 a_n9242_226.n7 a_n9242_226.n6 5.18724
R4122 a_n9242_226.n6 a_n9242_226.n2 0.3505
R4123 a_n9242_226.n6 a_n9242_226.n5 0.3505
R4124 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t10 134.734
R4125 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t13 134.734
R4126 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t9 134.734
R4127 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n6 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t8 134.734
R4128 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t11 134.734
R4129 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t15 134.734
R4130 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t14 134.734
R4131 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n7 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t12 134.734
R4132 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n11 79.7972
R4133 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n1 79.7972
R4134 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n0 79.7972
R4135 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n13 79.6389
R4136 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t4 9.23217
R4137 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n11 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t0 9.23217
R4138 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t5 9.23217
R4139 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t1 9.23217
R4140 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t2 9.23217
R4141 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t7 9.23217
R4142 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t3 9.23217
R4143 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n13 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t6 9.23217
R4144 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n3 9.2005
R4145 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n6 9.2005
R4146 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n5 6.63891
R4147 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n9 5.06405
R4148 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n5 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n4 4.5005
R4149 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n8 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n7 4.5005
R4150 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n9 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n8 4.43133
R4151 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n12 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n10 0.429667
R4152 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n10 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n2 0.429667
R4153 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n12 0.158833
R4154 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t1 231.236
R4155 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t0 231.129
R4156 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t2 230.782
R4157 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t3 230.272
R4158 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n0 1.03165
R4159 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n1 0.550258
R4160 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t3 146.001
R4161 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t2 144.221
R4162 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t0 143.886
R4163 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t1 143.494
R4164 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n1 0.424924
R4165 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n0 0.328076
R4166 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t1 231.016
R4167 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t0 230.996
R4168 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t2 230.959
R4169 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t3 230.272
R4170 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n0 0.968985
R4171 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n1 0.550258
C0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.22509f
C1 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.20881f
C2 P_IN[3] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.59591f
C3 a_n4955_n1462# opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.01975f
C4 a_n12122_4060# P_IN[4] 0.03952f
C5 opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_n1209_9323# 0.03145f
C6 P_IN[0] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.59672f
C7 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 P_IN[4] 0.06309f
C8 P_IN[2] P_IN[4] 0.43685f
C9 a_n1991_889# opa_folded_cascode_0.monticelli_top_0.A 0.02366f
C10 a_n5210_1510# a_n5758_1510# 0.0103f
C11 VDDA a_n1209_9323# 0.72706f
C12 a_n5758_3153# P_IN[0] 0.01212f
C13 a_n1613_4121# VDDA 0.54014f
C14 opa_folded_cascode_0.monticelli_top_0.Bx opa_folded_cascode_0.monticelli_top_0.A 0.4915f
C15 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 8.75672f
C16 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_folded_cascode_0.monticelli_top_0.A 0.37749f
C17 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_n5210_3153# 0.04959f
C18 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 8.23983f
C19 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.52521f
C20 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA N_IN 1.84784f
C21 a_n1209_n641# opa_folded_cascode_0.monticelli_top_0.Bx 0.05988f
C22 VDDA opa_folded_cascode_0.monticelli_top_0.A 3.89016f
C23 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 1.32033f
C24 VDDA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 2.24614f
C25 P_IN[1] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.59629f
C26 opa_folded_cascode_0.monticelli_top_0.B opa_folded_cascode_0.monticelli_top_0.A 5.08653f
C27 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.03879f
C28 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.48023f
C29 a_n5210_4060# N_IN 0.04644f
C30 a_n4030_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.01033f
C31 a_n5210_2008# N_IN 0.02204f
C32 a_n1991_10706# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.13435f
C33 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_folded_cascode_0.VB2 0.09525f
C34 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.0971f
C35 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_folded_cascode_0.VB2 0.16031f
C36 a_n5210_4060# VDDA 0.49886f
C37 a_n1209_5246# opa_folded_cascode_0.monticelli_top_0.A 0.0747f
C38 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA P_IN[4] 0.32156f
C39 opa_folded_cascode_0.VB1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.57726f
C40 a_n10394_1510# P_IN[3] 0.01061f
C41 a_n12122_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04134f
C42 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.44293f
C43 a_n7486_1510# N_IN 0.03463f
C44 P_IN[2] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.59606f
C45 P_IN[3] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.01305f
C46 a_n4030_4060# P_IN[0] 0.03029f
C47 opa_folded_cascode_0.VB2 opa_folded_cascode_0.monticelli_top_0.Ax 0.27696f
C48 a_n1613_3356# VDDA 0.53441f
C49 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_folded_cascode_0.VB2 0.06042f
C50 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.25263f
C51 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_folded_cascode_0.VB2 2.89603f
C52 a_n12122_1510# N_IN 0.04641f
C53 a_n1991_9323# a_n1209_9323# 0.02127f
C54 a_n1209_6513# a_n1991_6513# 0.02127f
C55 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.16361f
C56 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.56882f
C57 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 0.2177f
C58 a_n1209_6513# opa_folded_cascode_0.monticelli_top_0.Ax 0.01034f
C59 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 10.1642f
C60 a_n9214_1510# N_IN 0.03463f
C61 a_n5210_3153# N_IN 0.06743f
C62 P_IN[1] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.01667f
C63 a_n1209_1507# opa_folded_cascode_0.VB2 0.02948f
C64 a_n4030_2008# N_IN 0.0131f
C65 a_n1991_9323# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.05719f
C66 opa_folded_cascode_0.monticelli_top_0.Bx opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.12775f
C67 a_n12122_1510# P_IN[4] 0.01061f
C68 a_n5210_3153# VDDA 0.49013f
C69 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 6.01491f
C70 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 2.89925f
C71 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB N_IN 2.58453f
C72 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.05622f
C73 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 3.4882f
C74 VDDA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 2.32844f
C75 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.15175f
C76 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.33091f
C77 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.18445f
C78 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_folded_cascode_0.VB2 0.24606f
C79 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.43454f
C80 a_n10394_4060# a_n10942_4060# 0.0237f
C81 P_IN[1] a_n6938_2008# 0.03209f
C82 a_n12122_2008# N_IN 0.02119f
C83 a_n1991_10706# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.01199f
C84 a_n5210_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C85 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.17402f
C86 P_IN[2] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.66459f
C87 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.21785f
C88 a_n5210_1510# P_IN[0] 0.01061f
C89 a_n1613_4121# a_n949_4121# 0.01589f
C90 a_n10394_2008# N_IN 0.02203f
C91 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 1.39622f
C92 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 3.34137f
C93 a_n8666_3153# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.04959f
C94 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB P_IN[4] 0.07987f
C95 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 VOUT 0.03563f
C96 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 4.1684f
C97 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 12.2409f
C98 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_n1991_11973# 0.07653f
C99 a_n12122_3153# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.04134f
C100 a_n949_4121# opa_folded_cascode_0.monticelli_top_0.A 0.03043f
C101 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_folded_cascode_0.VB1 0.03137f
C102 VDDA opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 8.60419f
C103 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 5.28584f
C104 a_n5758_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.01033f
C105 a_n8666_4060# N_IN 0.04641f
C106 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 2.46853f
C107 a_n12122_2008# P_IN[4] 0.03389f
C108 a_n1209_11973# opa_folded_cascode_0.monticelli_top_0.Ax 0.09901f
C109 a_n10942_2008# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.0208f
C110 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.13043f
C111 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.13628f
C112 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.1736f
C113 a_n4030_1510# N_IN 0.039f
C114 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.57519f
C115 a_n1209_889# opa_folded_cascode_0.VB2 0.02948f
C116 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 10.1432f
C117 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.34329f
C118 a_n8666_4060# VDDA 0.49783f
C119 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.13217f
C120 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_folded_cascode_0.VB1 1.90588f
C121 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.09057f
C122 a_n4955_n34# opa_folded_cascode_0.VB2 0.0541f
C123 a_n4291_n1462# a_n4291_n2609# 0.015f
C124 a_n1613_2355# opa_folded_cascode_0.monticelli_top_0.B 0.03772f
C125 a_n10942_4060# N_IN 0.01454f
C126 opa_folded_cascode_0.VB1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 1.40678f
C127 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.61039f
C128 a_n6938_1510# N_IN 0.04471f
C129 a_n10942_4060# VDDA 0.49751f
C130 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.14299f
C131 P_IN[1] a_n5758_2008# 0.02844f
C132 a_n1991_6513# opa_folded_cascode_0.monticelli_top_0.Ax 0.06384f
C133 a_n8666_2008# P_IN[2] 0.03212f
C134 a_n1991_9323# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.01554f
C135 P_IN[0] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.01688f
C136 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_folded_cascode_0.VB2 4.37057f
C137 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_n1991_n23# 0.04394f
C138 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 7.06738f
C139 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.36581f
C140 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.0591f
C141 a_n5758_3153# a_n5210_3153# 0.0237f
C142 opa_folded_cascode_0.VB1 a_n4955_n2609# 0.10623f
C143 a_n6938_2008# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.0208f
C144 a_n10942_4060# P_IN[4] 0.03029f
C145 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.17799f
C146 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 0.13514f
C147 a_n949_3356# opa_folded_cascode_0.monticelli_top_0.A 0.03043f
C148 opa_folded_cascode_0.VB1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.22726f
C149 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.1193f
C150 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_folded_cascode_0.VB1 0.16742f
C151 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 2.84584f
C152 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.09533f
C153 a_n8666_1510# N_IN 0.04471f
C154 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_folded_cascode_0.monticelli_top_0.Bx 0.31237f
C155 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 1.27443f
C156 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 N_IN 0.09581f
C157 a_n8666_3153# N_IN 0.06741f
C158 P_IN[1] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.59788f
C159 a_n7486_4060# P_IN[1] 0.01175f
C160 VDDA opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 3.79805f
C161 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.78185f
C162 VDDA opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.1547f
C163 a_n12122_3153# N_IN 0.06888f
C164 a_n8666_3153# VDDA 0.49013f
C165 opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_n1209_8056# 0.03145f
C166 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.23878f
C167 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.63053f
C168 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.12567f
C169 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_folded_cascode_0.monticelli_top_0.B 0.26297f
C170 a_n12122_3153# VDDA 0.48f
C171 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 P_IN[3] 0.20612f
C172 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 1.57333f
C173 VDDA a_n1209_8056# 0.722f
C174 a_n8666_2008# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.0208f
C175 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.35096f
C176 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.11834f
C177 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.19454f
C178 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 1.09015f
C179 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 P_IN[0] 0.20524f
C180 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.14638f
C181 a_n7486_2008# P_IN[2] 0.02847f
C182 a_n8666_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C183 opa_folded_cascode_0.VB1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 3.43068f
C184 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.20768f
C185 P_IN[2] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.01317f
C186 a_n7486_4060# P_IN[2] 0.03029f
C187 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 1.88113f
C188 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_n1991_n641# 0.04179f
C189 a_n10942_3153# P_IN[3] 0.01201f
C190 a_n12122_3153# P_IN[4] 0.01862f
C191 a_n1613_3356# a_n949_3356# 0.01589f
C192 opa_folded_cascode_0.VB2 opa_folded_cascode_0.monticelli_top_0.A 0.35421f
C193 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_folded_cascode_0.monticelli_top_0.Bx 1.25574f
C194 a_n10394_1510# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.0208f
C195 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB N_IN 3.83784f
C196 N_IN opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.75441f
C197 opa_folded_cascode_0.monticelli_top_0.Bx VOUT 0.12771f
C198 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.20339f
C199 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.26862f
C200 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.20864f
C201 VDDA a_n4955_n2609# 0.72861f
C202 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 4.14638f
C203 a_n5758_2008# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.0208f
C204 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.63136f
C205 a_n10942_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C206 P_IN[3] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.01656f
C207 a_n1991_5246# opa_folded_cascode_0.monticelli_top_0.Ax 0.07145f
C208 a_n10394_3153# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.04959f
C209 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDA 1.85473f
C210 a_n4291_n34# opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.01297f
C211 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 P_IN[1] 0.20513f
C212 VDDA VOUT 1.08595f
C213 a_n10942_2008# a_n10394_2008# 0.0103f
C214 a_n1209_6513# opa_folded_cascode_0.monticelli_top_0.A 0.06525f
C215 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_folded_cascode_0.monticelli_top_0.B 0.01931f
C216 a_n6938_4060# N_IN 0.04641f
C217 opa_folded_cascode_0.monticelli_top_0.B VOUT 0.49893f
C218 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.98465f
C219 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.73274f
C220 a_n1209_889# opa_folded_cascode_0.monticelli_top_0.Ax 0.02366f
C221 a_n7486_3153# P_IN[1] 0.01208f
C222 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.61305f
C223 a_n5210_2008# a_n5758_2008# 0.0103f
C224 a_n6938_4060# VDDA 0.49751f
C225 a_n10394_4060# N_IN 0.04641f
C226 opa_folded_cascode_0.VB1 opa_folded_cascode_0.monticelli_top_0.Bx 1.1422f
C227 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 1.34502f
C228 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_folded_cascode_0.VB1 0.02575f
C229 opa_folded_cascode_0.VB1 N_IN 0.03415f
C230 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB P_IN[4] 0.05823f
C231 a_n10394_4060# VDDA 0.49886f
C232 VDDA opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 4.55333f
C233 VDDA opa_folded_cascode_0.VB1 7.28409f
C234 a_n7486_2008# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.0208f
C235 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.87726f
C236 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.11794f
C237 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 23.5069f
C238 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 P_IN[2] 0.20891f
C239 a_n4955_n1462# a_n4955_n2609# 0.015f
C240 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.28513f
C241 opa_folded_cascode_0.VB1 opa_folded_cascode_0.monticelli_top_0.B 0.38202f
C242 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.08235f
C243 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.21897f
C244 a_n10942_1510# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.02171f
C245 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 2.6115f
C246 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 1.24832f
C247 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.62163f
C248 a_n1991_8056# opa_folded_cascode_0.monticelli_top_0.A 0.06357f
C249 a_n9214_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.01035f
C250 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 8.67322f
C251 a_n5758_4060# P_IN[0] 0.01175f
C252 a_n1991_8056# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.0593f
C253 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.03344f
C254 P_IN[0] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.59734f
C255 opa_folded_cascode_0.monticelli_top_0.Bx a_n1991_n23# 0.02385f
C256 a_n9214_4060# P_IN[3] 0.03029f
C257 a_n8666_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.01034f
C258 a_n1209_10706# opa_folded_cascode_0.monticelli_top_0.Ax 0.0991f
C259 a_n7486_3153# a_n6938_3153# 0.0237f
C260 a_n1209_5246# opa_folded_cascode_0.VB1 0.0335f
C261 a_n1991_889# opa_folded_cascode_0.monticelli_top_0.Bx 0.0175f
C262 opa_folded_cascode_0.VB1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.23045f
C263 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.25378f
C264 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD a_n12122_4060# 0.01033f
C265 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 3.4669f
C266 P_IN[3] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.5977f
C267 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.18261f
C268 a_n5210_1510# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.0208f
C269 a_n4955_n1462# opa_folded_cascode_0.VB1 0.01613f
C270 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 3.39716f
C271 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 1.77943f
C272 opa_input_and_self_bias_0/cm_pcell3_0.VB2 N_IN 0.03859f
C273 P_IN[3] P_IN[0] 0.09964f
C274 P_IN[1] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.01299f
C275 a_n5758_4060# P_IN[1] 0.03029f
C276 VDDA opa_folded_cascode_0.monticelli_top_0.Bx 0.39566f
C277 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.15473f
C278 a_n1209_11973# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.06357f
C279 opa_input_and_self_bias_0/cm_pcell3_0.VB2 VDDA 25.2922f
C280 a_n10394_3153# N_IN 0.06741f
C281 VDDA N_IN 7.41634f
C282 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 11.2661f
C283 opa_folded_cascode_0.monticelli_top_0.B opa_folded_cascode_0.monticelli_top_0.Bx 2.34702f
C284 a_n10394_3153# VDDA 0.49013f
C285 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.84443f
C286 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT 24.2634f
C287 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.15608f
C288 a_n1209_9323# opa_folded_cascode_0.monticelli_top_0.Ax 0.06418f
C289 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_n5758_3153# 0.04994f
C290 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.3935f
C291 VDDA opa_folded_cascode_0.monticelli_top_0.B 2.19142f
C292 VDDA a_n1991_10706# 0.75792f
C293 VDDA opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.77292f
C294 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.32927f
C295 P_IN[4] N_IN 6.6392f
C296 a_n6938_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C297 P_IN[3] P_IN[1] 0.10582f
C298 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 1.05534f
C299 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.05844f
C300 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.14077f
C301 P_IN[1] P_IN[0] 4.11851f
C302 opa_folded_cascode_0.monticelli_top_0.A opa_folded_cascode_0.monticelli_top_0.Ax 4.43463f
C303 VDDA P_IN[4] 1.55121f
C304 a_n10394_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C305 VDDA a_n1209_5246# 0.72203f
C306 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.15777f
C307 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_folded_cascode_0.VB1 0.19101f
C308 opa_folded_cascode_0.monticelli_top_0.Ax opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 1.32808f
C309 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.70581f
C310 a_n9214_4060# P_IN[2] 0.01175f
C311 VDDA a_n1991_11973# 0.76867f
C312 a_n4291_464# a_n4291_n34# 0.015f
C313 a_n1209_5246# opa_folded_cascode_0.monticelli_top_0.B 0.08441f
C314 P_IN[0] opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.08765f
C315 opa_folded_cascode_0.monticelli_top_0.B a_n1991_n641# 0.02366f
C316 a_n949_4121# VOUT 0.01189f
C317 VDDA a_n4955_n1462# 0.79462f
C318 opa_input_and_self_bias_0/cm_pcell3_0.VB2 ROUT 0.02043f
C319 opa_folded_cascode_0.VB1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.0315f
C320 a_n1991_8056# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.01343f
C321 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.22101f
C322 P_IN[2] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.01655f
C323 P_IN[3] P_IN[2] 4.1241f
C324 VDDA ROUT 28.3503f
C325 a_n1209_1507# opa_folded_cascode_0.monticelli_top_0.A 0.06294f
C326 P_IN[2] P_IN[0] 0.09964f
C327 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_n1991_n23# 0.02444f
C328 a_n8666_2008# a_n9214_2008# 0.0103f
C329 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.13332f
C330 a_n5758_1510# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.02171f
C331 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 1.0059f
C332 opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_n1991_9323# 0.05095f
C333 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.16543f
C334 VDDA a_n1991_9323# 0.73351f
C335 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_folded_cascode_0.monticelli_top_0.Bx 1.70038f
C336 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA N_IN 1.91702f
C337 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 0.07698f
C338 P_IN[2] P_IN[1] 4.12484f
C339 VDDA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 1.90636f
C340 a_n5758_4060# a_n5210_4060# 0.0237f
C341 a_n5758_3153# N_IN 0.0409f
C342 a_n5210_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.01037f
C343 a_n1613_2711# a_n1613_2355# 0.02286f
C344 a_n9214_3153# P_IN[2] 0.01204f
C345 a_n6938_3153# P_IN[1] 0.01871f
C346 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.17446f
C347 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_folded_cascode_0.monticelli_top_0.B 0.33001f
C348 a_n5758_3153# VDDA 0.49013f
C349 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 2.81584f
C350 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 8.15945f
C351 P_IN[3] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.40148f
C352 a_n949_3356# VOUT 0.02398f
C353 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 3.9742f
C354 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_folded_cascode_0.VB2 0.19471f
C355 P_IN[0] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.40291f
C356 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA P_IN[4] 0.47247f
C357 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 0.79254f
C358 opa_folded_cascode_0.monticelli_top_0.Ax opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 1.33763f
C359 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_n1991_n641# 0.02628f
C360 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.39965f
C361 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.17464f
C362 a_n5210_4060# P_IN[0] 0.03805f
C363 a_n949_4121# VDDA 0.554f
C364 a_n5210_2008# P_IN[0] 0.03196f
C365 a_n949_2711# VOUT 0.0153f
C366 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_n4030_3153# 0.05017f
C367 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.07563f
C368 P_IN[1] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.40061f
C369 a_n10394_1510# N_IN 0.04471f
C370 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.21911f
C371 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 7.26391f
C372 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.5492f
C373 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD N_IN 0.67332f
C374 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.14677f
C375 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_folded_cascode_0.VB2 0.13276f
C376 a_n4030_4060# N_IN 0.0236f
C377 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 3.95069f
C378 opa_folded_cascode_0.VB2 VOUT 0.03299f
C379 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 2.35144f
C380 a_n1991_1507# opa_folded_cascode_0.VB2 0.04249f
C381 VDDA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.63708f
C382 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.07481f
C383 a_n4030_4060# VDDA 0.49013f
C384 a_n10942_2008# P_IN[4] 0.0287f
C385 a_n1991_8056# a_n1209_8056# 0.02127f
C386 P_IN[2] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.40094f
C387 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.08136f
C388 a_n6938_2008# N_IN 0.02203f
C389 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 opa_folded_cascode_0.VB1 0.16205f
C390 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 3.4847f
C391 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.39803f
C392 opa_folded_cascode_0.VB2 opa_folded_cascode_0.VB1 0.45991f
C393 a_n5210_3153# P_IN[0] 0.01852f
C394 a_n10942_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.01033f
C395 a_n949_3356# VDDA 0.53376f
C396 a_n4030_2008# P_IN[0] 0.02832f
C397 P_IN[3] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.20714f
C398 a_n10942_1510# N_IN 0.03463f
C399 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 3.18174f
C400 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 2.17542f
C401 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 1.00479f
C402 a_n949_2355# VOUT 0.01045f
C403 P_IN[0] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.20643f
C404 opa_folded_cascode_0.monticelli_top_0.A a_n1209_9323# 0.07342f
C405 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.32704f
C406 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.18431f
C407 a_n1209_6513# opa_folded_cascode_0.VB1 0.03145f
C408 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.3441f
C409 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.42152f
C410 a_n1613_4121# opa_folded_cascode_0.monticelli_top_0.A 0.04824f
C411 a_n8666_2008# N_IN 0.02203f
C412 a_n6938_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.01033f
C413 a_n7486_4060# a_n6938_4060# 0.0237f
C414 a_n4030_3153# N_IN 0.05095f
C415 a_n1991_889# opa_folded_cascode_0.VB2 0.04314f
C416 a_n5210_1510# N_IN 0.04473f
C417 opa_folded_cascode_0.monticelli_top_0.A opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.91896f
C418 P_IN[3] a_n10394_2008# 0.03215f
C419 a_n8666_4060# a_n9214_4060# 0.0237f
C420 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.11461f
C421 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.30956f
C422 a_n4030_3153# VDDA 0.48125f
C423 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 12.9813f
C424 a_n4291_464# opa_folded_cascode_0.VB2 0.06246f
C425 P_IN[1] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.20652f
C426 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 3.60244f
C427 a_n949_2711# opa_folded_cascode_0.monticelli_top_0.B 0.02725f
C428 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 N_IN 0.02759f
C429 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.53743f
C430 opa_folded_cascode_0.VB2 opa_folded_cascode_0.monticelli_top_0.Bx 1.48647f
C431 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_folded_cascode_0.VB2 1.16389f
C432 opa_folded_cascode_0.VB2 N_IN 0.05796f
C433 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.09585f
C434 VDDA opa_folded_cascode_0.VB2 4.40756f
C435 a_n1209_8056# opa_folded_cascode_0.monticelli_top_0.Ax 0.13749f
C436 a_n5210_2008# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.0208f
C437 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.96291f
C438 a_n1209_10706# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.06357f
C439 a_n4030_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C440 a_n1209_6513# opa_folded_cascode_0.monticelli_top_0.Bx 0.06357f
C441 opa_folded_cascode_0.VB2 opa_folded_cascode_0.monticelli_top_0.B 0.6182f
C442 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 opa_folded_cascode_0.VB1 0.3192f
C443 a_n1613_4121# a_n1613_3356# 0.02286f
C444 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.16159f
C445 a_n7486_3153# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.04994f
C446 VDDA a_n1209_6513# 0.722f
C447 P_IN[2] opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.20676f
C448 a_n10942_4060# P_IN[3] 0.01175f
C449 opa_folded_cascode_0.VB1 a_n4291_n1462# 0.11619f
C450 a_n10942_3153# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.04994f
C451 a_n1613_3356# opa_folded_cascode_0.monticelli_top_0.A 0.04784f
C452 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.20703f
C453 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 1.18645f
C454 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.22837f
C455 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 1.51685f
C456 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.13554f
C457 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.2482f
C458 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 1.8091f
C459 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD N_IN 0.6262f
C460 a_n7486_4060# N_IN 0.01454f
C461 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.92259f
C462 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 1.00408f
C463 a_n1991_1507# opa_folded_cascode_0.monticelli_top_0.Ax 0.05618f
C464 P_IN[3] a_n9214_2008# 0.02851f
C465 VDDA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.74227f
C466 a_n7486_4060# VDDA 0.49886f
C467 opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_n1991_8056# 0.05231f
C468 a_n4955_n2609# a_n4291_n2609# 0.02543f
C469 a_n949_2355# opa_folded_cascode_0.monticelli_top_0.B 0.02725f
C470 VDDA a_n1991_8056# 0.72849f
C471 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.41078f
C472 a_n1991_6513# opa_folded_cascode_0.VB1 0.0506f
C473 a_n1613_2711# opa_folded_cascode_0.monticelli_top_0.B 0.03745f
C474 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.32371f
C475 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.37208f
C476 a_n5758_1510# N_IN 0.03463f
C477 opa_folded_cascode_0.VB1 opa_folded_cascode_0.monticelli_top_0.Ax 1.45275f
C478 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 1.63629f
C479 P_IN[1] a_n6938_1510# 0.01061f
C480 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.37639f
C481 a_n4030_2008# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.02092f
C482 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 N_IN 0.02946f
C483 a_n8666_4060# P_IN[2] 0.03805f
C484 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 13.38f
C485 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_n1209_n23# 0.02981f
C486 a_n949_4121# a_n949_3356# 0.02286f
C487 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 1.00436f
C488 VDDA a_n4291_n1462# 0.73032f
C489 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 N_IN 0.21011f
C490 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 3.26761f
C491 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.46882f
C492 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.46005f
C493 VDDA a_n1209_11973# 0.73797f
C494 a_n4955_n34# opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.01106f
C495 a_n12122_2008# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.01625f
C496 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDA 11.2802f
C497 VDDA opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.65106f
C498 a_n7486_3153# N_IN 0.0409f
C499 a_n10394_2008# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.0208f
C500 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.06117f
C501 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.48886f
C502 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 1.00479f
C503 a_n8666_3153# a_n9214_3153# 0.0237f
C504 a_n7486_3153# VDDA 0.49013f
C505 a_n10942_3153# N_IN 0.0409f
C506 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB P_IN[3] 0.20421f
C507 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 2.48633f
C508 a_n10394_1510# a_n10942_1510# 0.0103f
C509 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.03331f
C510 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 3.04089f
C511 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 3.40713f
C512 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.54635f
C513 a_n7486_1510# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.02171f
C514 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 1.7781f
C515 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB P_IN[0] 0.2057f
C516 opa_folded_cascode_0.monticelli_top_0.Bx opa_folded_cascode_0.monticelli_top_0.Ax 4.04973f
C517 a_n10942_3153# a_n10394_3153# 0.0237f
C518 a_n10942_3153# VDDA 0.49013f
C519 VDDA a_n1991_6513# 0.72716f
C520 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_folded_cascode_0.monticelli_top_0.Ax 0.48335f
C521 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 10.7556f
C522 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD N_IN 0.61926f
C523 a_n1209_11973# a_n1991_11973# 0.02127f
C524 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 10.3151f
C525 a_n4955_n1462# a_n4291_n1462# 0.02543f
C526 VDDA opa_folded_cascode_0.monticelli_top_0.Ax 4.71077f
C527 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDA 48.6569f
C528 a_n1991_6513# opa_folded_cascode_0.monticelli_top_0.B 0.06357f
C529 VDDA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 2.42443f
C530 a_n8666_1510# P_IN[2] 0.01061f
C531 a_n12122_1510# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.01625f
C532 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.96164f
C533 a_n7486_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C534 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 4.44061f
C535 a_n10394_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.01033f
C536 opa_folded_cascode_0.monticelli_top_0.B opa_folded_cascode_0.monticelli_top_0.Ax 0.42504f
C537 a_n8666_3153# P_IN[2] 0.01867f
C538 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 1.03205f
C539 a_n10394_4060# P_IN[3] 0.03805f
C540 a_n1991_10706# opa_folded_cascode_0.monticelli_top_0.Ax 0.03151f
C541 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.4603f
C542 a_n1991_5246# opa_folded_cascode_0.VB1 0.0585f
C543 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.09063f
C544 a_n9214_1510# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.02171f
C545 VDDA a_n4291_n2609# 0.79433f
C546 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB P_IN[1] 0.20491f
C547 a_n4955_464# a_n4955_n34# 0.015f
C548 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 P_IN[4] 0.06879f
C549 a_n9214_3153# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.04994f
C550 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD P_IN[4] 0.59893f
C551 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN a_n4955_n2609# 0.01976f
C552 opa_folded_cascode_0.monticelli_top_0.Ax a_n1991_11973# 0.03145f
C553 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.08428f
C554 opa_folded_cascode_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 1.19048f
C555 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 5.81219f
C556 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VOUT 0.03648f
C557 a_n5758_4060# N_IN 0.01454f
C558 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.72782f
C559 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD N_IN 0.61932f
C560 a_n1209_1507# opa_folded_cascode_0.monticelli_top_0.B 0.01649f
C561 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 0.58085f
C562 a_n9214_2008# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.0208f
C563 a_n6938_4060# P_IN[1] 0.03805f
C564 a_n4955_464# opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 0.01003f
C565 a_n5758_4060# VDDA 0.49751f
C566 VDDA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 1.17943f
C567 a_n9214_4060# N_IN 0.01454f
C568 VDDA opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 1.40144f
C569 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 ROUT 0.0341f
C570 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB P_IN[2] 0.20447f
C571 a_n9214_4060# VDDA 0.49792f
C572 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.08957f
C573 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_n6938_3153# 0.04959f
C574 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.44079f
C575 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.08315f
C576 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.16693f
C577 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.09267f
C578 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_folded_cascode_0.VB1 0.45968f
C579 a_n7486_1510# a_n6938_1510# 0.0103f
C580 a_n1209_n641# opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.02965f
C581 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 1.2633f
C582 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD N_IN 0.62599f
C583 a_n1991_5246# opa_folded_cascode_0.monticelli_top_0.Bx 0.08404f
C584 opa_input_and_self_bias_0/cm_pcell3_0.VB2 P_IN[3] 0.01093f
C585 P_IN[3] N_IN 6.36642f
C586 a_n1209_8056# opa_folded_cascode_0.monticelli_top_0.A 0.02486f
C587 VDDA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 1.06003f
C588 opa_input_and_self_bias_0/cm_pcell3_0.VB2 P_IN[0] 0.0151f
C589 P_IN[0] N_IN 8.2946f
C590 opa_folded_cascode_0.monticelli_top_0.Bx a_n1209_n23# 0.02584f
C591 P_IN[3] VDDA 1.61008f
C592 a_n10394_3153# P_IN[3] 0.01864f
C593 a_n7486_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.01033f
C594 a_n1991_9323# opa_folded_cascode_0.monticelli_top_0.Ax 0.06368f
C595 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.04827f
C596 VDDA a_n1991_5246# 0.72637f
C597 P_IN[0] VDDA 1.99812f
C598 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.1884f
C599 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.1264f
C600 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.95801f
C601 opa_folded_cascode_0.monticelli_top_0.B a_n1209_n23# 0.03761f
C602 a_n4030_1510# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.02171f
C603 a_n7486_2008# a_n6938_2008# 0.0103f
C604 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD P_IN[4] 0.013f
C605 P_IN[3] P_IN[4] 4.45559f
C606 a_n1991_5246# a_n1209_5246# 0.02127f
C607 a_n1209_889# opa_folded_cascode_0.monticelli_top_0.B 0.02524f
C608 P_IN[1] N_IN 6.36674f
C609 P_IN[0] P_IN[4] 0.11402f
C610 opa_folded_cascode_0.monticelli_top_0.A VOUT 0.83749f
C611 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.61822f
C612 a_n9214_3153# N_IN 0.0409f
C613 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT 19.3099f
C614 P_IN[1] VDDA 1.61519f
C615 a_n6938_1510# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.0208f
C616 a_n9214_3153# VDDA 0.49013f
C617 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 2.66628f
C618 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN N_IN 0.31808f
C619 VDDA opa_input_and_self_bias_0/cm_ncell3_0.DRAIN 3.43281f
C620 a_n9214_1510# a_n8666_1510# 0.0103f
C621 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.1725f
C622 VDDA a_n1209_10706# 0.73997f
C623 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.0839f
C624 opa_folded_cascode_0.VB1 opa_folded_cascode_0.monticelli_top_0.A 0.6924f
C625 a_n5758_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C626 a_n12122_4060# N_IN 0.04557f
C627 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.95959f
C628 opa_folded_cascode_0.VB1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.69504f
C629 P_IN[1] P_IN[4] 0.43745f
C630 a_n949_2711# a_n949_2355# 0.02286f
C631 opa_input_and_self_bias_0/cm_pcell3_0.VB2 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 10.5012f
C632 opa_input_and_self_bias_0/cm_pcell3_0.VB2 P_IN[2] 0.01031f
C633 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 N_IN 0.03004f
C634 P_IN[2] N_IN 6.36553f
C635 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.15407f
C636 VDDA a_n12122_4060# 0.48931f
C637 a_n9214_4060# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C638 a_n6938_3153# N_IN 0.06741f
C639 a_n1991_10706# a_n1209_10706# 0.02127f
C640 VDDA opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 7.84417f
C641 a_n8666_1510# opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.0208f
C642 P_IN[2] VDDA 1.61107f
C643 a_n6938_3153# VDDA 0.49013f
C644 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.29164f
C645 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 1.16507f
C646 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.96164f
C647 VOUT GNDA 24.9907f
C648 P_IN[0] GNDA 5.34839f
C649 P_IN[1] GNDA 5.62173f
C650 P_IN[2] GNDA 5.55556f
C651 P_IN[3] GNDA 5.86506f
C652 N_IN GNDA 18.28604f
C653 P_IN[4] GNDA 6.82027f
C654 ROUT GNDA 13.44037f
C655 VDDA GNDA 0.3965p
C656 a_n1209_n641# GNDA 0.31627f $ **FLOATING
C657 a_n1991_n641# GNDA 0.3141f $ **FLOATING
C658 a_n1209_n23# GNDA 0.31363f $ **FLOATING
C659 a_n1991_n23# GNDA 0.31147f $ **FLOATING
C660 a_n4291_n2609# GNDA 0.10989f $ **FLOATING
C661 a_n4955_n2609# GNDA 0.11496f $ **FLOATING
C662 a_n4291_n1462# GNDA 0.10301f $ **FLOATING
C663 a_n4955_n1462# GNDA 0.11145f $ **FLOATING
C664 a_n1209_889# GNDA 0.31296f $ **FLOATING
C665 a_n1991_889# GNDA 0.31079f $ **FLOATING
C666 a_n1209_1507# GNDA 0.31297f $ **FLOATING
C667 a_n1991_1507# GNDA 0.31285f $ **FLOATING
C668 a_n4291_n34# GNDA 0.36693f $ **FLOATING
C669 a_n4955_n34# GNDA 0.35967f $ **FLOATING
C670 a_n4291_464# GNDA 0.34413f $ **FLOATING
C671 a_n4955_464# GNDA 0.38872f $ **FLOATING
C672 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 GNDA 1.37474f
C673 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 GNDA 1.32581f
C674 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 GNDA 1.4175f
C675 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GNDA 2.6963f
C676 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GNDA 3.3029f
C677 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GNDA 42.67636f
C678 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GNDA 8.84755f
C679 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GNDA 5.16437f
C680 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 GNDA 32.24463f
C681 a_n949_2355# GNDA 0.27787f $ **FLOATING
C682 a_n1613_2355# GNDA 0.27287f $ **FLOATING
C683 a_n949_2711# GNDA 0.26729f $ **FLOATING
C684 a_n1613_2711# GNDA 0.26729f $ **FLOATING
C685 a_n4030_1510# GNDA 0.23225f $ **FLOATING
C686 a_n5210_1510# GNDA 0.22396f $ **FLOATING
C687 a_n4030_2008# GNDA 0.23057f $ **FLOATING
C688 a_n5210_2008# GNDA 0.22049f $ **FLOATING
C689 a_n5758_1510# GNDA 0.22721f $ **FLOATING
C690 a_n6938_1510# GNDA 0.22504f $ **FLOATING
C691 a_n5758_2008# GNDA 0.2208f $ **FLOATING
C692 a_n6938_2008# GNDA 0.2208f $ **FLOATING
C693 a_n7486_1510# GNDA 0.22611f $ **FLOATING
C694 a_n8666_1510# GNDA 0.22485f $ **FLOATING
C695 a_n7486_2008# GNDA 0.2208f $ **FLOATING
C696 a_n8666_2008# GNDA 0.2208f $ **FLOATING
C697 a_n9214_1510# GNDA 0.22553f $ **FLOATING
C698 a_n10394_1510# GNDA 0.22626f $ **FLOATING
C699 a_n9214_2008# GNDA 0.2208f $ **FLOATING
C700 a_n10394_2008# GNDA 0.2208f $ **FLOATING
C701 a_n10942_1510# GNDA 0.2248f $ **FLOATING
C702 a_n12122_1510# GNDA 0.23775f $ **FLOATING
C703 a_n10942_2008# GNDA 0.2208f $ **FLOATING
C704 a_n12122_2008# GNDA 0.23134f $ **FLOATING
C705 a_n949_3356# GNDA 0.06968f $ **FLOATING
C706 a_n1613_3356# GNDA 0.06968f $ **FLOATING
C707 a_n949_4121# GNDA 0.06696f $ **FLOATING
C708 a_n1613_4121# GNDA 0.06696f $ **FLOATING
C709 a_n4030_3153# GNDA 0.03708f $ **FLOATING
C710 a_n4030_4060# GNDA 0.03501f $ **FLOATING
C711 a_n12122_3153# GNDA 0.03708f $ **FLOATING
C712 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB GNDA 5.37232f
C713 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA GNDA 11.80651f
C714 a_n12122_4060# GNDA 0.03439f $ **FLOATING
C715 a_n1209_5246# GNDA 0.04167f $ **FLOATING
C716 a_n1991_5246# GNDA 0.0358f $ **FLOATING
C717 a_n1209_6513# GNDA 0.04167f $ **FLOATING
C718 opa_folded_cascode_0.monticelli_top_0.Bx GNDA 10.82375f
C719 opa_folded_cascode_0.monticelli_top_0.B GNDA 6.70008f
C720 opa_folded_cascode_0.VB1 GNDA 5.83273f
C721 a_n1991_6513# GNDA 0.03283f $ **FLOATING
C722 a_n1209_8056# GNDA 0.04167f $ **FLOATING
C723 a_n1991_8056# GNDA 0.03182f $ **FLOATING
C724 a_n1209_9323# GNDA 0.04167f $ **FLOATING
C725 opa_folded_cascode_0.monticelli_top_0.A GNDA 2.77007f
C726 a_n1991_9323# GNDA 0.03182f $ **FLOATING
C727 a_n1209_10706# GNDA 0.04167f $ **FLOATING
C728 a_n1991_10706# GNDA 0.03283f $ **FLOATING
C729 a_n1209_11973# GNDA 0.04712f $ **FLOATING
C730 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GNDA 9.34486f
C731 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GNDA 4.56814f
C732 opa_folded_cascode_0.monticelli_top_0.Ax GNDA 2.79544f
C733 a_n1991_11973# GNDA 0.03804f $ **FLOATING
C734 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD GNDA 0.75655f
C735 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD GNDA 0.97515f
C736 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD GNDA 0.89487f
C737 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD GNDA 1.35942f
C738 opa_folded_cascode_0.VB2 GNDA 5.26252f
C739 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD GNDA 1.8513f
C740 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN GNDA 44.43706f
C741 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 GNDA 0.72361f
C742 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 GNDA 0.5471f
C743 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 GNDA 0.53866f
C744 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 GNDA 1.39706f
C745 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 GNDA 1.1991f
C746 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 GNDA 2.15001f
C747 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 GNDA 1.69093f
C748 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 GNDA 1.65173f
C749 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 GNDA 16.20341f
C750 opa_input_and_self_bias_0/cm_pcell3_0.VB2 GNDA 17.05692f
C751 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t1 GNDA 0.05654f
C752 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t0 GNDA 0.05718f
C753 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n0 GNDA 1.04424f
C754 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t2 GNDA 0.05624f
C755 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.t3 GNDA 0.0538f
C756 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0.n1 GNDA 0.81076f
C757 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t1 GNDA 0.19229f
C758 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t0 GNDA 0.20585f
C759 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n0 GNDA 1.53847f
C760 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t3 GNDA 0.22982f
C761 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.t2 GNDA 0.21285f
C762 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0.n1 GNDA 2.80418f
C763 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t0 GNDA 0.05778f
C764 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t1 GNDA 0.05865f
C765 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n0 GNDA 1.04124f
C766 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t2 GNDA 0.05535f
C767 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.t3 GNDA 0.054f
C768 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1.n1 GNDA 0.78821f
C769 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t2 GNDA 0.04627f
C770 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t7 GNDA 0.04627f
C771 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n0 GNDA 0.10972f
C772 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t5 GNDA 0.04627f
C773 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t1 GNDA 0.04627f
C774 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n1 GNDA 0.10972f
C775 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n2 GNDA 0.63006f
C776 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t15 GNDA 0.10271f
C777 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t11 GNDA 0.10271f
C778 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n3 GNDA 0.61687f
C779 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t13 GNDA 0.10271f
C780 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t10 GNDA 0.10271f
C781 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n4 GNDA 0.42623f
C782 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n5 GNDA 0.92706f
C783 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t8 GNDA 0.10271f
C784 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t9 GNDA 0.10271f
C785 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n6 GNDA 0.61598f
C786 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t12 GNDA 0.10271f
C787 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t14 GNDA 0.10271f
C788 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n7 GNDA 0.42711f
C789 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n8 GNDA 0.68929f
C790 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n9 GNDA 1.50345f
C791 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n10 GNDA 0.20317f
C792 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t4 GNDA 0.04627f
C793 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t0 GNDA 0.04627f
C794 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n11 GNDA 0.10972f
C795 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n12 GNDA 0.34359f
C796 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t3 GNDA 0.04627f
C797 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.t6 GNDA 0.04627f
C798 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD.n13 GNDA 0.10915f
C799 a_n9242_226.t2 GNDA 0.02366f
C800 a_n9242_226.t9 GNDA 0.02366f
C801 a_n9242_226.n0 GNDA 0.05487f
C802 a_n9242_226.t7 GNDA 0.02366f
C803 a_n9242_226.t4 GNDA 0.02366f
C804 a_n9242_226.n1 GNDA 0.05487f
C805 a_n9242_226.n2 GNDA 0.40357f
C806 a_n9242_226.t6 GNDA 0.02366f
C807 a_n9242_226.t5 GNDA 0.02366f
C808 a_n9242_226.n3 GNDA 0.05487f
C809 a_n9242_226.t3 GNDA 0.02366f
C810 a_n9242_226.t8 GNDA 0.02366f
C811 a_n9242_226.n4 GNDA 0.05487f
C812 a_n9242_226.n5 GNDA 0.40357f
C813 a_n9242_226.n6 GNDA 0.32667f
C814 a_n9242_226.t1 GNDA 0.11399f
C815 a_n9242_226.n7 GNDA 5.31895f
C816 a_n9242_226.t0 GNDA 0.12455f
C817 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t0 GNDA 0.12074f
C818 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t1 GNDA 0.12074f
C819 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n0 GNDA 0.65062f
C820 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t3 GNDA 0.12074f
C821 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t2 GNDA 0.12074f
C822 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n1 GNDA 0.70506f
C823 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n2 GNDA 0.74687f
C824 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t4 GNDA 0.13368f
C825 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t7 GNDA 0.13005f
C826 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n3 GNDA 1.04458f
C827 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t5 GNDA 0.13368f
C828 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.t6 GNDA 0.13005f
C829 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n4 GNDA 0.85678f
C830 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2.n5 GNDA 0.82256f
C831 a_n11843_11539.t5 GNDA 0.08912f
C832 a_n11843_11539.t4 GNDA 0.23322f
C833 a_n11843_11539.n0 GNDA 2.67545f
C834 a_n11843_11539.t0 GNDA 8.34107f
C835 a_n11843_11539.t7 GNDA 6.50682f
C836 a_n11843_11539.n1 GNDA 3.76814f
C837 a_n11843_11539.n2 GNDA 0.53672f
C838 a_n11843_11539.t6 GNDA 8.34107f
C839 a_n11843_11539.t2 GNDA 6.50682f
C840 a_n11843_11539.n3 GNDA 3.96571f
C841 a_n11843_11539.n4 GNDA 0.57813f
C842 a_n11843_11539.t1 GNDA 0.30099f
C843 a_n11843_11539.n5 GNDA 2.46761f
C844 a_n11843_11539.t3 GNDA 0.08912f
C845 ROUT.t4 GNDA 7.10369f
C846 ROUT.t2 GNDA 5.54155f
C847 ROUT.n0 GNDA 3.3774f
C848 ROUT.t3 GNDA 0.0759f
C849 ROUT.t1 GNDA 0.25634f
C850 ROUT.n1 GNDA 2.1133f
C851 ROUT.t0 GNDA 7.10369f
C852 ROUT.t5 GNDA 5.54155f
C853 ROUT.n2 GNDA 3.20579f
C854 ROUT.n3 GNDA 0.38258f
C855 ROUT.n4 GNDA 0.48914f
C856 P_IN[3].t7 GNDA 0.92458f
C857 P_IN[3].t3 GNDA 0.91882f
C858 P_IN[3].n0 GNDA 1.42783f
C859 P_IN[3].t5 GNDA 0.37774f
C860 P_IN[3].t0 GNDA 0.37592f
C861 P_IN[3].n1 GNDA 0.99837f
C862 P_IN[3].t6 GNDA 0.38397f
C863 P_IN[3].t2 GNDA 0.37748f
C864 P_IN[3].n2 GNDA 1.11206f
C865 P_IN[3].n3 GNDA 0.51849f
C866 P_IN[3].n4 GNDA 1.54154f
C867 P_IN[3].t1 GNDA 0.91943f
C868 P_IN[3].t4 GNDA 0.91775f
C869 P_IN[3].n5 GNDA 1.1838f
C870 P_IN[3].n6 GNDA 0.35605f
C871 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t0 GNDA 0.199f
C872 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t1 GNDA 0.21007f
C873 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n0 GNDA 1.52173f
C874 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t2 GNDA 0.24388f
C875 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.t3 GNDA 0.22393f
C876 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1.n1 GNDA 3.07321f
C877 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t4 GNDA 0.02214f
C878 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t0 GNDA 0.02214f
C879 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n0 GNDA 0.0525f
C880 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t1 GNDA 0.02214f
C881 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t5 GNDA 0.02214f
C882 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n1 GNDA 0.0525f
C883 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n2 GNDA 0.3015f
C884 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t9 GNDA 0.07201f
C885 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t8 GNDA 0.06819f
C886 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n3 GNDA 1.29541f
C887 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n4 GNDA 0.07426f
C888 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t2 GNDA 0.02214f
C889 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t6 GNDA 0.02214f
C890 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n5 GNDA 0.0525f
C891 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n6 GNDA 0.16442f
C892 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t7 GNDA 0.02214f
C893 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.t3 GNDA 0.02214f
C894 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD.n7 GNDA 0.05223f
C895 opa_folded_cascode_0.VB1.t8 GNDA 0.57153f
C896 opa_folded_cascode_0.VB1.t10 GNDA 0.57173f
C897 opa_folded_cascode_0.VB1.t15 GNDA 0.57394f
C898 opa_folded_cascode_0.VB1.t13 GNDA 0.57311f
C899 opa_folded_cascode_0.VB1.n0 GNDA 0.57028f
C900 opa_folded_cascode_0.VB1.t12 GNDA 0.57394f
C901 opa_folded_cascode_0.VB1.t14 GNDA 0.57311f
C902 opa_folded_cascode_0.VB1.n1 GNDA 0.5671f
C903 opa_folded_cascode_0.VB1.n2 GNDA 1.86177f
C904 opa_folded_cascode_0.VB1.n3 GNDA 2.60622f
C905 opa_folded_cascode_0.VB1.t11 GNDA 0.17341f
C906 opa_folded_cascode_0.VB1.n4 GNDA 0.23921f
C907 opa_folded_cascode_0.VB1.t5 GNDA 0.02203f
C908 opa_folded_cascode_0.VB1.t1 GNDA 0.02203f
C909 opa_folded_cascode_0.VB1.n5 GNDA 0.45415f
C910 opa_folded_cascode_0.VB1.n6 GNDA 0.47964f
C911 opa_folded_cascode_0.VB1.t7 GNDA 0.02201f
C912 opa_folded_cascode_0.VB1.n7 GNDA 0.07372f
C913 opa_folded_cascode_0.VB1.t3 GNDA 0.02201f
C914 opa_folded_cascode_0.VB1.n8 GNDA 0.07372f
C915 opa_folded_cascode_0.VB1.n9 GNDA 0.32363f
C916 opa_folded_cascode_0.VB1.t2 GNDA 0.02203f
C917 opa_folded_cascode_0.VB1.t6 GNDA 0.02203f
C918 opa_folded_cascode_0.VB1.n10 GNDA 0.45415f
C919 opa_folded_cascode_0.VB1.n11 GNDA 0.47964f
C920 opa_folded_cascode_0.VB1.t4 GNDA 0.02201f
C921 opa_folded_cascode_0.VB1.n12 GNDA 0.07372f
C922 opa_folded_cascode_0.VB1.t0 GNDA 0.02201f
C923 opa_folded_cascode_0.VB1.n13 GNDA 0.07372f
C924 opa_folded_cascode_0.VB1.n14 GNDA 0.19305f
C925 opa_folded_cascode_0.VB1.n15 GNDA 0.64379f
C926 opa_folded_cascode_0.VB1.n16 GNDA 0.22337f
C927 opa_folded_cascode_0.VB1.t9 GNDA 0.17341f
C928 opa_folded_cascode_0.VB1.n17 GNDA 0.20786f
C929 opa_folded_cascode_0.VB1.n18 GNDA 0.22442f
C930 a_n10488_226.t4 GNDA 0.02333f
C931 a_n10488_226.t1 GNDA 0.02333f
C932 a_n10488_226.n0 GNDA 0.21448f
C933 a_n10488_226.t8 GNDA 0.01041f
C934 a_n10488_226.t12 GNDA 0.01041f
C935 a_n10488_226.n1 GNDA 0.02413f
C936 a_n10488_226.t14 GNDA 0.01041f
C937 a_n10488_226.t10 GNDA 0.01041f
C938 a_n10488_226.n2 GNDA 0.02413f
C939 a_n10488_226.n3 GNDA 0.17752f
C940 a_n10488_226.t11 GNDA 0.01041f
C941 a_n10488_226.t9 GNDA 0.01041f
C942 a_n10488_226.n4 GNDA 0.02413f
C943 a_n10488_226.t15 GNDA 0.01041f
C944 a_n10488_226.t13 GNDA 0.01041f
C945 a_n10488_226.n5 GNDA 0.02413f
C946 a_n10488_226.n6 GNDA 0.17752f
C947 a_n10488_226.n7 GNDA 0.07503f
C948 a_n10488_226.t0 GNDA 0.02333f
C949 a_n10488_226.t5 GNDA 0.02333f
C950 a_n10488_226.n8 GNDA 0.35392f
C951 a_n10488_226.n9 GNDA 0.34189f
C952 a_n10488_226.t2 GNDA 0.0233f
C953 a_n10488_226.n10 GNDA 0.09101f
C954 a_n10488_226.t6 GNDA 0.0233f
C955 a_n10488_226.n11 GNDA 0.09101f
C956 a_n10488_226.n12 GNDA 0.08577f
C957 a_n10488_226.n13 GNDA 0.63923f
C958 a_n10488_226.n14 GNDA 0.38663f
C959 a_n10488_226.t3 GNDA 0.02333f
C960 a_n10488_226.n15 GNDA 0.29964f
C961 a_n10488_226.t7 GNDA 0.02333f
C962 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t3 GNDA 0.03385f
C963 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t2 GNDA 0.03293f
C964 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n0 GNDA 0.67533f
C965 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t0 GNDA 0.03385f
C966 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t1 GNDA 0.03293f
C967 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n1 GNDA 0.52074f
C968 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n2 GNDA 0.64975f
C969 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t4 GNDA 0.02952f
C970 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t6 GNDA 0.02948f
C971 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n3 GNDA 0.2736f
C972 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t5 GNDA 0.02952f
C973 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.t7 GNDA 0.02948f
C974 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n4 GNDA 0.29926f
C975 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2.n5 GNDA 0.58174f
C976 opa_folded_cascode_0.monticelli_top_0.Ax.t1 GNDA 0.28451f
C977 opa_folded_cascode_0.monticelli_top_0.Ax.t8 GNDA 0.87667f
C978 opa_folded_cascode_0.monticelli_top_0.Ax.t6 GNDA 0.86819f
C979 opa_folded_cascode_0.monticelli_top_0.Ax.n0 GNDA 1.06648f
C980 opa_folded_cascode_0.monticelli_top_0.Ax.t7 GNDA 0.86819f
C981 opa_folded_cascode_0.monticelli_top_0.Ax.t9 GNDA 0.87667f
C982 opa_folded_cascode_0.monticelli_top_0.Ax.n1 GNDA 0.71078f
C983 opa_folded_cascode_0.monticelli_top_0.Ax.n2 GNDA 0.54423f
C984 opa_folded_cascode_0.monticelli_top_0.Ax.t3 GNDA 0.27375f
C985 opa_folded_cascode_0.monticelli_top_0.Ax.t2 GNDA 0.28821f
C986 opa_folded_cascode_0.monticelli_top_0.Ax.n3 GNDA 1.07924f
C987 opa_folded_cascode_0.monticelli_top_0.Ax.n4 GNDA 0.81885f
C988 opa_folded_cascode_0.monticelli_top_0.Ax.t0 GNDA 0.36911f
C989 opa_folded_cascode_0.monticelli_top_0.Ax.n5 GNDA 1.30848f
C990 opa_folded_cascode_0.monticelli_top_0.Ax.n6 GNDA 1.17185f
C991 opa_folded_cascode_0.monticelli_top_0.Ax.t4 GNDA 0.08638f
C992 opa_folded_cascode_0.monticelli_top_0.Ax.t5 GNDA 0.09208f
C993 opa_folded_cascode_0.monticelli_top_0.Ax.n7 GNDA 0.92476f
C994 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t0 GNDA 0.18452f
C995 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t5 GNDA 0.18452f
C996 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n0 GNDA 1.4305f
C997 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t1 GNDA 0.18452f
C998 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t2 GNDA 0.18452f
C999 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n1 GNDA 1.05912f
C1000 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n2 GNDA 2.27113f
C1001 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t6 GNDA 0.18452f
C1002 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t7 GNDA 0.18452f
C1003 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n3 GNDA 1.25158f
C1004 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t3 GNDA 0.18452f
C1005 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t4 GNDA 0.18452f
C1006 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n4 GNDA 1.22182f
C1007 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n5 GNDA 2.22498f
C1008 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n6 GNDA 0.81562f
C1009 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t12 GNDA 0.20184f
C1010 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t9 GNDA 0.19632f
C1011 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n7 GNDA 1.73221f
C1012 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t11 GNDA 0.20184f
C1013 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t10 GNDA 0.19673f
C1014 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n8 GNDA 1.70817f
C1015 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n9 GNDA 1.43567f
C1016 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t13 GNDA 0.20184f
C1017 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t8 GNDA 0.19673f
C1018 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n10 GNDA 1.96104f
C1019 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t15 GNDA 0.20184f
C1020 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.t14 GNDA 0.19632f
C1021 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n11 GNDA 1.47934f
C1022 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n12 GNDA 1.32744f
C1023 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2.n13 GNDA 1.11227f
C1024 P_IN[0].t0 GNDA 0.76432f
C1025 P_IN[0].t4 GNDA 0.75955f
C1026 P_IN[0].n0 GNDA 1.18034f
C1027 P_IN[0].t1 GNDA 0.31227f
C1028 P_IN[0].t6 GNDA 0.31076f
C1029 P_IN[0].n1 GNDA 0.82532f
C1030 P_IN[0].t7 GNDA 0.31742f
C1031 P_IN[0].t3 GNDA 0.31205f
C1032 P_IN[0].n2 GNDA 0.9193f
C1033 P_IN[0].n3 GNDA 0.48205f
C1034 P_IN[0].n4 GNDA 1.2493f
C1035 P_IN[0].t5 GNDA 0.76006f
C1036 P_IN[0].t2 GNDA 0.75867f
C1037 P_IN[0].n5 GNDA 0.97861f
C1038 P_IN[0].n6 GNDA 0.24091f
C1039 a_n9242_n890.t2 GNDA 0.01193f
C1040 a_n9242_n890.t7 GNDA 0.01193f
C1041 a_n9242_n890.n0 GNDA 0.02768f
C1042 a_n9242_n890.t8 GNDA 0.01193f
C1043 a_n9242_n890.t5 GNDA 0.01193f
C1044 a_n9242_n890.n1 GNDA 0.02768f
C1045 a_n9242_n890.n2 GNDA 0.2036f
C1046 a_n9242_n890.t6 GNDA 0.01193f
C1047 a_n9242_n890.t3 GNDA 0.01193f
C1048 a_n9242_n890.n3 GNDA 0.02768f
C1049 a_n9242_n890.t4 GNDA 0.01193f
C1050 a_n9242_n890.t9 GNDA 0.01193f
C1051 a_n9242_n890.n4 GNDA 0.02768f
C1052 a_n9242_n890.n5 GNDA 0.2036f
C1053 a_n9242_n890.n6 GNDA 0.11865f
C1054 a_n9242_n890.t1 GNDA 0.05399f
C1055 a_n9242_n890.n7 GNDA 2.06772f
C1056 a_n9242_n890.t0 GNDA 0.04624f
C1057 P_IN[1].t5 GNDA 0.89992f
C1058 P_IN[1].t4 GNDA 0.89431f
C1059 P_IN[1].n0 GNDA 1.38976f
C1060 P_IN[1].t2 GNDA 0.36767f
C1061 P_IN[1].t1 GNDA 0.3659f
C1062 P_IN[1].n1 GNDA 0.97175f
C1063 P_IN[1].t3 GNDA 0.37373f
C1064 P_IN[1].t0 GNDA 0.36742f
C1065 P_IN[1].n2 GNDA 1.0824f
C1066 P_IN[1].n3 GNDA 0.5466f
C1067 P_IN[1].n4 GNDA 1.66914f
C1068 P_IN[1].t7 GNDA 0.89491f
C1069 P_IN[1].t6 GNDA 0.89327f
C1070 P_IN[1].n5 GNDA 1.15223f
C1071 P_IN[1].n6 GNDA 0.30462f
C1072 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t0 GNDA 0.09331f
C1073 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t6 GNDA 0.09112f
C1074 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n0 GNDA 1.29109f
C1075 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t4 GNDA 0.09331f
C1076 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t3 GNDA 0.09112f
C1077 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n1 GNDA 1.44549f
C1078 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n2 GNDA 1.38567f
C1079 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t2 GNDA 0.09331f
C1080 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t1 GNDA 0.09112f
C1081 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n3 GNDA 1.60154f
C1082 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t7 GNDA 0.09331f
C1083 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t5 GNDA 0.09112f
C1084 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n4 GNDA 1.13504f
C1085 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n5 GNDA 1.29052f
C1086 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n6 GNDA 1.36983f
C1087 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t8 GNDA 0.08941f
C1088 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t13 GNDA 0.08941f
C1089 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n7 GNDA 0.95504f
C1090 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t14 GNDA 0.08941f
C1091 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t11 GNDA 0.08941f
C1092 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n8 GNDA 0.62001f
C1093 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n9 GNDA 2.44269f
C1094 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t12 GNDA 0.08941f
C1095 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t9 GNDA 0.08941f
C1096 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n10 GNDA 0.7235f
C1097 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t10 GNDA 0.08941f
C1098 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.t15 GNDA 0.08941f
C1099 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n11 GNDA 0.83514f
C1100 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n12 GNDA 2.41198f
C1101 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1.n13 GNDA 0.91107f
C1102 opa_folded_cascode_0.monticelli_top_0.Bx.t2 GNDA 0.18007f
C1103 opa_folded_cascode_0.monticelli_top_0.Bx.t3 GNDA 0.13294f
C1104 opa_folded_cascode_0.monticelli_top_0.Bx.n0 GNDA 0.61683f
C1105 opa_folded_cascode_0.monticelli_top_0.Bx.t5 GNDA 0.04257f
C1106 opa_folded_cascode_0.monticelli_top_0.Bx.t12 GNDA 0.16546f
C1107 opa_folded_cascode_0.monticelli_top_0.Bx.t11 GNDA 0.1651f
C1108 opa_folded_cascode_0.monticelli_top_0.Bx.n1 GNDA 0.19224f
C1109 opa_folded_cascode_0.monticelli_top_0.Bx.t14 GNDA 0.1651f
C1110 opa_folded_cascode_0.monticelli_top_0.Bx.n2 GNDA 0.09113f
C1111 opa_folded_cascode_0.monticelli_top_0.Bx.t10 GNDA 0.16546f
C1112 opa_folded_cascode_0.monticelli_top_0.Bx.t6 GNDA 0.1651f
C1113 opa_folded_cascode_0.monticelli_top_0.Bx.n3 GNDA 0.19224f
C1114 opa_folded_cascode_0.monticelli_top_0.Bx.t16 GNDA 0.1651f
C1115 opa_folded_cascode_0.monticelli_top_0.Bx.n4 GNDA 0.09113f
C1116 opa_folded_cascode_0.monticelli_top_0.Bx.n5 GNDA 0.08771f
C1117 opa_folded_cascode_0.monticelli_top_0.Bx.t9 GNDA 0.16546f
C1118 opa_folded_cascode_0.monticelli_top_0.Bx.t8 GNDA 0.1651f
C1119 opa_folded_cascode_0.monticelli_top_0.Bx.n6 GNDA 0.19224f
C1120 opa_folded_cascode_0.monticelli_top_0.Bx.t13 GNDA 0.1651f
C1121 opa_folded_cascode_0.monticelli_top_0.Bx.n7 GNDA 0.09113f
C1122 opa_folded_cascode_0.monticelli_top_0.Bx.t7 GNDA 0.16546f
C1123 opa_folded_cascode_0.monticelli_top_0.Bx.t17 GNDA 0.1651f
C1124 opa_folded_cascode_0.monticelli_top_0.Bx.n8 GNDA 0.19224f
C1125 opa_folded_cascode_0.monticelli_top_0.Bx.t15 GNDA 0.1651f
C1126 opa_folded_cascode_0.monticelli_top_0.Bx.n9 GNDA 0.09113f
C1127 opa_folded_cascode_0.monticelli_top_0.Bx.n10 GNDA 0.21002f
C1128 opa_folded_cascode_0.monticelli_top_0.Bx.t0 GNDA 0.04195f
C1129 opa_folded_cascode_0.monticelli_top_0.Bx.t1 GNDA 0.04451f
C1130 opa_folded_cascode_0.monticelli_top_0.Bx.n11 GNDA 0.29215f
C1131 opa_folded_cascode_0.monticelli_top_0.Bx.n12 GNDA 0.21628f
C1132 opa_folded_cascode_0.monticelli_top_0.Bx.n13 GNDA 0.28139f
C1133 opa_folded_cascode_0.monticelli_top_0.Bx.t4 GNDA 0.06193f
C1134 opa_folded_cascode_0.monticelli_top_0.Bx.n14 GNDA 0.50309f
C1135 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t5 GNDA 0.09798f
C1136 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t2 GNDA 0.09517f
C1137 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n0 GNDA 0.98853f
C1138 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t0 GNDA 0.09798f
C1139 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t7 GNDA 0.09517f
C1140 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n1 GNDA 1.57121f
C1141 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n2 GNDA 0.81058f
C1142 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t3 GNDA 0.09798f
C1143 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t1 GNDA 0.09517f
C1144 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n3 GNDA 1.30559f
C1145 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t4 GNDA 0.09798f
C1146 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t6 GNDA 0.09517f
C1147 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n4 GNDA 1.25415f
C1148 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n5 GNDA 0.68388f
C1149 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n6 GNDA 1.49193f
C1150 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t11 GNDA 0.09131f
C1151 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t9 GNDA 0.09131f
C1152 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n7 GNDA 0.63869f
C1153 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t13 GNDA 0.09131f
C1154 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t10 GNDA 0.09131f
C1155 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n8 GNDA 0.60876f
C1156 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n9 GNDA 1.68727f
C1157 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t8 GNDA 0.09131f
C1158 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t14 GNDA 0.09131f
C1159 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n10 GNDA 0.48631f
C1160 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t15 GNDA 0.09131f
C1161 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.t12 GNDA 0.09131f
C1162 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n11 GNDA 0.81419f
C1163 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n12 GNDA 1.56335f
C1164 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3.n13 GNDA 1.03015f
C1165 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t5 GNDA 0.07931f
C1166 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t1 GNDA 0.07931f
C1167 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n0 GNDA 0.18806f
C1168 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t2 GNDA 0.07931f
C1169 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t4 GNDA 0.07931f
C1170 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n1 GNDA 0.18806f
C1171 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n2 GNDA 1.07994f
C1172 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t20 GNDA 0.19984f
C1173 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t17 GNDA 0.176f
C1174 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t21 GNDA 0.176f
C1175 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n3 GNDA 0.72684f
C1176 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n4 GNDA 2.09379f
C1177 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t22 GNDA 0.176f
C1178 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t13 GNDA 0.176f
C1179 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n5 GNDA 0.72829f
C1180 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n6 GNDA 1.44342f
C1181 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t14 GNDA 0.176f
C1182 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t15 GNDA 0.176f
C1183 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n7 GNDA 0.72829f
C1184 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n8 GNDA 0.60469f
C1185 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t19 GNDA 0.18546f
C1186 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n9 GNDA 0.5189f
C1187 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t8 GNDA 0.19033f
C1188 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t10 GNDA 0.176f
C1189 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t16 GNDA 0.176f
C1190 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n10 GNDA 0.72829f
C1191 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n11 GNDA 1.0751f
C1192 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t9 GNDA 0.176f
C1193 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t18 GNDA 0.176f
C1194 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n12 GNDA 0.72829f
C1195 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n13 GNDA 1.44342f
C1196 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t11 GNDA 0.176f
C1197 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t12 GNDA 0.176f
C1198 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n14 GNDA 0.72684f
C1199 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n15 GNDA 1.42725f
C1200 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t23 GNDA 0.18546f
C1201 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n16 GNDA 0.69316f
C1202 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n17 GNDA 1.65076f
C1203 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n18 GNDA 0.36304f
C1204 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t0 GNDA 0.07931f
C1205 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t6 GNDA 0.07931f
C1206 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n19 GNDA 0.18806f
C1207 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n20 GNDA 0.58892f
C1208 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t7 GNDA 0.07931f
C1209 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.t3 GNDA 0.07931f
C1210 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD.n21 GNDA 0.18708f
C1211 P_IN[4].t4 GNDA 0.68419f
C1212 P_IN[4].t0 GNDA 0.67992f
C1213 P_IN[4].n0 GNDA 1.0566f
C1214 P_IN[4].t7 GNDA 0.27953f
C1215 P_IN[4].t6 GNDA 0.27818f
C1216 P_IN[4].n1 GNDA 0.73879f
C1217 P_IN[4].t3 GNDA 0.28414f
C1218 P_IN[4].t5 GNDA 0.27934f
C1219 P_IN[4].n2 GNDA 0.82292f
C1220 P_IN[4].n3 GNDA 0.36774f
C1221 P_IN[4].n4 GNDA 0.18382f
C1222 P_IN[4].t2 GNDA 0.68038f
C1223 P_IN[4].t1 GNDA 0.67913f
C1224 P_IN[4].n5 GNDA 0.87601f
C1225 P_IN[4].n6 GNDA 0.27942f
C1226 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t1 GNDA 0.10578f
C1227 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t10 GNDA 0.17177f
C1228 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t11 GNDA 0.04571f
C1229 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t12 GNDA 0.04571f
C1230 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n0 GNDA 0.09572f
C1231 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t9 GNDA 0.17177f
C1232 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t6 GNDA 0.17177f
C1233 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t3 GNDA 0.04571f
C1234 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t5 GNDA 0.04571f
C1235 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n1 GNDA 0.09572f
C1236 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t4 GNDA 0.17177f
C1237 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t13 GNDA 0.17177f
C1238 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t16 GNDA 0.04571f
C1239 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t14 GNDA 0.04571f
C1240 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n2 GNDA 0.09572f
C1241 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t7 GNDA 0.17177f
C1242 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t18 GNDA 0.17177f
C1243 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t17 GNDA 0.04571f
C1244 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t8 GNDA 0.04571f
C1245 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n3 GNDA 0.09572f
C1246 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t15 GNDA 0.17177f
C1247 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t19 GNDA 0.17177f
C1248 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t20 GNDA 0.04571f
C1249 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t21 GNDA 0.04571f
C1250 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n4 GNDA 0.09572f
C1251 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t22 GNDA 0.21282f
C1252 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n5 GNDA 0.8214f
C1253 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n6 GNDA 0.42217f
C1254 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n7 GNDA 0.53295f
C1255 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n8 GNDA 0.46949f
C1256 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n9 GNDA 0.42217f
C1257 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n10 GNDA 0.53295f
C1258 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n11 GNDA 0.46949f
C1259 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n12 GNDA 0.42217f
C1260 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n13 GNDA 0.53295f
C1261 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n14 GNDA 0.46949f
C1262 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n15 GNDA 0.42217f
C1263 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n16 GNDA 0.53295f
C1264 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n17 GNDA 0.46949f
C1265 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n18 GNDA 1.09712f
C1266 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n19 GNDA 1.35128f
C1267 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t0 GNDA 0.11063f
C1268 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t23 GNDA 0.02438f
C1269 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t25 GNDA 0.02438f
C1270 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n20 GNDA 0.05278f
C1271 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t2 GNDA 0.02438f
C1272 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t24 GNDA 0.02438f
C1273 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n21 GNDA 0.05278f
C1274 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t27 GNDA 0.02438f
C1275 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.t26 GNDA 0.02438f
C1276 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n22 GNDA 0.05805f
C1277 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n23 GNDA 0.63042f
C1278 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n24 GNDA 0.57189f
C1279 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB.n25 GNDA 0.8575f
C1280 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t5 GNDA 0.01854f
C1281 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t2 GNDA 0.01854f
C1282 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n0 GNDA 0.04396f
C1283 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t0 GNDA 0.01854f
C1284 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t4 GNDA 0.01854f
C1285 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n1 GNDA 0.04396f
C1286 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t9 GNDA 0.01854f
C1287 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t1 GNDA 0.01854f
C1288 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n2 GNDA 0.04396f
C1289 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n3 GNDA 0.25242f
C1290 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t6 GNDA 0.07589f
C1291 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t7 GNDA 0.0695f
C1292 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n4 GNDA 1.46047f
C1293 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n5 GNDA 0.06518f
C1294 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n6 GNDA 0.13765f
C1295 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t3 GNDA 0.01854f
C1296 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.t8 GNDA 0.01854f
C1297 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD.n7 GNDA 0.04373f
C1298 P_IN[2].t7 GNDA 0.89992f
C1299 P_IN[2].t3 GNDA 0.89431f
C1300 P_IN[2].n0 GNDA 1.38976f
C1301 P_IN[2].t0 GNDA 0.36767f
C1302 P_IN[2].t2 GNDA 0.3659f
C1303 P_IN[2].n1 GNDA 0.97175f
C1304 P_IN[2].t6 GNDA 0.37373f
C1305 P_IN[2].t1 GNDA 0.36742f
C1306 P_IN[2].n2 GNDA 1.0824f
C1307 P_IN[2].n3 GNDA 0.52564f
C1308 P_IN[2].n4 GNDA 1.73661f
C1309 P_IN[2].t4 GNDA 0.89491f
C1310 P_IN[2].t5 GNDA 0.89327f
C1311 P_IN[2].n5 GNDA 1.15223f
C1312 P_IN[2].n6 GNDA 0.32559f
C1313 a_n11789_1598.t23 GNDA 0.02477f
C1314 a_n11789_1598.t17 GNDA 0.02477f
C1315 a_n11789_1598.n0 GNDA 0.05745f
C1316 a_n11789_1598.t18 GNDA 0.02477f
C1317 a_n11789_1598.t21 GNDA 0.02477f
C1318 a_n11789_1598.n1 GNDA 0.05745f
C1319 a_n11789_1598.n2 GNDA 0.42255f
C1320 a_n11789_1598.t20 GNDA 0.02477f
C1321 a_n11789_1598.t16 GNDA 0.02477f
C1322 a_n11789_1598.n3 GNDA 0.05745f
C1323 a_n11789_1598.t22 GNDA 0.02477f
C1324 a_n11789_1598.t19 GNDA 0.02477f
C1325 a_n11789_1598.n4 GNDA 0.05745f
C1326 a_n11789_1598.n5 GNDA 0.42255f
C1327 a_n11789_1598.n6 GNDA 0.12609f
C1328 a_n11789_1598.t13 GNDA 0.05554f
C1329 a_n11789_1598.t4 GNDA 0.05553f
C1330 a_n11789_1598.n7 GNDA 0.75856f
C1331 a_n11789_1598.n8 GNDA 0.61998f
C1332 a_n11789_1598.t0 GNDA 0.05546f
C1333 a_n11789_1598.n9 GNDA 0.2593f
C1334 a_n11789_1598.t5 GNDA 0.05546f
C1335 a_n11789_1598.n10 GNDA 0.2593f
C1336 a_n11789_1598.n11 GNDA 0.39892f
C1337 a_n11789_1598.n12 GNDA 0.39892f
C1338 a_n11789_1598.t1 GNDA 0.05546f
C1339 a_n11789_1598.n13 GNDA 0.2593f
C1340 a_n11789_1598.t10 GNDA 0.05546f
C1341 a_n11789_1598.n14 GNDA 0.2593f
C1342 a_n11789_1598.n15 GNDA 0.39892f
C1343 a_n11789_1598.n16 GNDA 0.37714f
C1344 a_n11789_1598.t3 GNDA 0.05546f
C1345 a_n11789_1598.n17 GNDA 0.2593f
C1346 a_n11789_1598.t11 GNDA 0.05546f
C1347 a_n11789_1598.n18 GNDA 0.26103f
C1348 a_n11789_1598.n19 GNDA 0.08229f
C1349 a_n11789_1598.n20 GNDA 1.80716f
C1350 a_n11789_1598.n21 GNDA 0.58376f
C1351 a_n11789_1598.t12 GNDA 0.05546f
C1352 a_n11789_1598.n22 GNDA 0.2593f
C1353 a_n11789_1598.t14 GNDA 0.05546f
C1354 a_n11789_1598.n23 GNDA 0.2593f
C1355 a_n11789_1598.n24 GNDA 0.39892f
C1356 a_n11789_1598.n25 GNDA 0.39892f
C1357 a_n11789_1598.t2 GNDA 0.05546f
C1358 a_n11789_1598.n26 GNDA 0.2593f
C1359 a_n11789_1598.t9 GNDA 0.05546f
C1360 a_n11789_1598.n27 GNDA 0.2593f
C1361 a_n11789_1598.n28 GNDA 0.39892f
C1362 a_n11789_1598.n29 GNDA 0.39892f
C1363 a_n11789_1598.t6 GNDA 0.05546f
C1364 a_n11789_1598.n30 GNDA 0.2593f
C1365 a_n11789_1598.t7 GNDA 0.05546f
C1366 a_n11789_1598.n31 GNDA 0.2593f
C1367 a_n11789_1598.n32 GNDA 0.61998f
C1368 a_n11789_1598.t8 GNDA 0.05553f
C1369 a_n11789_1598.n33 GNDA 0.75856f
C1370 a_n11789_1598.t15 GNDA 0.05554f
C1371 opa_folded_cascode_0.monticelli_top_0.A.t2 GNDA 0.33267f
C1372 opa_folded_cascode_0.monticelli_top_0.A.t1 GNDA 0.44805f
C1373 opa_folded_cascode_0.monticelli_top_0.A.n0 GNDA 1.42513f
C1374 opa_folded_cascode_0.monticelli_top_0.A.t3 GNDA 0.45415f
C1375 opa_folded_cascode_0.monticelli_top_0.A.n1 GNDA 1.80267f
C1376 opa_folded_cascode_0.monticelli_top_0.A.t0 GNDA 0.33485f
C1377 opa_folded_cascode_0.monticelli_top_0.A.n2 GNDA 1.63869f
C1378 opa_folded_cascode_0.monticelli_top_0.A.t7 GNDA 0.70113f
C1379 opa_folded_cascode_0.monticelli_top_0.A.t6 GNDA 0.70026f
C1380 opa_folded_cascode_0.monticelli_top_0.A.n3 GNDA 0.57805f
C1381 opa_folded_cascode_0.monticelli_top_0.A.t9 GNDA 0.70113f
C1382 opa_folded_cascode_0.monticelli_top_0.A.t8 GNDA 0.70026f
C1383 opa_folded_cascode_0.monticelli_top_0.A.n4 GNDA 0.57843f
C1384 opa_folded_cascode_0.monticelli_top_0.A.n5 GNDA 0.37163f
C1385 opa_folded_cascode_0.monticelli_top_0.A.n6 GNDA 0.43001f
C1386 opa_folded_cascode_0.monticelli_top_0.A.t5 GNDA 0.10488f
C1387 opa_folded_cascode_0.monticelli_top_0.A.t4 GNDA 0.1592f
C1388 opa_folded_cascode_0.monticelli_top_0.A.n7 GNDA 1.27842f
C1389 opa_folded_cascode_0.VB2.t10 GNDA 0.39693f
C1390 opa_folded_cascode_0.VB2.t0 GNDA 0.11669f
C1391 opa_folded_cascode_0.VB2.t4 GNDA 0.11669f
C1392 opa_folded_cascode_0.VB2.n0 GNDA 1.17006f
C1393 opa_folded_cascode_0.VB2.t5 GNDA 0.11669f
C1394 opa_folded_cascode_0.VB2.t1 GNDA 0.11669f
C1395 opa_folded_cascode_0.VB2.n1 GNDA 0.48525f
C1396 opa_folded_cascode_0.VB2.n2 GNDA 1.72063f
C1397 opa_folded_cascode_0.VB2.t7 GNDA 0.11669f
C1398 opa_folded_cascode_0.VB2.t2 GNDA 0.11669f
C1399 opa_folded_cascode_0.VB2.n3 GNDA 1.17107f
C1400 opa_folded_cascode_0.VB2.t3 GNDA 0.11669f
C1401 opa_folded_cascode_0.VB2.t6 GNDA 0.11669f
C1402 opa_folded_cascode_0.VB2.n4 GNDA 0.48425f
C1403 opa_folded_cascode_0.VB2.n5 GNDA 1.8498f
C1404 opa_folded_cascode_0.VB2.n6 GNDA 3.18521f
C1405 opa_folded_cascode_0.VB2.t12 GNDA 0.40061f
C1406 opa_folded_cascode_0.VB2.t14 GNDA 0.3992f
C1407 opa_folded_cascode_0.VB2.n7 GNDA 0.64417f
C1408 opa_folded_cascode_0.VB2.t13 GNDA 0.40061f
C1409 opa_folded_cascode_0.VB2.t15 GNDA 0.3992f
C1410 opa_folded_cascode_0.VB2.n8 GNDA 0.63961f
C1411 opa_folded_cascode_0.VB2.n9 GNDA 3.47383f
C1412 opa_folded_cascode_0.VB2.n10 GNDA 0.24736f
C1413 opa_folded_cascode_0.VB2.t8 GNDA 0.3978f
C1414 opa_folded_cascode_0.VB2.t9 GNDA 0.10005f
C1415 opa_folded_cascode_0.VB2.n11 GNDA 0.45496f
C1416 opa_folded_cascode_0.VB2.t11 GNDA 0.10005f
C1417 opa_folded_cascode_0.VB2.n12 GNDA 0.25966f
C1418 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t15 GNDA 0.02428f
C1419 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t16 GNDA 0.02428f
C1420 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n0 GNDA 0.05333f
C1421 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t18 GNDA 0.08653f
C1422 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t10 GNDA 0.02428f
C1423 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t7 GNDA 0.02428f
C1424 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n1 GNDA 0.05333f
C1425 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t6 GNDA 0.08653f
C1426 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t19 GNDA 0.02428f
C1427 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t5 GNDA 0.02428f
C1428 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n2 GNDA 0.05333f
C1429 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t8 GNDA 0.08653f
C1430 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t21 GNDA 0.52705f
C1431 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t23 GNDA 0.46697f
C1432 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t20 GNDA 0.44522f
C1433 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n3 GNDA 2.3024f
C1434 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t22 GNDA 0.52635f
C1435 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n4 GNDA 1.50121f
C1436 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n5 GNDA 3.10193f
C1437 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n6 GNDA 2.17073f
C1438 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n7 GNDA 0.34173f
C1439 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n8 GNDA 0.511f
C1440 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t9 GNDA 0.08653f
C1441 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n9 GNDA 0.42483f
C1442 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n10 GNDA 0.33613f
C1443 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n11 GNDA 0.34173f
C1444 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n12 GNDA 0.511f
C1445 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t4 GNDA 0.08653f
C1446 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n13 GNDA 0.42483f
C1447 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n14 GNDA 0.33613f
C1448 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n15 GNDA 0.34173f
C1449 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n16 GNDA 0.511f
C1450 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t17 GNDA 0.08653f
C1451 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n17 GNDA 0.42483f
C1452 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t2 GNDA 0.08653f
C1453 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t1 GNDA 0.02428f
C1454 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t3 GNDA 0.02428f
C1455 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n18 GNDA 0.05333f
C1456 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t0 GNDA 0.08653f
C1457 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t13 GNDA 0.08653f
C1458 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t14 GNDA 0.02428f
C1459 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t11 GNDA 0.02428f
C1460 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n19 GNDA 0.05333f
C1461 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.t12 GNDA 0.12342f
C1462 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n20 GNDA 0.8221f
C1463 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n21 GNDA 0.31986f
C1464 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n22 GNDA 0.33613f
C1465 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n23 GNDA 0.42483f
C1466 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n24 GNDA 0.511f
C1467 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n25 GNDA 0.34173f
C1468 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB.n26 GNDA 0.33613f
C1469 N_IN.n0 GNDA 0.32968f
C1470 N_IN.t1 GNDA 0.70518f
C1471 N_IN.n1 GNDA 0.37997f
C1472 N_IN.t19 GNDA 0.70518f
C1473 N_IN.n2 GNDA 0.68365f
C1474 N_IN.t39 GNDA 0.29005f
C1475 N_IN.n3 GNDA 0.585f
C1476 N_IN.t7 GNDA 0.28885f
C1477 N_IN.n4 GNDA 0.35254f
C1478 N_IN.t25 GNDA 0.29005f
C1479 N_IN.n5 GNDA 0.39393f
C1480 N_IN.t28 GNDA 0.29005f
C1481 N_IN.n6 GNDA 0.4639f
C1482 N_IN.t5 GNDA 0.28885f
C1483 N_IN.n7 GNDA 0.28257f
C1484 N_IN.t31 GNDA 0.28885f
C1485 N_IN.n8 GNDA 0.35254f
C1486 N_IN.t15 GNDA 0.29005f
C1487 N_IN.n9 GNDA 0.39393f
C1488 N_IN.t29 GNDA 0.29005f
C1489 N_IN.n10 GNDA 0.4639f
C1490 N_IN.t9 GNDA 0.28885f
C1491 N_IN.n11 GNDA 0.28257f
C1492 N_IN.t35 GNDA 0.29005f
C1493 N_IN.n12 GNDA 0.69416f
C1494 N_IN.t37 GNDA 0.28885f
C1495 N_IN.n13 GNDA 0.6023f
C1496 N_IN.t38 GNDA 0.28885f
C1497 N_IN.n14 GNDA 0.35254f
C1498 N_IN.n15 GNDA 0.46348f
C1499 N_IN.n16 GNDA 0.36114f
C1500 N_IN.t22 GNDA 0.29005f
C1501 N_IN.n17 GNDA 0.39393f
C1502 N_IN.t32 GNDA 0.29005f
C1503 N_IN.n18 GNDA 0.4639f
C1504 N_IN.n19 GNDA 0.36114f
C1505 N_IN.n20 GNDA 0.46348f
C1506 N_IN.t17 GNDA 0.28885f
C1507 N_IN.n21 GNDA 0.28257f
C1508 N_IN.t0 GNDA 0.28885f
C1509 N_IN.n22 GNDA 0.35254f
C1510 N_IN.n23 GNDA 0.46348f
C1511 N_IN.n24 GNDA 0.36114f
C1512 N_IN.t3 GNDA 0.29005f
C1513 N_IN.n25 GNDA 0.39393f
C1514 N_IN.t10 GNDA 0.29005f
C1515 N_IN.n26 GNDA 0.4639f
C1516 N_IN.n27 GNDA 0.36114f
C1517 N_IN.n28 GNDA 0.46348f
C1518 N_IN.t34 GNDA 0.28885f
C1519 N_IN.n29 GNDA 0.28257f
C1520 N_IN.t13 GNDA 0.28885f
C1521 N_IN.n30 GNDA 0.45601f
C1522 N_IN.n31 GNDA 0.42512f
C1523 N_IN.n32 GNDA 0.64866f
C1524 N_IN.t23 GNDA 0.706f
C1525 N_IN.n33 GNDA 0.63649f
C1526 N_IN.t33 GNDA 0.706f
C1527 N_IN.n34 GNDA 0.48998f
C1528 N_IN.t6 GNDA 0.706f
C1529 N_IN.n35 GNDA 0.55995f
C1530 N_IN.t14 GNDA 0.70518f
C1531 N_IN.n36 GNDA 0.44995f
C1532 N_IN.t12 GNDA 0.70518f
C1533 N_IN.n37 GNDA 0.37997f
C1534 N_IN.t36 GNDA 0.70518f
C1535 N_IN.n38 GNDA 0.44995f
C1536 N_IN.t27 GNDA 0.706f
C1537 N_IN.n39 GNDA 0.48998f
C1538 N_IN.t11 GNDA 0.706f
C1539 N_IN.n40 GNDA 0.55995f
C1540 N_IN.t16 GNDA 0.70518f
C1541 N_IN.n41 GNDA 0.37997f
C1542 N_IN.t20 GNDA 0.706f
C1543 N_IN.n42 GNDA 0.62591f
C1544 N_IN.t2 GNDA 0.70518f
C1545 N_IN.n43 GNDA 0.55128f
C1546 N_IN.t4 GNDA 0.70518f
C1547 N_IN.n44 GNDA 0.44995f
C1548 N_IN.n45 GNDA 0.32968f
C1549 N_IN.n46 GNDA 0.22719f
C1550 N_IN.t30 GNDA 0.706f
C1551 N_IN.n47 GNDA 0.48998f
C1552 N_IN.t18 GNDA 0.706f
C1553 N_IN.n48 GNDA 0.55995f
C1554 N_IN.n49 GNDA 0.22719f
C1555 N_IN.n50 GNDA 0.32968f
C1556 N_IN.t21 GNDA 0.70518f
C1557 N_IN.n51 GNDA 0.37997f
C1558 N_IN.t8 GNDA 0.70518f
C1559 N_IN.n52 GNDA 0.44995f
C1560 N_IN.n53 GNDA 0.32968f
C1561 N_IN.n54 GNDA 0.22719f
C1562 N_IN.t24 GNDA 0.706f
C1563 N_IN.n55 GNDA 0.48998f
C1564 N_IN.t26 GNDA 0.706f
C1565 N_IN.n56 GNDA 0.55995f
C1566 N_IN.n57 GNDA 0.22719f
C1567 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t1 GNDA 0.01191f
C1568 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t9 GNDA 0.01191f
C1569 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n0 GNDA 0.02616f
C1570 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t0 GNDA 0.04245f
C1571 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t5 GNDA 0.01191f
C1572 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t13 GNDA 0.01191f
C1573 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n1 GNDA 0.02616f
C1574 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t17 GNDA 0.04245f
C1575 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t18 GNDA 0.01191f
C1576 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t12 GNDA 0.01191f
C1577 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n2 GNDA 0.02616f
C1578 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t11 GNDA 0.04245f
C1579 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t16 GNDA 0.01191f
C1580 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t3 GNDA 0.01191f
C1581 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n3 GNDA 0.02616f
C1582 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t23 GNDA 0.04245f
C1583 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t15 GNDA 0.26016f
C1584 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t14 GNDA 0.26166f
C1585 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t21 GNDA 0.21835f
C1586 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t20 GNDA 0.29634f
C1587 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n4 GNDA 1.07628f
C1588 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n5 GNDA 0.67911f
C1589 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n6 GNDA 1.21166f
C1590 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t26 GNDA 0.78859f
C1591 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t28 GNDA 0.89044f
C1592 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t34 GNDA 0.65724f
C1593 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n7 GNDA 0.85404f
C1594 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t39 GNDA 0.65724f
C1595 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n8 GNDA 0.5153f
C1596 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n9 GNDA 0.46821f
C1597 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t37 GNDA 0.78859f
C1598 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t40 GNDA 0.89044f
C1599 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t27 GNDA 0.65724f
C1600 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n10 GNDA 0.85404f
C1601 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t32 GNDA 0.65724f
C1602 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n11 GNDA 0.5153f
C1603 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n12 GNDA 0.44059f
C1604 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n13 GNDA 0.46078f
C1605 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t41 GNDA 0.78859f
C1606 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t43 GNDA 0.89044f
C1607 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t29 GNDA 0.65724f
C1608 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n14 GNDA 0.85404f
C1609 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t35 GNDA 0.65724f
C1610 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n15 GNDA 0.5153f
C1611 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n16 GNDA 0.46836f
C1612 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t42 GNDA 0.78859f
C1613 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t25 GNDA 0.89044f
C1614 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t31 GNDA 0.65724f
C1615 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n17 GNDA 0.85404f
C1616 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t36 GNDA 0.65724f
C1617 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n18 GNDA 0.5153f
C1618 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n19 GNDA 0.44059f
C1619 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n20 GNDA 0.59017f
C1620 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t30 GNDA 0.78859f
C1621 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t33 GNDA 0.89044f
C1622 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t38 GNDA 0.65724f
C1623 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n21 GNDA 0.85404f
C1624 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t24 GNDA 0.65724f
C1625 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n22 GNDA 0.5153f
C1626 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n23 GNDA 0.44059f
C1627 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n24 GNDA 0.3281f
C1628 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n25 GNDA 1.89782f
C1629 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n26 GNDA 1.7696f
C1630 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n27 GNDA 0.30404f
C1631 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n28 GNDA 0.1836f
C1632 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n29 GNDA 0.25007f
C1633 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t6 GNDA 0.04245f
C1634 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n30 GNDA 0.19307f
C1635 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n31 GNDA 0.1649f
C1636 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n32 GNDA 0.1836f
C1637 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n33 GNDA 0.25007f
C1638 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t10 GNDA 0.04245f
C1639 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n34 GNDA 0.19307f
C1640 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n35 GNDA 0.1649f
C1641 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n36 GNDA 0.1836f
C1642 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n37 GNDA 0.25007f
C1643 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t8 GNDA 0.04245f
C1644 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n38 GNDA 0.19307f
C1645 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n39 GNDA 0.1649f
C1646 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n40 GNDA 0.1836f
C1647 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n41 GNDA 0.24032f
C1648 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t2 GNDA 0.04245f
C1649 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n42 GNDA 0.19049f
C1650 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t22 GNDA 0.04245f
C1651 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t4 GNDA 0.01191f
C1652 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t19 GNDA 0.01191f
C1653 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n43 GNDA 0.02616f
C1654 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.t7 GNDA 0.04448f
C1655 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n44 GNDA 0.39269f
C1656 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n45 GNDA 0.1836f
C1657 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA.n46 GNDA 0.1649f
C1658 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t11 GNDA 0.08659f
C1659 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t2 GNDA 0.08376f
C1660 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n0 GNDA 1.26472f
C1661 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t12 GNDA 0.08376f
C1662 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n1 GNDA 0.63996f
C1663 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t5 GNDA 0.08659f
C1664 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t1 GNDA 0.08376f
C1665 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n2 GNDA 1.26472f
C1666 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t4 GNDA 0.08376f
C1667 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n3 GNDA 0.77891f
C1668 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t13 GNDA 0.08376f
C1669 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n4 GNDA 0.77891f
C1670 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t3 GNDA 0.08376f
C1671 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n5 GNDA 0.68725f
C1672 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n6 GNDA 0.54086f
C1673 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t15 GNDA 0.08659f
C1674 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t6 GNDA 0.08376f
C1675 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n7 GNDA 1.26472f
C1676 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t9 GNDA 0.08376f
C1677 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n8 GNDA 0.77891f
C1678 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t8 GNDA 0.08376f
C1679 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n9 GNDA 0.59704f
C1680 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t10 GNDA 0.08659f
C1681 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t14 GNDA 0.08376f
C1682 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n10 GNDA 1.26472f
C1683 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t0 GNDA 0.08376f
C1684 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n11 GNDA 0.77891f
C1685 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t7 GNDA 0.08376f
C1686 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n12 GNDA 0.64432f
C1687 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n13 GNDA 0.31646f
C1688 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n14 GNDA 1.724f
C1689 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t19 GNDA 0.07878f
C1690 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t28 GNDA 0.07878f
C1691 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n15 GNDA 0.5907f
C1692 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t27 GNDA 0.07878f
C1693 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t25 GNDA 0.07878f
C1694 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n16 GNDA 0.35538f
C1695 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n17 GNDA 1.13493f
C1696 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t18 GNDA 0.07878f
C1697 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t30 GNDA 0.07878f
C1698 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n18 GNDA 0.5907f
C1699 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t29 GNDA 0.07878f
C1700 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t21 GNDA 0.07878f
C1701 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n19 GNDA 0.35538f
C1702 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n20 GNDA 1.18222f
C1703 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n21 GNDA 0.65639f
C1704 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t20 GNDA 0.07878f
C1705 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t17 GNDA 0.07878f
C1706 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n22 GNDA 0.57514f
C1707 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t23 GNDA 0.07878f
C1708 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t16 GNDA 0.07878f
C1709 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n23 GNDA 0.5907f
C1710 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t31 GNDA 0.07878f
C1711 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t24 GNDA 0.07878f
C1712 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n24 GNDA 0.35538f
C1713 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n25 GNDA 1.43212f
C1714 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t22 GNDA 0.07878f
C1715 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.t26 GNDA 0.07878f
C1716 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n26 GNDA 0.35538f
C1717 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n27 GNDA 0.57073f
C1718 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n28 GNDA 0.87695f
C1719 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4.n29 GNDA 1.05186f
C1720 opa_folded_cascode_0.monticelli_top_0.B.t2 GNDA 0.33786f
C1721 opa_folded_cascode_0.monticelli_top_0.B.t3 GNDA 0.35366f
C1722 opa_folded_cascode_0.monticelli_top_0.B.n0 GNDA 1.69903f
C1723 opa_folded_cascode_0.monticelli_top_0.B.t1 GNDA 0.10661f
C1724 opa_folded_cascode_0.monticelli_top_0.B.t0 GNDA 0.1615f
C1725 opa_folded_cascode_0.monticelli_top_0.B.n1 GNDA 0.80656f
C1726 opa_folded_cascode_0.monticelli_top_0.B.t4 GNDA 0.16175f
C1727 opa_folded_cascode_0.monticelli_top_0.B.n2 GNDA 1.08345f
C1728 opa_folded_cascode_0.monticelli_top_0.B.t5 GNDA 0.1574f
C1729 opa_folded_cascode_0.monticelli_top_0.B.n3 GNDA 0.91132f
C1730 opa_folded_cascode_0.monticelli_top_0.B.t6 GNDA 0.29079f
C1731 opa_folded_cascode_0.monticelli_top_0.B.t9 GNDA 0.29006f
C1732 opa_folded_cascode_0.monticelli_top_0.B.n4 GNDA 0.31276f
C1733 opa_folded_cascode_0.monticelli_top_0.B.t8 GNDA 0.29079f
C1734 opa_folded_cascode_0.monticelli_top_0.B.t7 GNDA 0.29006f
C1735 opa_folded_cascode_0.monticelli_top_0.B.n5 GNDA 0.31276f
C1736 opa_folded_cascode_0.monticelli_top_0.B.n6 GNDA 0.20481f
C1737 opa_folded_cascode_0.monticelli_top_0.B.n7 GNDA 0.56015f
C1738 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t0 GNDA 0.2583f
C1739 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t9 GNDA 0.23142f
C1740 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t1 GNDA 0.23142f
C1741 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n0 GNDA 1.02719f
C1742 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n1 GNDA 1.97426f
C1743 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t13 GNDA 0.24661f
C1744 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t6 GNDA 0.23142f
C1745 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t7 GNDA 0.23142f
C1746 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n2 GNDA 1.02719f
C1747 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n3 GNDA 1.33348f
C1748 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t3 GNDA 0.23136f
C1749 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t5 GNDA 0.23136f
C1750 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n4 GNDA 0.73738f
C1751 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n5 GNDA 1.24044f
C1752 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n6 GNDA 1.40802f
C1753 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t10 GNDA 0.24661f
C1754 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t12 GNDA 0.23142f
C1755 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t2 GNDA 0.23142f
C1756 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n7 GNDA 1.02719f
C1757 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n8 GNDA 1.33348f
C1758 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t11 GNDA 0.23136f
C1759 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t4 GNDA 0.23136f
C1760 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n9 GNDA 0.73738f
C1761 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n10 GNDA 0.92337f
C1762 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t8 GNDA 0.2583f
C1763 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t14 GNDA 0.23142f
C1764 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t15 GNDA 0.23142f
C1765 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n11 GNDA 1.02719f
C1766 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n12 GNDA 2.29133f
C1767 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n13 GNDA 1.35167f
C1768 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n14 GNDA 0.94014f
C1769 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t20 GNDA 0.2335f
C1770 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t25 GNDA 0.23352f
C1771 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n15 GNDA 1.21388f
C1772 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t29 GNDA 0.2503f
C1773 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n16 GNDA 1.2622f
C1774 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t19 GNDA 0.2503f
C1775 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n17 GNDA 1.05359f
C1776 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t17 GNDA 0.2503f
C1777 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n18 GNDA 1.01045f
C1778 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t26 GNDA 0.26105f
C1779 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t16 GNDA 0.2503f
C1780 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n19 GNDA 1.89151f
C1781 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t31 GNDA 0.2503f
C1782 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n20 GNDA 1.59785f
C1783 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n21 GNDA 1.13336f
C1784 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t23 GNDA 0.26105f
C1785 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t27 GNDA 0.2503f
C1786 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n22 GNDA 1.89151f
C1787 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t18 GNDA 0.2503f
C1788 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n23 GNDA 1.28078f
C1789 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t24 GNDA 0.23352f
C1790 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t28 GNDA 0.2335f
C1791 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n24 GNDA 1.21388f
C1792 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t30 GNDA 0.2503f
C1793 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n25 GNDA 1.2622f
C1794 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t21 GNDA 0.2503f
C1795 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n26 GNDA 1.05359f
C1796 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.t22 GNDA 0.2503f
C1797 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n27 GNDA 1.32752f
C1798 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n28 GNDA 1.12088f
C1799 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4.n29 GNDA 0.89148f
C1800 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t19 GNDA 0.08748f
C1801 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t4 GNDA 0.08248f
C1802 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t10 GNDA 0.07822f
C1803 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n0 GNDA 1.08605f
C1804 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t9 GNDA 0.07822f
C1805 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n1 GNDA 0.46201f
C1806 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n2 GNDA 1.08984f
C1807 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t0 GNDA 0.0844f
C1808 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n3 GNDA 0.82131f
C1809 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t12 GNDA 0.0844f
C1810 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n4 GNDA 0.82131f
C1811 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t8 GNDA 0.0844f
C1812 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n5 GNDA 0.68473f
C1813 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t18 GNDA 0.08748f
C1814 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t7 GNDA 0.0844f
C1815 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n6 GNDA 1.3512f
C1816 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t13 GNDA 0.0844f
C1817 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n7 GNDA 0.72881f
C1818 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n8 GNDA 0.57528f
C1819 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t1 GNDA 0.08748f
C1820 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t17 GNDA 0.0844f
C1821 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n9 GNDA 1.3512f
C1822 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t2 GNDA 0.0844f
C1823 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n10 GNDA 0.82131f
C1824 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t11 GNDA 0.0844f
C1825 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n11 GNDA 0.64209f
C1826 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t16 GNDA 0.08748f
C1827 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t14 GNDA 0.08248f
C1828 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t3 GNDA 0.07822f
C1829 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n12 GNDA 1.08605f
C1830 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t5 GNDA 0.07822f
C1831 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n13 GNDA 0.46201f
C1832 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n14 GNDA 1.08984f
C1833 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t6 GNDA 0.0844f
C1834 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n15 GNDA 0.82131f
C1835 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t15 GNDA 0.0844f
C1836 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n16 GNDA 0.68617f
C1837 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n17 GNDA 0.31437f
C1838 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n18 GNDA 1.77552f
C1839 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t31 GNDA 0.07826f
C1840 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t32 GNDA 0.07826f
C1841 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n19 GNDA 0.70457f
C1842 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t39 GNDA 0.07826f
C1843 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t24 GNDA 0.07826f
C1844 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n20 GNDA 0.47705f
C1845 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n21 GNDA 1.14431f
C1846 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t21 GNDA 0.07832f
C1847 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t25 GNDA 0.07822f
C1848 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n22 GNDA 0.41842f
C1849 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t22 GNDA 0.07822f
C1850 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n23 GNDA 0.19934f
C1851 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t36 GNDA 0.07826f
C1852 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n24 GNDA 0.57069f
C1853 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t37 GNDA 0.07826f
C1854 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t23 GNDA 0.07826f
C1855 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n25 GNDA 0.47705f
C1856 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n26 GNDA 1.18839f
C1857 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n27 GNDA 0.71001f
C1858 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t33 GNDA 0.07826f
C1859 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t28 GNDA 0.07832f
C1860 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t20 GNDA 0.07822f
C1861 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n28 GNDA 0.41842f
C1862 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t27 GNDA 0.07822f
C1863 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n29 GNDA 0.19934f
C1864 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n30 GNDA 0.57069f
C1865 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t26 GNDA 0.07826f
C1866 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t29 GNDA 0.07826f
C1867 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n31 GNDA 0.47705f
C1868 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n32 GNDA 1.41604f
C1869 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t34 GNDA 0.07826f
C1870 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t35 GNDA 0.07826f
C1871 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n33 GNDA 0.70457f
C1872 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t30 GNDA 0.07826f
C1873 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.t38 GNDA 0.07826f
C1874 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n34 GNDA 0.47705f
C1875 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n35 GNDA 0.91667f
C1876 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n36 GNDA 0.54346f
C1877 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0.n37 GNDA 1.19678f
C1878 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t9 GNDA 0.03763f
C1879 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t2 GNDA 0.03762f
C1880 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t10 GNDA 0.03758f
C1881 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n0 GNDA 0.26539f
C1882 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t15 GNDA 0.03758f
C1883 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n1 GNDA 0.29049f
C1884 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n2 GNDA 0.35844f
C1885 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n3 GNDA 0.43211f
C1886 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t4 GNDA 0.03758f
C1887 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n4 GNDA 0.19468f
C1888 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t16 GNDA 0.03758f
C1889 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n5 GNDA 0.19468f
C1890 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n6 GNDA 0.27467f
C1891 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n7 GNDA 0.27467f
C1892 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t14 GNDA 0.03758f
C1893 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n8 GNDA 0.19468f
C1894 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t17 GNDA 0.03758f
C1895 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n9 GNDA 0.19468f
C1896 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n10 GNDA 0.03513f
C1897 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t1 GNDA 0.03763f
C1898 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t8 GNDA 0.03763f
C1899 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n11 GNDA 0.55219f
C1900 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n12 GNDA 0.60467f
C1901 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t7 GNDA 0.03763f
C1902 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t5 GNDA 0.03763f
C1903 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n13 GNDA 0.55306f
C1904 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n14 GNDA 0.43211f
C1905 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t12 GNDA 0.03758f
C1906 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n15 GNDA 0.19468f
C1907 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t3 GNDA 0.03758f
C1908 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n16 GNDA 0.19468f
C1909 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n17 GNDA 0.16566f
C1910 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t6 GNDA 0.03763f
C1911 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t13 GNDA 0.03762f
C1912 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t18 GNDA 0.03758f
C1913 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n18 GNDA 0.26539f
C1914 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t11 GNDA 0.03758f
C1915 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n19 GNDA 0.29049f
C1916 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n20 GNDA 0.35844f
C1917 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n21 GNDA 0.43211f
C1918 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t0 GNDA 0.03758f
C1919 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n22 GNDA 0.19468f
C1920 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t19 GNDA 0.03758f
C1921 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n23 GNDA 0.19468f
C1922 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n24 GNDA 0.1431f
C1923 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n25 GNDA 0.24058f
C1924 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n26 GNDA 0.91514f
C1925 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n27 GNDA 0.18865f
C1926 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t72 GNDA 0.1893f
C1927 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t33 GNDA 0.18766f
C1928 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n28 GNDA 0.46608f
C1929 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t67 GNDA 0.18766f
C1930 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n29 GNDA 0.23386f
C1931 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t77 GNDA 0.18766f
C1932 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n30 GNDA 0.23386f
C1933 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t34 GNDA 0.18766f
C1934 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n31 GNDA 0.23386f
C1935 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t46 GNDA 0.18766f
C1936 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n32 GNDA 0.23386f
C1937 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t62 GNDA 0.18766f
C1938 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n33 GNDA 0.23386f
C1939 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t39 GNDA 0.18766f
C1940 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n34 GNDA 0.23386f
C1941 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t30 GNDA 0.18766f
C1942 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n35 GNDA 0.21251f
C1943 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t21 GNDA 0.03764f
C1944 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t20 GNDA 0.14431f
C1945 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n36 GNDA 3.02766f
C1946 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n37 GNDA 0.32533f
C1947 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t69 GNDA 0.19022f
C1948 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t44 GNDA 0.18766f
C1949 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n38 GNDA 0.5957f
C1950 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t51 GNDA 0.18766f
C1951 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n39 GNDA 0.23386f
C1952 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t70 GNDA 0.18766f
C1953 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n40 GNDA 0.23386f
C1954 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t80 GNDA 0.18766f
C1955 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n41 GNDA 0.23386f
C1956 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t41 GNDA 0.18766f
C1957 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n42 GNDA 0.23386f
C1958 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t73 GNDA 0.18766f
C1959 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n43 GNDA 0.23386f
C1960 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t66 GNDA 0.18766f
C1961 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n44 GNDA 0.21251f
C1962 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t74 GNDA 0.1893f
C1963 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t35 GNDA 0.18766f
C1964 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n45 GNDA 0.46608f
C1965 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t68 GNDA 0.18766f
C1966 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n46 GNDA 0.23386f
C1967 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t78 GNDA 0.18766f
C1968 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n47 GNDA 0.23386f
C1969 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t36 GNDA 0.18766f
C1970 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n48 GNDA 0.23386f
C1971 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t47 GNDA 0.18766f
C1972 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n49 GNDA 0.23386f
C1973 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t64 GNDA 0.18766f
C1974 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n50 GNDA 0.23386f
C1975 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t40 GNDA 0.18766f
C1976 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n51 GNDA 0.23386f
C1977 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t31 GNDA 0.18766f
C1978 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n52 GNDA 0.21251f
C1979 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t81 GNDA 0.18766f
C1980 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n53 GNDA 0.35069f
C1981 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t59 GNDA 0.18766f
C1982 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n54 GNDA 0.23386f
C1983 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t27 GNDA 0.18766f
C1984 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n55 GNDA 0.23386f
C1985 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t76 GNDA 0.18766f
C1986 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n56 GNDA 0.23386f
C1987 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t58 GNDA 0.18766f
C1988 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n57 GNDA 0.23386f
C1989 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t23 GNDA 0.18766f
C1990 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n58 GNDA 0.23386f
C1991 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t65 GNDA 0.18766f
C1992 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n59 GNDA 0.18995f
C1993 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n60 GNDA 0.0734f
C1994 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n61 GNDA 0.27713f
C1995 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n62 GNDA 0.06527f
C1996 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t42 GNDA 0.18766f
C1997 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n63 GNDA 0.18995f
C1998 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t55 GNDA 0.18766f
C1999 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n64 GNDA 0.23386f
C2000 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t37 GNDA 0.18766f
C2001 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n65 GNDA 0.23386f
C2002 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t49 GNDA 0.18766f
C2003 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n66 GNDA 0.23386f
C2004 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t60 GNDA 0.18766f
C2005 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n67 GNDA 0.23386f
C2006 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t38 GNDA 0.18766f
C2007 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n68 GNDA 0.44501f
C2008 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n69 GNDA 0.25344f
C2009 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t53 GNDA 0.19022f
C2010 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t32 GNDA 0.18766f
C2011 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n70 GNDA 0.5957f
C2012 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t45 GNDA 0.18766f
C2013 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n71 GNDA 0.23386f
C2014 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t54 GNDA 0.18766f
C2015 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n72 GNDA 0.23386f
C2016 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t71 GNDA 0.18766f
C2017 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n73 GNDA 0.23386f
C2018 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t28 GNDA 0.18766f
C2019 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n74 GNDA 0.23386f
C2020 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t61 GNDA 0.18766f
C2021 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n75 GNDA 0.23386f
C2022 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t52 GNDA 0.18766f
C2023 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n76 GNDA 0.21251f
C2024 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n77 GNDA 0.06527f
C2025 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t29 GNDA 0.18766f
C2026 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n78 GNDA 0.18995f
C2027 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t48 GNDA 0.18766f
C2028 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n79 GNDA 0.23386f
C2029 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t24 GNDA 0.18766f
C2030 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n80 GNDA 0.23386f
C2031 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t43 GNDA 0.18766f
C2032 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n81 GNDA 0.23386f
C2033 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t50 GNDA 0.18766f
C2034 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n82 GNDA 0.23386f
C2035 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t25 GNDA 0.18766f
C2036 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n83 GNDA 0.44501f
C2037 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n84 GNDA 0.3724f
C2038 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t79 GNDA 0.18766f
C2039 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n85 GNDA 0.35885f
C2040 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t57 GNDA 0.18766f
C2041 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n86 GNDA 0.23386f
C2042 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t26 GNDA 0.18766f
C2043 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n87 GNDA 0.23386f
C2044 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t75 GNDA 0.18766f
C2045 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n88 GNDA 0.23386f
C2046 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t56 GNDA 0.18766f
C2047 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n89 GNDA 0.23386f
C2048 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t22 GNDA 0.18766f
C2049 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n90 GNDA 0.23386f
C2050 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.t63 GNDA 0.18766f
C2051 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n91 GNDA 0.18995f
C2052 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n92 GNDA 0.06527f
C2053 opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1.n93 GNDA 0.1306f
C2054 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n0 GNDA 0.01746f
C2055 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n1 GNDA 0.0906f
C2056 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n2 GNDA 0.08269f
C2057 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n3 GNDA 0.08287f
C2058 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t4 GNDA 0.15492f
C2059 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t43 GNDA 0.15358f
C2060 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n4 GNDA 0.38143f
C2061 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t19 GNDA 0.15358f
C2062 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n5 GNDA 0.19139f
C2063 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t40 GNDA 0.15358f
C2064 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n6 GNDA 0.19139f
C2065 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t66 GNDA 0.15358f
C2066 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n7 GNDA 0.16326f
C2067 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t24 GNDA 0.15492f
C2068 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t46 GNDA 0.15358f
C2069 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n8 GNDA 0.38143f
C2070 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t6 GNDA 0.15358f
C2071 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n9 GNDA 0.19139f
C2072 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t47 GNDA 0.15358f
C2073 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n10 GNDA 0.19139f
C2074 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t26 GNDA 0.15358f
C2075 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n11 GNDA 0.19139f
C2076 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t58 GNDA 0.15358f
C2077 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n12 GNDA 0.19139f
C2078 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t25 GNDA 0.15358f
C2079 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n13 GNDA 0.19139f
C2080 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t45 GNDA 0.15358f
C2081 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n14 GNDA 0.19139f
C2082 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t39 GNDA 0.15358f
C2083 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n15 GNDA 0.19139f
C2084 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t62 GNDA 0.15358f
C2085 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n16 GNDA 0.19139f
C2086 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t29 GNDA 0.15358f
C2087 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n17 GNDA 0.1661f
C2088 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n18 GNDA 0.06574f
C2089 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t9 GNDA 0.31403f
C2090 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t8 GNDA 0.31286f
C2091 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n19 GNDA 0.49793f
C2092 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t15 GNDA 0.31403f
C2093 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t41 GNDA 0.31286f
C2094 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n20 GNDA 0.5037f
C2095 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n21 GNDA 0.53799f
C2096 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t52 GNDA 0.15358f
C2097 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n22 GNDA 0.94496f
C2098 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t34 GNDA 0.15358f
C2099 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n23 GNDA 0.19139f
C2100 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t51 GNDA 0.15358f
C2101 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n24 GNDA 0.19139f
C2102 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t16 GNDA 0.15358f
C2103 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n25 GNDA 0.16326f
C2104 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t60 GNDA 0.15567f
C2105 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t23 GNDA 0.15358f
C2106 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n26 GNDA 0.4875f
C2107 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t61 GNDA 0.15358f
C2108 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n27 GNDA 0.19139f
C2109 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t36 GNDA 0.15358f
C2110 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n28 GNDA 0.19139f
C2111 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t11 GNDA 0.15358f
C2112 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n29 GNDA 0.19139f
C2113 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t35 GNDA 0.15358f
C2114 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n30 GNDA 0.19139f
C2115 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t57 GNDA 0.15358f
C2116 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n31 GNDA 0.19139f
C2117 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t48 GNDA 0.15358f
C2118 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n32 GNDA 0.19139f
C2119 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t13 GNDA 0.15358f
C2120 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n33 GNDA 0.19139f
C2121 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t38 GNDA 0.15358f
C2122 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n34 GNDA 0.1661f
C2123 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n35 GNDA 0.05341f
C2124 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n36 GNDA 0.33285f
C2125 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t63 GNDA 0.15567f
C2126 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t30 GNDA 0.15358f
C2127 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n37 GNDA 0.4875f
C2128 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t28 GNDA 0.15358f
C2129 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n38 GNDA 0.19139f
C2130 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t65 GNDA 0.15358f
C2131 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n39 GNDA 0.16326f
C2132 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t20 GNDA 0.15567f
C2133 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t53 GNDA 0.15358f
C2134 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n40 GNDA 0.4875f
C2135 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t54 GNDA 0.15358f
C2136 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n41 GNDA 0.19139f
C2137 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t18 GNDA 0.15358f
C2138 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n42 GNDA 0.19139f
C2139 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t22 GNDA 0.15358f
C2140 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n43 GNDA 0.19139f
C2141 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t44 GNDA 0.15358f
C2142 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n44 GNDA 0.19139f
C2143 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t17 GNDA 0.15358f
C2144 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n45 GNDA 0.19139f
C2145 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t67 GNDA 0.15358f
C2146 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n46 GNDA 0.19139f
C2147 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t42 GNDA 0.15358f
C2148 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n47 GNDA 0.19139f
C2149 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t64 GNDA 0.15358f
C2150 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n48 GNDA 0.1661f
C2151 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n49 GNDA 0.05341f
C2152 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n50 GNDA 0.23704f
C2153 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t5 GNDA 0.15492f
C2154 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t31 GNDA 0.15358f
C2155 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n51 GNDA 0.38143f
C2156 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t59 GNDA 0.15358f
C2157 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n52 GNDA 0.19139f
C2158 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t10 GNDA 0.15358f
C2159 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n53 GNDA 0.19139f
C2160 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t32 GNDA 0.15358f
C2161 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n54 GNDA 0.16326f
C2162 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t12 GNDA 0.15492f
C2163 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t50 GNDA 0.15358f
C2164 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n55 GNDA 0.38143f
C2165 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t21 GNDA 0.15358f
C2166 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n56 GNDA 0.19139f
C2167 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t7 GNDA 0.15358f
C2168 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n57 GNDA 0.19139f
C2169 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t49 GNDA 0.15358f
C2170 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n58 GNDA 0.19139f
C2171 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t14 GNDA 0.15358f
C2172 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n59 GNDA 0.19139f
C2173 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t56 GNDA 0.15358f
C2174 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n60 GNDA 0.19139f
C2175 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t27 GNDA 0.15358f
C2176 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n61 GNDA 0.19139f
C2177 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t33 GNDA 0.15358f
C2178 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n62 GNDA 0.19139f
C2179 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t55 GNDA 0.15358f
C2180 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n63 GNDA 0.19139f
C2181 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.t37 GNDA 0.15358f
C2182 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n64 GNDA 0.1661f
C2183 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n65 GNDA 0.05341f
C2184 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n66 GNDA 0.5305f
C2185 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n67 GNDA 0.01746f
C2186 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n68 GNDA 0.19226f
C2187 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n69 GNDA 0.0829f
C2188 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n70 GNDA 0.07458f
C2189 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n71 GNDA 0.53524f
C2190 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n72 GNDA 0.07796f
C2191 opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2.n73 GNDA 0.08175f
C2192 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t2 GNDA 0.22296f
C2193 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t16 GNDA 0.22296f
C2194 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n0 GNDA 1.07167f
C2195 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t1 GNDA 0.22296f
C2196 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t6 GNDA 0.22296f
C2197 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n1 GNDA 0.84762f
C2198 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n2 GNDA 1.29878f
C2199 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t3 GNDA 0.22296f
C2200 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t17 GNDA 0.22296f
C2201 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n3 GNDA 1.07167f
C2202 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t15 GNDA 0.22296f
C2203 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t4 GNDA 0.22296f
C2204 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n4 GNDA 0.84762f
C2205 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n5 GNDA 1.36355f
C2206 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t19 GNDA 0.22296f
C2207 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t9 GNDA 0.22296f
C2208 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n6 GNDA 0.84762f
C2209 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n7 GNDA 0.58565f
C2210 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n8 GNDA 0.70528f
C2211 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t5 GNDA 0.22296f
C2212 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t11 GNDA 0.22296f
C2213 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n9 GNDA 1.07167f
C2214 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t8 GNDA 0.22296f
C2215 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t10 GNDA 0.22296f
C2216 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n10 GNDA 0.84762f
C2217 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n11 GNDA 1.36355f
C2218 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t7 GNDA 0.22296f
C2219 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t14 GNDA 0.22296f
C2220 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n12 GNDA 0.84762f
C2221 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n13 GNDA 0.71657f
C2222 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t12 GNDA 0.22296f
C2223 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t0 GNDA 0.22296f
C2224 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n14 GNDA 1.07167f
C2225 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t18 GNDA 0.22296f
C2226 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t13 GNDA 0.22296f
C2227 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n15 GNDA 0.84762f
C2228 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n16 GNDA 1.16787f
C2229 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n17 GNDA 0.52089f
C2230 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n18 GNDA 1.27853f
C2231 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t31 GNDA 0.2513f
C2232 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t35 GNDA 0.24374f
C2233 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n19 GNDA 1.86562f
C2234 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t33 GNDA 0.24374f
C2235 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n20 GNDA 1.07339f
C2236 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t34 GNDA 0.24374f
C2237 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n21 GNDA 1.07339f
C2238 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t32 GNDA 0.24374f
C2239 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n22 GNDA 1.07339f
C2240 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t39 GNDA 0.24374f
C2241 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n23 GNDA 0.85936f
C2242 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t23 GNDA 0.2513f
C2243 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t36 GNDA 0.24374f
C2244 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n24 GNDA 1.86562f
C2245 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t37 GNDA 0.24374f
C2246 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n25 GNDA 1.07339f
C2247 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t21 GNDA 0.24374f
C2248 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n26 GNDA 0.98889f
C2249 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n27 GNDA 0.79614f
C2250 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t22 GNDA 0.2513f
C2251 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t28 GNDA 0.24374f
C2252 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n28 GNDA 1.86562f
C2253 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t25 GNDA 0.24374f
C2254 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n29 GNDA 1.07339f
C2255 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t38 GNDA 0.24374f
C2256 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n30 GNDA 1.07339f
C2257 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t24 GNDA 0.24374f
C2258 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n31 GNDA 0.89746f
C2259 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t30 GNDA 0.2513f
C2260 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t27 GNDA 0.24374f
C2261 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n32 GNDA 1.86562f
C2262 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t20 GNDA 0.24374f
C2263 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n33 GNDA 1.07339f
C2264 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t26 GNDA 0.24374f
C2265 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n34 GNDA 1.07339f
C2266 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.t29 GNDA 0.24374f
C2267 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n35 GNDA 1.02698f
C2268 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n36 GNDA 0.22235f
C2269 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0.n37 GNDA 1.98784f
C2270 VOUT.t45 GNDA 0.01909f
C2271 VOUT.t12 GNDA 0.01909f
C2272 VOUT.n0 GNDA 0.04f
C2273 VOUT.t0 GNDA 0.01909f
C2274 VOUT.t9 GNDA 0.01909f
C2275 VOUT.n1 GNDA 0.04001f
C2276 VOUT.n2 GNDA 0.26526f
C2277 VOUT.n3 GNDA 0.01399f
C2278 VOUT.n4 GNDA 0.01399f
C2279 VOUT.n5 GNDA 0.12211f
C2280 VOUT.t31 GNDA 0.84012f
C2281 VOUT.t38 GNDA 0.79329f
C2282 VOUT.n6 GNDA 0.26836f
C2283 VOUT.t23 GNDA 0.79329f
C2284 VOUT.n7 GNDA 0.13358f
C2285 VOUT.t29 GNDA 0.81388f
C2286 VOUT.n8 GNDA 0.17585f
C2287 VOUT.t24 GNDA 0.84012f
C2288 VOUT.t30 GNDA 0.79329f
C2289 VOUT.n9 GNDA 0.26836f
C2290 VOUT.t36 GNDA 0.79329f
C2291 VOUT.n10 GNDA 0.13358f
C2292 VOUT.t21 GNDA 0.81388f
C2293 VOUT.n11 GNDA 0.16101f
C2294 VOUT.n12 GNDA 0.31526f
C2295 VOUT.t34 GNDA 0.84012f
C2296 VOUT.t40 GNDA 0.79329f
C2297 VOUT.n13 GNDA 0.26836f
C2298 VOUT.t26 GNDA 0.79329f
C2299 VOUT.n14 GNDA 0.13358f
C2300 VOUT.t32 GNDA 0.81388f
C2301 VOUT.n15 GNDA 0.16101f
C2302 VOUT.n16 GNDA 0.21318f
C2303 VOUT.t27 GNDA 0.84012f
C2304 VOUT.t33 GNDA 0.79329f
C2305 VOUT.n17 GNDA 0.26836f
C2306 VOUT.t39 GNDA 0.79329f
C2307 VOUT.n18 GNDA 0.13358f
C2308 VOUT.t25 GNDA 0.81388f
C2309 VOUT.n19 GNDA 0.16101f
C2310 VOUT.n20 GNDA 0.21318f
C2311 VOUT.t37 GNDA 0.84012f
C2312 VOUT.t22 GNDA 0.79329f
C2313 VOUT.n21 GNDA 0.26836f
C2314 VOUT.t28 GNDA 0.79329f
C2315 VOUT.n22 GNDA 0.13358f
C2316 VOUT.t35 GNDA 0.81388f
C2317 VOUT.n23 GNDA 0.16101f
C2318 VOUT.n24 GNDA 0.31977f
C2319 VOUT.t19 GNDA 0.84012f
C2320 VOUT.t13 GNDA 0.79329f
C2321 VOUT.n25 GNDA 0.26836f
C2322 VOUT.t20 GNDA 0.79329f
C2323 VOUT.n26 GNDA 0.13358f
C2324 VOUT.t10 GNDA 0.81388f
C2325 VOUT.n27 GNDA 0.16101f
C2326 VOUT.n28 GNDA 0.31977f
C2327 VOUT.t7 GNDA 0.84012f
C2328 VOUT.t4 GNDA 0.79329f
C2329 VOUT.n29 GNDA 0.26836f
C2330 VOUT.t18 GNDA 0.79329f
C2331 VOUT.n30 GNDA 0.13358f
C2332 VOUT.t5 GNDA 0.81388f
C2333 VOUT.n31 GNDA 0.16101f
C2334 VOUT.n32 GNDA 0.21318f
C2335 VOUT.t46 GNDA 0.84012f
C2336 VOUT.t1 GNDA 0.79329f
C2337 VOUT.n33 GNDA 0.26836f
C2338 VOUT.t43 GNDA 0.79329f
C2339 VOUT.n34 GNDA 0.13358f
C2340 VOUT.t17 GNDA 0.81388f
C2341 VOUT.n35 GNDA 0.16101f
C2342 VOUT.n36 GNDA 0.21318f
C2343 VOUT.t6 GNDA 0.84012f
C2344 VOUT.t11 GNDA 0.79329f
C2345 VOUT.n37 GNDA 0.26836f
C2346 VOUT.t8 GNDA 0.79329f
C2347 VOUT.n38 GNDA 0.13358f
C2348 VOUT.t41 GNDA 0.81388f
C2349 VOUT.n39 GNDA 0.16101f
C2350 VOUT.n40 GNDA 0.21318f
C2351 VOUT.t47 GNDA 0.84012f
C2352 VOUT.t3 GNDA 0.79329f
C2353 VOUT.n41 GNDA 0.26836f
C2354 VOUT.t44 GNDA 0.79329f
C2355 VOUT.n42 GNDA 0.13358f
C2356 VOUT.t14 GNDA 0.81388f
C2357 VOUT.n43 GNDA 0.16101f
C2358 VOUT.n44 GNDA 1.9746f
C2359 VOUT.n45 GNDA 0.66811f
C2360 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t3 GNDA 0.12328f
C2361 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t4 GNDA 0.12328f
C2362 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t24 GNDA 0.03281f
C2363 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t9 GNDA 0.03281f
C2364 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n0 GNDA 0.0687f
C2365 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t26 GNDA 0.12328f
C2366 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t6 GNDA 0.03281f
C2367 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t27 GNDA 0.03281f
C2368 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n1 GNDA 0.0687f
C2369 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t10 GNDA 0.12328f
C2370 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t17 GNDA 0.03281f
C2371 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t22 GNDA 0.03281f
C2372 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n2 GNDA 0.0687f
C2373 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t18 GNDA 0.12328f
C2374 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t37 GNDA 0.81745f
C2375 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t30 GNDA 0.60337f
C2376 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n3 GNDA 0.72202f
C2377 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t39 GNDA 0.81745f
C2378 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t45 GNDA 0.60337f
C2379 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n4 GNDA 0.72202f
C2380 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n5 GNDA 0.14952f
C2381 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t44 GNDA 0.81745f
C2382 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t38 GNDA 0.60337f
C2383 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n6 GNDA 0.72202f
C2384 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t47 GNDA 0.81745f
C2385 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t32 GNDA 0.60337f
C2386 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n7 GNDA 0.72202f
C2387 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n8 GNDA 0.12403f
C2388 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n9 GNDA 0.5418f
C2389 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t34 GNDA 0.81745f
C2390 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t28 GNDA 0.60337f
C2391 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n10 GNDA 0.72202f
C2392 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t36 GNDA 0.81745f
C2393 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t42 GNDA 0.60337f
C2394 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n11 GNDA 0.72202f
C2395 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n12 GNDA 0.12403f
C2396 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n13 GNDA 0.36636f
C2397 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t41 GNDA 0.81745f
C2398 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t35 GNDA 0.60337f
C2399 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n14 GNDA 0.72202f
C2400 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t43 GNDA 0.81745f
C2401 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t29 GNDA 0.60337f
C2402 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n15 GNDA 0.72202f
C2403 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n16 GNDA 0.12403f
C2404 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n17 GNDA 0.36636f
C2405 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t31 GNDA 0.81745f
C2406 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t46 GNDA 0.60337f
C2407 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n18 GNDA 0.72202f
C2408 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t33 GNDA 0.81745f
C2409 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t40 GNDA 0.60337f
C2410 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n19 GNDA 0.72202f
C2411 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n20 GNDA 0.12403f
C2412 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n21 GNDA 3.44672f
C2413 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t16 GNDA 0.07878f
C2414 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t12 GNDA 0.07506f
C2415 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t15 GNDA 0.0175f
C2416 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t7 GNDA 0.0175f
C2417 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n22 GNDA 0.03823f
C2418 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t25 GNDA 0.0175f
C2419 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t20 GNDA 0.0175f
C2420 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n23 GNDA 0.03788f
C2421 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t13 GNDA 0.0175f
C2422 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t19 GNDA 0.0175f
C2423 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n24 GNDA 0.07175f
C2424 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n25 GNDA 0.44438f
C2425 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n26 GNDA 0.39495f
C2426 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n27 GNDA 0.62226f
C2427 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n28 GNDA 0.38487f
C2428 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n29 GNDA 2.15985f
C2429 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n30 GNDA 0.63358f
C2430 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n31 GNDA 0.34778f
C2431 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t21 GNDA 0.12328f
C2432 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n32 GNDA 0.36842f
C2433 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n33 GNDA 0.303f
C2434 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n34 GNDA 0.34778f
C2435 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t14 GNDA 0.12328f
C2436 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n35 GNDA 0.36842f
C2437 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n36 GNDA 0.303f
C2438 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n37 GNDA 0.34778f
C2439 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t11 GNDA 0.12328f
C2440 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n38 GNDA 0.36842f
C2441 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n39 GNDA 0.303f
C2442 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t2 GNDA 0.03281f
C2443 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t0 GNDA 0.03281f
C2444 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n40 GNDA 0.0687f
C2445 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n41 GNDA 0.33884f
C2446 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t1 GNDA 0.12328f
C2447 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n42 GNDA 0.36605f
C2448 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n43 GNDA 0.303f
C2449 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t23 GNDA 0.03281f
C2450 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t8 GNDA 0.03281f
C2451 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n44 GNDA 0.0687f
C2452 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.t5 GNDA 0.12673f
C2453 opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA.n45 GNDA 0.60098f
C2454 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t14 GNDA 0.23722f
C2455 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t16 GNDA 0.23722f
C2456 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n0 GNDA 1.14024f
C2457 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t11 GNDA 0.23722f
C2458 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t10 GNDA 0.23722f
C2459 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n1 GNDA 0.90185f
C2460 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n2 GNDA 1.45079f
C2461 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t6 GNDA 0.23722f
C2462 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t7 GNDA 0.23722f
C2463 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n3 GNDA 0.90185f
C2464 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n4 GNDA 0.80884f
C2465 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t15 GNDA 0.23722f
C2466 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t9 GNDA 0.23722f
C2467 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n5 GNDA 1.14024f
C2468 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t1 GNDA 0.23722f
C2469 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t3 GNDA 0.23722f
C2470 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n6 GNDA 0.90185f
C2471 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n7 GNDA 1.19616f
C2472 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n8 GNDA 0.71788f
C2473 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t17 GNDA 0.23722f
C2474 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t4 GNDA 0.23722f
C2475 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n9 GNDA 1.14024f
C2476 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t19 GNDA 0.23722f
C2477 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t12 GNDA 0.23722f
C2478 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n10 GNDA 0.90185f
C2479 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n11 GNDA 1.42831f
C2480 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t2 GNDA 0.23722f
C2481 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t8 GNDA 0.23722f
C2482 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n12 GNDA 1.14024f
C2483 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t0 GNDA 0.23722f
C2484 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t13 GNDA 0.23722f
C2485 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n13 GNDA 0.90185f
C2486 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n14 GNDA 1.45079f
C2487 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t18 GNDA 0.23722f
C2488 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t5 GNDA 0.23722f
C2489 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n15 GNDA 0.90185f
C2490 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n16 GNDA 0.57669f
C2491 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n17 GNDA 0.55421f
C2492 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n18 GNDA 1.28584f
C2493 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t26 GNDA 0.26404f
C2494 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t33 GNDA 0.25657f
C2495 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n19 GNDA 1.86139f
C2496 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t28 GNDA 0.25657f
C2497 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n20 GNDA 1.07998f
C2498 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t36 GNDA 0.25657f
C2499 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n21 GNDA 1.07998f
C2500 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t27 GNDA 0.25657f
C2501 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n22 GNDA 0.93922f
C2502 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t35 GNDA 0.26404f
C2503 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t31 GNDA 0.25657f
C2504 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n23 GNDA 1.86139f
C2505 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t38 GNDA 0.25657f
C2506 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n24 GNDA 1.07998f
C2507 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t30 GNDA 0.25657f
C2508 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n25 GNDA 1.07998f
C2509 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t34 GNDA 0.25657f
C2510 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n26 GNDA 0.98418f
C2511 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n27 GNDA 0.71895f
C2512 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t37 GNDA 0.26404f
C2513 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t22 GNDA 0.25657f
C2514 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n28 GNDA 1.86139f
C2515 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t20 GNDA 0.25657f
C2516 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n29 GNDA 1.07998f
C2517 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t21 GNDA 0.25657f
C2518 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n30 GNDA 1.07998f
C2519 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t39 GNDA 0.25657f
C2520 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n31 GNDA 1.07998f
C2521 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t25 GNDA 0.25657f
C2522 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n32 GNDA 0.89869f
C2523 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t32 GNDA 0.26404f
C2524 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t23 GNDA 0.25657f
C2525 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n33 GNDA 1.86139f
C2526 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t24 GNDA 0.25657f
C2527 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n34 GNDA 1.07998f
C2528 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.t29 GNDA 0.25657f
C2529 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n35 GNDA 0.94364f
C2530 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n36 GNDA 0.31764f
C2531 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1.n37 GNDA 2.05101f
C2532 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t24 GNDA 2.8674f
C2533 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t2 GNDA 1.93769f
C2534 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n0 GNDA 1.77419f
C2535 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t3 GNDA 0.02043f
C2536 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t1 GNDA 0.09f
C2537 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t7 GNDA 0.06067f
C2538 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t20 GNDA 0.06067f
C2539 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n1 GNDA 0.31327f
C2540 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t22 GNDA 0.06067f
C2541 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t10 GNDA 0.06067f
C2542 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n2 GNDA 0.2523f
C2543 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n3 GNDA 0.37106f
C2544 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t13 GNDA 0.06067f
C2545 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t16 GNDA 0.06067f
C2546 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n4 GNDA 0.2523f
C2547 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n5 GNDA 0.2835f
C2548 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t12 GNDA 0.06067f
C2549 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t11 GNDA 0.06067f
C2550 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n6 GNDA 0.2523f
C2551 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n7 GNDA 0.2835f
C2552 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t8 GNDA 0.06067f
C2553 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t6 GNDA 0.06067f
C2554 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n8 GNDA 0.23066f
C2555 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n9 GNDA 0.38691f
C2556 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t19 GNDA 0.06067f
C2557 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t15 GNDA 0.06067f
C2558 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n10 GNDA 0.29163f
C2559 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t4 GNDA 0.06067f
C2560 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t9 GNDA 0.06067f
C2561 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n11 GNDA 0.2523f
C2562 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n12 GNDA 0.37106f
C2563 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t18 GNDA 0.06067f
C2564 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t14 GNDA 0.06067f
C2565 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n13 GNDA 0.2523f
C2566 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n14 GNDA 0.2835f
C2567 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t21 GNDA 0.06067f
C2568 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t5 GNDA 0.06067f
C2569 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n15 GNDA 0.2523f
C2570 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n16 GNDA 0.2835f
C2571 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t17 GNDA 0.06067f
C2572 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t23 GNDA 0.06067f
C2573 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n17 GNDA 0.2523f
C2574 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n18 GNDA 0.39811f
C2575 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n19 GNDA 4.90173f
C2576 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n20 GNDA 2.44547f
C2577 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n21 GNDA 0.21829f
C2578 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n22 GNDA 0.28717f
C2579 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t0 GNDA 2.8674f
C2580 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.t25 GNDA 1.93769f
C2581 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n23 GNDA 1.76738f
C2582 opa_input_and_self_bias_0/cm_ncell3_0.DRAIN.n24 GNDA 0.20492f
C2583 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t0 GNDA 0.03483f
C2584 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t3 GNDA 0.03483f
C2585 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n0 GNDA 0.07139f
C2586 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n1 GNDA 0.28435f
C2587 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t1 GNDA 0.03483f
C2588 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t2 GNDA 0.03483f
C2589 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n2 GNDA 0.07139f
C2590 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t21 GNDA 0.49404f
C2591 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t11 GNDA 0.49225f
C2592 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n3 GNDA 0.65036f
C2593 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t63 GNDA 0.49225f
C2594 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n4 GNDA 0.32608f
C2595 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t38 GNDA 0.49225f
C2596 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n5 GNDA 0.32608f
C2597 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t13 GNDA 0.49225f
C2598 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n6 GNDA 0.32608f
C2599 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t12 GNDA 0.49225f
C2600 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n7 GNDA 0.32608f
C2601 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t59 GNDA 0.49225f
C2602 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n8 GNDA 0.32608f
C2603 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t17 GNDA 0.49225f
C2604 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n9 GNDA 0.32548f
C2605 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t32 GNDA 0.49404f
C2606 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t54 GNDA 0.49225f
C2607 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n10 GNDA 0.65036f
C2608 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t56 GNDA 0.49225f
C2609 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n11 GNDA 0.32608f
C2610 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t8 GNDA 0.49225f
C2611 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n12 GNDA 0.32608f
C2612 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t9 GNDA 0.49225f
C2613 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n13 GNDA 0.32608f
C2614 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t55 GNDA 0.49225f
C2615 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n14 GNDA 0.32608f
C2616 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t7 GNDA 0.49225f
C2617 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n15 GNDA 0.32608f
C2618 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t61 GNDA 0.49225f
C2619 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n16 GNDA 0.32608f
C2620 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t35 GNDA 0.49225f
C2621 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n17 GNDA 0.32608f
C2622 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t60 GNDA 0.49225f
C2623 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n18 GNDA 0.32608f
C2624 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t5 GNDA 0.49225f
C2625 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n19 GNDA 0.32608f
C2626 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t14 GNDA 0.49225f
C2627 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n20 GNDA 0.25142f
C2628 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n21 GNDA 0.12706f
C2629 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t86 GNDA 0.49404f
C2630 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t73 GNDA 0.49225f
C2631 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n22 GNDA 0.65036f
C2632 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t51 GNDA 0.49225f
C2633 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n23 GNDA 0.32608f
C2634 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t30 GNDA 0.49225f
C2635 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n24 GNDA 0.32608f
C2636 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t76 GNDA 0.49225f
C2637 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n25 GNDA 0.32608f
C2638 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t74 GNDA 0.49225f
C2639 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n26 GNDA 0.32608f
C2640 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t44 GNDA 0.49225f
C2641 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n27 GNDA 0.32608f
C2642 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t81 GNDA 0.49225f
C2643 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n28 GNDA 0.32548f
C2644 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t15 GNDA 0.49404f
C2645 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t39 GNDA 0.49225f
C2646 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n29 GNDA 0.65036f
C2647 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t40 GNDA 0.49225f
C2648 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n30 GNDA 0.32608f
C2649 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t69 GNDA 0.49225f
C2650 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n31 GNDA 0.32608f
C2651 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t71 GNDA 0.49225f
C2652 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n32 GNDA 0.32608f
C2653 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t41 GNDA 0.49225f
C2654 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n33 GNDA 0.32608f
C2655 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t68 GNDA 0.49225f
C2656 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n34 GNDA 0.32608f
C2657 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t50 GNDA 0.49225f
C2658 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n35 GNDA 0.32608f
C2659 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t23 GNDA 0.49225f
C2660 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n36 GNDA 0.32608f
C2661 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t45 GNDA 0.49225f
C2662 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n37 GNDA 0.32608f
C2663 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t67 GNDA 0.49225f
C2664 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n38 GNDA 0.32608f
C2665 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t79 GNDA 0.49225f
C2666 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n39 GNDA 0.25142f
C2667 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n40 GNDA 0.07526f
C2668 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n41 GNDA 0.58913f
C2669 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t33 GNDA 0.49404f
C2670 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t25 GNDA 0.49225f
C2671 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n42 GNDA 0.65036f
C2672 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t82 GNDA 0.49225f
C2673 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n43 GNDA 0.32608f
C2674 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t49 GNDA 0.49225f
C2675 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n44 GNDA 0.32608f
C2676 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t27 GNDA 0.49225f
C2677 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n45 GNDA 0.32608f
C2678 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t26 GNDA 0.49225f
C2679 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n46 GNDA 0.32608f
C2680 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t70 GNDA 0.49225f
C2681 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n47 GNDA 0.32608f
C2682 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t29 GNDA 0.49225f
C2683 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n48 GNDA 0.32548f
C2684 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t37 GNDA 0.49404f
C2685 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t62 GNDA 0.49225f
C2686 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n49 GNDA 0.65036f
C2687 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t64 GNDA 0.49225f
C2688 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n50 GNDA 0.32608f
C2689 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t20 GNDA 0.49225f
C2690 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n51 GNDA 0.32608f
C2691 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t22 GNDA 0.49225f
C2692 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n52 GNDA 0.32608f
C2693 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t65 GNDA 0.49225f
C2694 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n53 GNDA 0.32608f
C2695 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t19 GNDA 0.49225f
C2696 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n54 GNDA 0.32608f
C2697 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t78 GNDA 0.49225f
C2698 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n55 GNDA 0.32608f
C2699 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t43 GNDA 0.49225f
C2700 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n56 GNDA 0.32608f
C2701 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t72 GNDA 0.49225f
C2702 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n57 GNDA 0.32608f
C2703 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t18 GNDA 0.49225f
C2704 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n58 GNDA 0.32608f
C2705 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t28 GNDA 0.49225f
C2706 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n59 GNDA 0.25142f
C2707 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n60 GNDA 0.07526f
C2708 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n61 GNDA 0.37231f
C2709 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t36 GNDA 1.13006f
C2710 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t66 GNDA 1.12853f
C2711 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n62 GNDA 0.96689f
C2712 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t16 GNDA 1.13006f
C2713 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t42 GNDA 1.12853f
C2714 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n63 GNDA 1.14066f
C2715 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n64 GNDA 0.56996f
C2716 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t10 GNDA 0.49225f
C2717 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n65 GNDA 0.6695f
C2718 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t84 GNDA 0.49225f
C2719 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n66 GNDA 0.32608f
C2720 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t58 GNDA 0.49225f
C2721 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n67 GNDA 0.32608f
C2722 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t34 GNDA 0.49225f
C2723 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n68 GNDA 0.32608f
C2724 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t87 GNDA 0.49225f
C2725 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n69 GNDA 0.32608f
C2726 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t85 GNDA 0.49225f
C2727 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n70 GNDA 0.32608f
C2728 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t52 GNDA 0.49225f
C2729 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n71 GNDA 0.32608f
C2730 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t6 GNDA 0.49225f
C2731 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n72 GNDA 0.32548f
C2732 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t24 GNDA 0.49404f
C2733 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t46 GNDA 0.49225f
C2734 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n73 GNDA 0.65036f
C2735 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t47 GNDA 0.49225f
C2736 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n74 GNDA 0.32608f
C2737 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t80 GNDA 0.49225f
C2738 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n75 GNDA 0.32608f
C2739 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t83 GNDA 0.49225f
C2740 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n76 GNDA 0.32608f
C2741 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t48 GNDA 0.49225f
C2742 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n77 GNDA 0.32608f
C2743 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t77 GNDA 0.49225f
C2744 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n78 GNDA 0.32608f
C2745 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t57 GNDA 0.49225f
C2746 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n79 GNDA 0.32608f
C2747 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t31 GNDA 0.49225f
C2748 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n80 GNDA 0.32608f
C2749 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t53 GNDA 0.49225f
C2750 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n81 GNDA 0.32608f
C2751 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t75 GNDA 0.49225f
C2752 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n82 GNDA 0.32608f
C2753 opa_input_and_self_bias_0/cm_pcell3_0.VB2.t4 GNDA 0.49225f
C2754 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n83 GNDA 0.25142f
C2755 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n84 GNDA 0.07526f
C2756 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n85 GNDA 1.44386f
C2757 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n86 GNDA 0.54115f
C2758 opa_input_and_self_bias_0/cm_pcell3_0.VB2.n87 GNDA 0.45905f
C2759 VDDA.n0 GNDA 0.09148f
C2760 VDDA.t255 GNDA 0.04388f
C2761 VDDA.t264 GNDA 0.04388f
C2762 VDDA.n1 GNDA 0.0951f
C2763 VDDA.n2 GNDA 0.03029f
C2764 VDDA.n3 GNDA 0.0995f
C2765 VDDA.n4 GNDA 0.05177f
C2766 VDDA.n5 GNDA 0.63705f
C2767 VDDA.n6 GNDA 0.0461f
C2768 VDDA.t29 GNDA 0.04388f
C2769 VDDA.n7 GNDA 0.14148f
C2770 VDDA.n8 GNDA 0.02759f
C2771 VDDA.n9 GNDA 0.63705f
C2772 VDDA.n10 GNDA 3.45163f
C2773 VDDA.n11 GNDA 0.06008f
C2774 VDDA.n12 GNDA 0.17348f
C2775 VDDA.t254 GNDA 4.15639f
C2776 VDDA.n13 GNDA 0.06008f
C2777 VDDA.n14 GNDA 0.12841f
C2778 VDDA.n15 GNDA 0.12841f
C2779 VDDA.n16 GNDA 0.07313f
C2780 VDDA.n17 GNDA 0.07313f
C2781 VDDA.n18 GNDA 0.17289f
C2782 VDDA.t263 GNDA 0.06841f
C2783 VDDA.t267 GNDA 0.06841f
C2784 VDDA.n19 GNDA 0.2762f
C2785 VDDA.n20 GNDA 0.07725f
C2786 VDDA.n21 GNDA 0.01873f
C2787 VDDA.n22 GNDA 0.05124f
C2788 VDDA.n23 GNDA 0.06346f
C2789 VDDA.n24 GNDA 0.13632f
C2790 VDDA.n25 GNDA 0.14118f
C2791 VDDA.n26 GNDA 0.14274f
C2792 VDDA.n27 GNDA 0.11029f
C2793 VDDA.n28 GNDA 0.06309f
C2794 VDDA.n29 GNDA 0.08088f
C2795 VDDA.n30 GNDA 0.03404f
C2796 VDDA.n31 GNDA 0.08088f
C2797 VDDA.n32 GNDA 0.13632f
C2798 VDDA.n33 GNDA 0.14274f
C2799 VDDA.n34 GNDA 0.07744f
C2800 VDDA.n35 GNDA 0.14118f
C2801 VDDA.n36 GNDA 4.17859f
C2802 VDDA.n37 GNDA 0.11029f
C2803 VDDA.n38 GNDA 0.06309f
C2804 VDDA.n39 GNDA 0.07725f
C2805 VDDA.n40 GNDA 0.03404f
C2806 VDDA.n41 GNDA 0.151f
C2807 VDDA.n42 GNDA 0.09479f
C2808 VDDA.n43 GNDA 0.06244f
C2809 VDDA.n44 GNDA 0.01386f
C2810 VDDA.n45 GNDA 0.41914f
C2811 VDDA.n46 GNDA 0.11897f
C2812 VDDA.t213 GNDA 0.02581f
C2813 VDDA.t202 GNDA 0.02581f
C2814 VDDA.n47 GNDA 0.10025f
C2815 VDDA.n48 GNDA 0.21436f
C2816 VDDA.t203 GNDA 0.02581f
C2817 VDDA.t244 GNDA 0.02581f
C2818 VDDA.n49 GNDA 0.10025f
C2819 VDDA.t221 GNDA 0.02581f
C2820 VDDA.t175 GNDA 0.02581f
C2821 VDDA.n50 GNDA 0.10025f
C2822 VDDA.n51 GNDA 0.21732f
C2823 VDDA.n52 GNDA 0.11762f
C2824 VDDA.n53 GNDA 0.41333f
C2825 VDDA.n55 GNDA 0.01202f
C2826 VDDA.n56 GNDA 0.0642f
C2827 VDDA.n57 GNDA 0.04992f
C2828 VDDA.t61 GNDA 0.02596f
C2829 VDDA.t64 GNDA 0.02601f
C2830 VDDA.t62 GNDA 0.09806f
C2831 VDDA.t65 GNDA 0.02601f
C2832 VDDA.t98 GNDA 0.02581f
C2833 VDDA.t133 GNDA 0.02581f
C2834 VDDA.t92 GNDA 0.02581f
C2835 VDDA.t94 GNDA 0.02581f
C2836 VDDA.n58 GNDA 0.11165f
C2837 VDDA.t132 GNDA 0.02596f
C2838 VDDA.t91 GNDA 0.02596f
C2839 VDDA.t180 GNDA 0.02581f
C2840 VDDA.t193 GNDA 0.02581f
C2841 VDDA.n59 GNDA 0.12108f
C2842 VDDA.t240 GNDA 0.02581f
C2843 VDDA.t172 GNDA 0.02581f
C2844 VDDA.n60 GNDA 0.12108f
C2845 VDDA.n61 GNDA 0.12061f
C2846 VDDA.n62 GNDA 0.1292f
C2847 VDDA.n63 GNDA 0.36793f
C2848 VDDA.n64 GNDA 0.01306f
C2849 VDDA.n65 GNDA 0.22653f
C2850 VDDA.n66 GNDA 0.23956f
C2851 VDDA.n67 GNDA 0.02104f
C2852 VDDA.n68 GNDA 0.24729f
C2853 VDDA.n69 GNDA 0.24855f
C2854 VDDA.n70 GNDA 0.0197f
C2855 VDDA.n71 GNDA 0.01829f
C2856 VDDA.n72 GNDA 0.20849f
C2857 VDDA.n73 GNDA 0.1048f
C2858 VDDA.n74 GNDA 0.06314f
C2859 VDDA.n75 GNDA 0.10684f
C2860 VDDA.n76 GNDA 0.14669f
C2861 VDDA.t11 GNDA 1.05196f
C2862 VDDA.n77 GNDA 0.10809f
C2863 VDDA.n78 GNDA 0.23482f
C2864 VDDA.n79 GNDA 0.41914f
C2865 VDDA.n80 GNDA 0.23405f
C2866 VDDA.n81 GNDA 0.11956f
C2867 VDDA.n82 GNDA 0.01416f
C2868 VDDA.n83 GNDA 0.01386f
C2869 VDDA.n84 GNDA 0.13265f
C2870 VDDA.t169 GNDA 0.02601f
C2871 VDDA.t168 GNDA 0.09806f
C2872 VDDA.t170 GNDA 0.02601f
C2873 VDDA.t154 GNDA 0.02601f
C2874 VDDA.t152 GNDA 0.09806f
C2875 VDDA.t155 GNDA 0.02601f
C2876 VDDA.n85 GNDA 0.14912f
C2877 VDDA.n86 GNDA 0.30962f
C2878 VDDA.n87 GNDA 0.34527f
C2879 VDDA.n88 GNDA 0.23409f
C2880 VDDA.t13 GNDA 1.15015f
C2881 VDDA.n89 GNDA 0.36793f
C2882 VDDA.t265 GNDA 1.31846f
C2883 VDDA.n90 GNDA 0.43674f
C2884 VDDA.n91 GNDA 0.23956f
C2885 VDDA.n92 GNDA 0.13624f
C2886 VDDA.t217 GNDA 0.02581f
C2887 VDDA.t219 GNDA 0.02581f
C2888 VDDA.n93 GNDA 0.10464f
C2889 VDDA.n94 GNDA 0.10838f
C2890 VDDA.t231 GNDA 0.02581f
C2891 VDDA.t249 GNDA 0.02581f
C2892 VDDA.n95 GNDA 0.10464f
C2893 VDDA.t199 GNDA 0.02581f
C2894 VDDA.t239 GNDA 0.02581f
C2895 VDDA.n96 GNDA 0.10464f
C2896 VDDA.t230 GNDA 0.02581f
C2897 VDDA.t173 GNDA 0.02581f
C2898 VDDA.n97 GNDA 0.10464f
C2899 VDDA.t225 GNDA 0.02581f
C2900 VDDA.t229 GNDA 0.02581f
C2901 VDDA.n98 GNDA 0.10464f
C2902 VDDA.t174 GNDA 0.02581f
C2903 VDDA.t176 GNDA 0.02581f
C2904 VDDA.n99 GNDA 0.10464f
C2905 VDDA.t204 GNDA 0.02581f
C2906 VDDA.t45 GNDA 0.02581f
C2907 VDDA.n100 GNDA 0.10058f
C2908 VDDA.t46 GNDA 0.02581f
C2909 VDDA.t49 GNDA 0.02581f
C2910 VDDA.n101 GNDA 0.12009f
C2911 VDDA.t111 GNDA 0.02608f
C2912 VDDA.t109 GNDA 0.09806f
C2913 VDDA.n102 GNDA 0.0795f
C2914 VDDA.t107 GNDA 0.02608f
C2915 VDDA.t106 GNDA 0.09806f
C2916 VDDA.n103 GNDA 0.0795f
C2917 VDDA.t108 GNDA 0.02581f
C2918 VDDA.t110 GNDA 0.02581f
C2919 VDDA.n104 GNDA 0.09466f
C2920 VDDA.n105 GNDA 0.06659f
C2921 VDDA.t50 GNDA 0.02596f
C2922 VDDA.n106 GNDA 0.08404f
C2923 VDDA.n107 GNDA 0.13153f
C2924 VDDA.t16 GNDA 0.07161f
C2925 VDDA.n108 GNDA 0.20069f
C2926 VDDA.n109 GNDA 0.07269f
C2927 VDDA.n110 GNDA 0.12999f
C2928 VDDA.n111 GNDA 0.92691f
C2929 VDDA.n112 GNDA 0.92691f
C2930 VDDA.t258 GNDA 0.77166f
C2931 VDDA.t15 GNDA 0.77166f
C2932 VDDA.n113 GNDA 0.43907f
C2933 VDDA.n114 GNDA 0.12999f
C2934 VDDA.n115 GNDA 0.0734f
C2935 VDDA.t262 GNDA 0.07161f
C2936 VDDA.n116 GNDA 0.20069f
C2937 VDDA.n117 GNDA 0.10069f
C2938 VDDA.n118 GNDA 0.15553f
C2939 VDDA.n119 GNDA 0.07269f
C2940 VDDA.n120 GNDA 0.0734f
C2941 VDDA.n121 GNDA 0.03663f
C2942 VDDA.n122 GNDA 0.70391f
C2943 VDDA.n123 GNDA 0.72582f
C2944 VDDA.n124 GNDA 0.01884f
C2945 VDDA.n125 GNDA 0.06314f
C2946 VDDA.n126 GNDA 0.10872f
C2947 VDDA.n127 GNDA 0.14669f
C2948 VDDA.n128 GNDA 0.10684f
C2949 VDDA.n129 GNDA 0.23486f
C2950 VDDA.n130 GNDA 0.23738f
C2951 VDDA.t163 GNDA 0.02597f
C2952 VDDA.t164 GNDA 0.02597f
C2953 VDDA.t144 GNDA 0.02597f
C2954 VDDA.t145 GNDA 0.02597f
C2955 VDDA.t147 GNDA 0.02601f
C2956 VDDA.t146 GNDA 0.09806f
C2957 VDDA.t148 GNDA 0.02601f
C2958 VDDA.t101 GNDA 0.02601f
C2959 VDDA.t99 GNDA 0.09806f
C2960 VDDA.t102 GNDA 0.02601f
C2961 VDDA.n131 GNDA 0.30958f
C2962 VDDA.n132 GNDA 0.14912f
C2963 VDDA.n133 GNDA 0.06244f
C2964 VDDA.n134 GNDA 0.05824f
C2965 VDDA.n135 GNDA 0.08993f
C2966 VDDA.t143 GNDA 0.09806f
C2967 VDDA.n136 GNDA 0.03789f
C2968 VDDA.n137 GNDA 0.2247f
C2969 VDDA.n138 GNDA 0.34025f
C2970 VDDA.n139 GNDA 0.22478f
C2971 VDDA.t162 GNDA 0.09806f
C2972 VDDA.n140 GNDA 0.03789f
C2973 VDDA.n141 GNDA 0.06878f
C2974 VDDA.n142 GNDA 0.08302f
C2975 VDDA.n143 GNDA 0.03662f
C2976 VDDA.n144 GNDA 0.11959f
C2977 VDDA.n145 GNDA 0.01386f
C2978 VDDA.n146 GNDA 0.23486f
C2979 VDDA.n147 GNDA -0.53185f
C2980 VDDA.n148 GNDA 0.05443f
C2981 VDDA.n149 GNDA 0.06518f
C2982 VDDA.t166 GNDA 0.02596f
C2983 VDDA.t80 GNDA 0.02581f
C2984 VDDA.t211 GNDA 0.02581f
C2985 VDDA.n150 GNDA 0.10058f
C2986 VDDA.t224 GNDA 0.02581f
C2987 VDDA.t241 GNDA 0.02581f
C2988 VDDA.n151 GNDA 0.10464f
C2989 VDDA.t195 GNDA 0.02581f
C2990 VDDA.t220 GNDA 0.02581f
C2991 VDDA.n152 GNDA 0.10464f
C2992 VDDA.t223 GNDA 0.02581f
C2993 VDDA.t250 GNDA 0.02581f
C2994 VDDA.n153 GNDA 0.10464f
C2995 VDDA.n154 GNDA 0.10838f
C2996 VDDA.n155 GNDA 0.10838f
C2997 VDDA.n156 GNDA 0.1097f
C2998 VDDA.n157 GNDA 0.09058f
C2999 VDDA.t78 GNDA 0.09806f
C3000 VDDA.n158 GNDA 0.04809f
C3001 VDDA.t123 GNDA 0.02601f
C3002 VDDA.t121 GNDA 0.09806f
C3003 VDDA.t124 GNDA 0.02601f
C3004 VDDA.t116 GNDA 0.02596f
C3005 VDDA.n159 GNDA 0.08145f
C3006 VDDA.n160 GNDA 0.15917f
C3007 VDDA.t115 GNDA 0.09806f
C3008 VDDA.n161 GNDA 0.05955f
C3009 VDDA.t58 GNDA 0.02581f
C3010 VDDA.t226 GNDA 0.02581f
C3011 VDDA.n162 GNDA 0.09214f
C3012 VDDA.t228 GNDA 0.02581f
C3013 VDDA.t188 GNDA 0.02581f
C3014 VDDA.n163 GNDA 0.10025f
C3015 VDDA.t238 GNDA 0.02581f
C3016 VDDA.t214 GNDA 0.02581f
C3017 VDDA.n164 GNDA 0.10025f
C3018 VDDA.t207 GNDA 0.02581f
C3019 VDDA.t181 GNDA 0.02581f
C3020 VDDA.n165 GNDA 0.10025f
C3021 VDDA.n166 GNDA 0.21732f
C3022 VDDA.n167 GNDA 0.21732f
C3023 VDDA.n168 GNDA 0.21498f
C3024 VDDA.n169 GNDA 0.15958f
C3025 VDDA.t55 GNDA 0.09806f
C3026 VDDA.n170 GNDA 0.0911f
C3027 VDDA.n171 GNDA 0.08907f
C3028 VDDA.t117 GNDA 0.02581f
C3029 VDDA.t57 GNDA 0.02581f
C3030 VDDA.n172 GNDA 0.11165f
C3031 VDDA.t120 GNDA 0.02581f
C3032 VDDA.t160 GNDA 0.02581f
C3033 VDDA.n173 GNDA 0.11165f
C3034 VDDA.t119 GNDA 0.02596f
C3035 VDDA.t76 GNDA 0.02596f
C3036 VDDA.n174 GNDA 0.11347f
C3037 VDDA.t75 GNDA 0.09806f
C3038 VDDA.t118 GNDA 0.09806f
C3039 VDDA.n175 GNDA 0.10084f
C3040 VDDA.t140 GNDA 0.09806f
C3041 VDDA.t161 GNDA 0.02596f
C3042 VDDA.t142 GNDA 0.02596f
C3043 VDDA.t177 GNDA 0.02581f
C3044 VDDA.t185 GNDA 0.02581f
C3045 VDDA.n176 GNDA 0.12108f
C3046 VDDA.t234 GNDA 0.02581f
C3047 VDDA.t246 GNDA 0.02581f
C3048 VDDA.n177 GNDA 0.12108f
C3049 VDDA.t206 GNDA 0.02581f
C3050 VDDA.t233 GNDA 0.02581f
C3051 VDDA.n178 GNDA 0.12108f
C3052 VDDA.t187 GNDA 0.02581f
C3053 VDDA.t212 GNDA 0.02581f
C3054 VDDA.n179 GNDA 0.12108f
C3055 VDDA.t182 GNDA 0.02581f
C3056 VDDA.t183 GNDA 0.02581f
C3057 VDDA.n180 GNDA 0.12108f
C3058 VDDA.t242 GNDA 0.02581f
C3059 VDDA.t245 GNDA 0.02581f
C3060 VDDA.n181 GNDA 0.12108f
C3061 VDDA.t210 GNDA 0.02581f
C3062 VDDA.t178 GNDA 0.02581f
C3063 VDDA.n182 GNDA 0.12108f
C3064 VDDA.t197 GNDA 0.02581f
C3065 VDDA.t237 GNDA 0.02581f
C3066 VDDA.n183 GNDA 0.12108f
C3067 VDDA.n184 GNDA 0.13633f
C3068 VDDA.n185 GNDA 0.13633f
C3069 VDDA.n186 GNDA 0.13633f
C3070 VDDA.n187 GNDA 0.12304f
C3071 VDDA.n188 GNDA 0.12532f
C3072 VDDA.t159 GNDA 0.09806f
C3073 VDDA.n189 GNDA 0.10084f
C3074 VDDA.n190 GNDA 0.10575f
C3075 VDDA.t77 GNDA 0.02581f
C3076 VDDA.t141 GNDA 0.02581f
C3077 VDDA.n191 GNDA 0.11165f
C3078 VDDA.t167 GNDA 0.02581f
C3079 VDDA.t79 GNDA 0.02581f
C3080 VDDA.n192 GNDA 0.12009f
C3081 VDDA.t151 GNDA 0.02608f
C3082 VDDA.t149 GNDA 0.09806f
C3083 VDDA.n193 GNDA 0.0795f
C3084 VDDA.t85 GNDA 0.02608f
C3085 VDDA.t84 GNDA 0.09806f
C3086 VDDA.n194 GNDA 0.0795f
C3087 VDDA.t86 GNDA 0.02581f
C3088 VDDA.t150 GNDA 0.02581f
C3089 VDDA.n195 GNDA 0.09466f
C3090 VDDA.n196 GNDA 0.06659f
C3091 VDDA.n197 GNDA 0.08781f
C3092 VDDA.t165 GNDA 0.09806f
C3093 VDDA.n198 GNDA 0.05045f
C3094 VDDA.n199 GNDA 0.0639f
C3095 VDDA.n200 GNDA 0.08015f
C3096 VDDA.n201 GNDA 0.05443f
C3097 VDDA.n202 GNDA 0.01268f
C3098 VDDA.n203 GNDA 0.01239f
C3099 VDDA.n204 GNDA 0.04125f
C3100 VDDA.n205 GNDA 0.24729f
C3101 VDDA.n206 GNDA 0.24855f
C3102 VDDA.n207 GNDA 0.01914f
C3103 VDDA.n208 GNDA 0.14211f
C3104 VDDA.n209 GNDA 0.01884f
C3105 VDDA.n210 GNDA 0.06327f
C3106 VDDA.n211 GNDA 0.22653f
C3107 VDDA.n212 GNDA 0.01239f
C3108 VDDA.n213 GNDA 0.22596f
C3109 VDDA.n214 GNDA 1.71059f
C3110 VDDA.t153 GNDA 1.45654f
C3111 VDDA.t122 GNDA 0.03387f
C3112 VDDA.t52 GNDA 1.51971f
C3113 VDDA.n215 GNDA 2.56306f
C3114 VDDA.t56 GNDA 3.34525f
C3115 VDDA.t260 GNDA 2.63692f
C3116 VDDA.t23 GNDA 1.80938f
C3117 VDDA.t256 GNDA 2.63692f
C3118 VDDA.t32 GNDA 0.90469f
C3119 VDDA.n216 GNDA 0.10809f
C3120 VDDA.t38 GNDA 1.90756f
C3121 VDDA.n217 GNDA 0.10684f
C3122 VDDA.n218 GNDA 0.06124f
C3123 VDDA.n219 GNDA 0.06084f
C3124 VDDA.n220 GNDA 0.10684f
C3125 VDDA.t26 GNDA 0.1052f
C3126 VDDA.t253 GNDA 1.43768f
C3127 VDDA.t30 GNDA 2.53173f
C3128 VDDA.t33 GNDA 1.80938f
C3129 VDDA.t14 GNDA 1.61301f
C3130 VDDA.t37 GNDA 1.02391f
C3131 VDDA.n221 GNDA 0.10684f
C3132 VDDA.t21 GNDA 1.80938f
C3133 VDDA.t36 GNDA 2.63692f
C3134 VDDA.t25 GNDA 3.34525f
C3135 VDDA.t171 GNDA 3.1068f
C3136 VDDA.t179 GNDA 2.87537f
C3137 VDDA.n222 GNDA 2.63692f
C3138 VDDA.n223 GNDA 0.07508f
C3139 VDDA.n224 GNDA 0.04313f
C3140 VDDA.t136 GNDA 0.02608f
C3141 VDDA.t134 GNDA 0.09806f
C3142 VDDA.n225 GNDA 0.0795f
C3143 VDDA.t73 GNDA 0.02608f
C3144 VDDA.t72 GNDA 0.09806f
C3145 VDDA.n226 GNDA 0.0795f
C3146 VDDA.t74 GNDA 0.02581f
C3147 VDDA.t135 GNDA 0.02581f
C3148 VDDA.n227 GNDA 0.09466f
C3149 VDDA.n228 GNDA 0.06254f
C3150 VDDA.n229 GNDA 0.27366f
C3151 VDDA.t89 GNDA 0.02608f
C3152 VDDA.t87 GNDA 0.09806f
C3153 VDDA.n230 GNDA 0.0795f
C3154 VDDA.t82 GNDA 0.02608f
C3155 VDDA.t81 GNDA 0.09806f
C3156 VDDA.n231 GNDA 0.0795f
C3157 VDDA.t83 GNDA 0.02581f
C3158 VDDA.t88 GNDA 0.02581f
C3159 VDDA.n232 GNDA 0.09466f
C3160 VDDA.n233 GNDA 0.06254f
C3161 VDDA.n234 GNDA 0.32012f
C3162 VDDA.n235 GNDA 0.43357f
C3163 VDDA.n236 GNDA 0.10872f
C3164 VDDA.n237 GNDA 0.10684f
C3165 VDDA.t22 GNDA 0.90469f
C3166 VDDA.n238 GNDA 0.0693f
C3167 VDDA.t7 GNDA 3.34525f
C3168 VDDA.n239 GNDA 0.10684f
C3169 VDDA.n240 GNDA 0.03927f
C3170 VDDA.n241 GNDA 0.06124f
C3171 VDDA.n242 GNDA 0.06084f
C3172 VDDA.n243 GNDA 0.10684f
C3173 VDDA.t6 GNDA 2.63692f
C3174 VDDA.t41 GNDA 1.80938f
C3175 VDDA.t4 GNDA 2.11796f
C3176 VDDA.t35 GNDA 0.07714f
C3177 VDDA.t257 GNDA 0.44884f
C3178 VDDA.t9 GNDA 0.82754f
C3179 VDDA.t2 GNDA 2.1951f
C3180 VDDA.t3 GNDA 2.2512f
C3181 VDDA.t8 GNDA 3.07875f
C3182 VDDA.t20 GNDA 2.90342f
C3183 VDDA.t42 GNDA 1.80938f
C3184 VDDA.t5 GNDA 2.63692f
C3185 VDDA.t40 GNDA 3.34525f
C3186 VDDA.n244 GNDA 2.63692f
C3187 VDDA.n245 GNDA 0.07508f
C3188 VDDA.n246 GNDA 0.04313f
C3189 VDDA.n247 GNDA 0.10872f
C3190 VDDA.n248 GNDA 0.16926f
C3191 VDDA.n249 GNDA 0.0693f
C3192 VDDA.n250 GNDA 0.97482f
C3193 VDDA.n251 GNDA 0.0693f
C3194 VDDA.n252 GNDA 0.03927f
C3195 VDDA.n253 GNDA 0.06084f
C3196 VDDA.n254 GNDA 0.04313f
C3197 VDDA.n255 GNDA 0.07508f
C3198 VDDA.n256 GNDA 2.63692f
C3199 VDDA.t39 GNDA 3.34525f
C3200 VDDA.t31 GNDA 2.63692f
C3201 VDDA.t34 GNDA 1.80938f
C3202 VDDA.t27 GNDA 2.0899f
C3203 VDDA.n257 GNDA 1.45171f
C3204 VDDA.n258 GNDA 0.0693f
C3205 VDDA.n259 GNDA 0.11179f
C3206 VDDA.n260 GNDA 0.08379f
C3207 VDDA.n261 GNDA 0.10872f
C3208 VDDA.n262 GNDA 0.16926f
C3209 VDDA.n263 GNDA 0.0693f
C3210 VDDA.n264 GNDA 1.80938f
C3211 VDDA.n265 GNDA 0.0693f
C3212 VDDA.n266 GNDA 0.03927f
C3213 VDDA.n267 GNDA 0.06084f
C3214 VDDA.n268 GNDA 0.04313f
C3215 VDDA.n269 GNDA 0.07508f
C3216 VDDA.n270 GNDA 2.63692f
C3217 VDDA.t24 GNDA 3.34525f
C3218 VDDA.t18 GNDA 2.63692f
C3219 VDDA.t19 GNDA 1.80938f
C3220 VDDA.t261 GNDA 2.59485f
C3221 VDDA.n271 GNDA 0.94677f
C3222 VDDA.n272 GNDA 0.10809f
C3223 VDDA.n273 GNDA 0.17095f
C3224 VDDA.n274 GNDA 0.14135f
C3225 VDDA.n275 GNDA 0.03125f
C3226 VDDA.n276 GNDA 0.07967f
C3227 VDDA.n277 GNDA 0.10795f
C3228 VDDA.t114 GNDA 0.02608f
C3229 VDDA.t112 GNDA 0.09806f
C3230 VDDA.n278 GNDA 0.0795f
C3231 VDDA.t53 GNDA 0.02608f
C3232 VDDA.t51 GNDA 0.09806f
C3233 VDDA.n279 GNDA 0.0795f
C3234 VDDA.t54 GNDA 0.02581f
C3235 VDDA.t113 GNDA 0.02581f
C3236 VDDA.n280 GNDA 0.09466f
C3237 VDDA.n281 GNDA 0.06254f
C3238 VDDA.t158 GNDA 0.02608f
C3239 VDDA.t156 GNDA 0.09806f
C3240 VDDA.n282 GNDA 0.0795f
C3241 VDDA.t104 GNDA 0.02608f
C3242 VDDA.t103 GNDA 0.09806f
C3243 VDDA.n283 GNDA 0.0795f
C3244 VDDA.t105 GNDA 0.02581f
C3245 VDDA.t157 GNDA 0.02581f
C3246 VDDA.n284 GNDA 0.09466f
C3247 VDDA.n285 GNDA 0.06254f
C3248 VDDA.n286 GNDA 0.29505f
C3249 VDDA.n287 GNDA 0.43357f
C3250 VDDA.t71 GNDA 0.02608f
C3251 VDDA.t69 GNDA 0.09806f
C3252 VDDA.n288 GNDA 0.0795f
C3253 VDDA.t67 GNDA 0.02608f
C3254 VDDA.t66 GNDA 0.09806f
C3255 VDDA.n289 GNDA 0.0795f
C3256 VDDA.t68 GNDA 0.02581f
C3257 VDDA.t70 GNDA 0.02581f
C3258 VDDA.n290 GNDA 0.09466f
C3259 VDDA.n291 GNDA 0.06254f
C3260 VDDA.t130 GNDA 0.02608f
C3261 VDDA.t128 GNDA 0.09806f
C3262 VDDA.n292 GNDA 0.0795f
C3263 VDDA.t126 GNDA 0.02608f
C3264 VDDA.t125 GNDA 0.09806f
C3265 VDDA.n293 GNDA 0.0795f
C3266 VDDA.t127 GNDA 0.02581f
C3267 VDDA.t129 GNDA 0.02581f
C3268 VDDA.n294 GNDA 0.09466f
C3269 VDDA.n295 GNDA 0.06254f
C3270 VDDA.n296 GNDA 0.295f
C3271 VDDA.n297 GNDA 0.10719f
C3272 VDDA.n298 GNDA 0.08485f
C3273 VDDA.n299 GNDA 0.05525f
C3274 VDDA.n300 GNDA 0.07907f
C3275 VDDA.n301 GNDA 0.06417f
C3276 VDDA.t47 GNDA 0.09806f
C3277 VDDA.n302 GNDA 0.05045f
C3278 VDDA.n303 GNDA 0.08781f
C3279 VDDA.t43 GNDA 0.09806f
C3280 VDDA.n304 GNDA 0.04809f
C3281 VDDA.n305 GNDA 0.09058f
C3282 VDDA.n306 GNDA 0.1097f
C3283 VDDA.n307 GNDA 0.10838f
C3284 VDDA.n308 GNDA 0.10838f
C3285 VDDA.n309 GNDA 0.10838f
C3286 VDDA.n310 GNDA 0.10838f
C3287 VDDA.n311 GNDA 0.13622f
C3288 VDDA.n312 GNDA 0.20849f
C3289 VDDA.n313 GNDA 0.36793f
C3290 VDDA.n314 GNDA 1.12911f
C3291 VDDA.n315 GNDA 0.84859f
C3292 VDDA.n316 GNDA 0.36965f
C3293 VDDA.n317 GNDA 0.20947f
C3294 VDDA.n318 GNDA 0.13263f
C3295 VDDA.n319 GNDA 0.01386f
C3296 VDDA.n320 GNDA 0.23482f
C3297 VDDA.n321 GNDA 1.83743f
C3298 VDDA.t48 GNDA 2.12497f
C3299 VDDA.t63 GNDA 0.30858f
C3300 VDDA.t100 GNDA 1.20625f
C3301 VDDA.t10 GNDA 2.32835f
C3302 VDDA.t44 GNDA 1.80938f
C3303 VDDA.t17 GNDA 1.58496f
C3304 VDDA.n322 GNDA 1.80938f
C3305 VDDA.n323 GNDA 0.10809f
C3306 VDDA.n324 GNDA 0.16926f
C3307 VDDA.n325 GNDA 0.1135f
C3308 VDDA.n326 GNDA 0.01361f
C3309 VDDA.n327 GNDA 0.0197f
C3310 VDDA.n329 GNDA 0.14061f
C3311 VDDA.n330 GNDA 0.01829f
C3312 VDDA.n331 GNDA 0.06327f
C3313 VDDA.n332 GNDA 0.22596f
C3314 VDDA.n333 GNDA 1.29041f
C3315 VDDA.n334 GNDA 0.04125f
C3316 VDDA.n335 GNDA 0.01202f
C3317 VDDA.n336 GNDA 0.12808f
C3318 VDDA.n337 GNDA 0.20849f
C3319 VDDA.n338 GNDA 0.03144f
C3320 VDDA.t209 GNDA 0.02581f
C3321 VDDA.t236 GNDA 0.02581f
C3322 VDDA.n339 GNDA 0.12108f
C3323 VDDA.t196 GNDA 0.02581f
C3324 VDDA.t222 GNDA 0.02581f
C3325 VDDA.n340 GNDA 0.12108f
C3326 VDDA.n341 GNDA 0.12061f
C3327 VDDA.t208 GNDA 0.02581f
C3328 VDDA.t190 GNDA 0.02581f
C3329 VDDA.n342 GNDA 0.12108f
C3330 VDDA.t191 GNDA 0.02581f
C3331 VDDA.t252 GNDA 0.02581f
C3332 VDDA.n343 GNDA 0.12108f
C3333 VDDA.n344 GNDA 0.13633f
C3334 VDDA.t215 GNDA 0.02581f
C3335 VDDA.t186 GNDA 0.02581f
C3336 VDDA.n345 GNDA 0.12108f
C3337 VDDA.t200 GNDA 0.02581f
C3338 VDDA.t248 GNDA 0.02581f
C3339 VDDA.n346 GNDA 0.12108f
C3340 VDDA.n347 GNDA 0.13633f
C3341 VDDA.t189 GNDA 0.02581f
C3342 VDDA.t216 GNDA 0.02581f
C3343 VDDA.n348 GNDA 0.12108f
C3344 VDDA.t251 GNDA 0.02581f
C3345 VDDA.t201 GNDA 0.02581f
C3346 VDDA.n349 GNDA 0.12108f
C3347 VDDA.n350 GNDA 0.13633f
C3348 VDDA.t218 GNDA 0.02581f
C3349 VDDA.t247 GNDA 0.02581f
C3350 VDDA.n351 GNDA 0.12108f
C3351 VDDA.t194 GNDA 0.02581f
C3352 VDDA.t232 GNDA 0.02581f
C3353 VDDA.n352 GNDA 0.12108f
C3354 VDDA.n353 GNDA 0.12304f
C3355 VDDA.n354 GNDA 0.12532f
C3356 VDDA.t90 GNDA 0.09806f
C3357 VDDA.t131 GNDA 0.09806f
C3358 VDDA.n355 GNDA 0.10084f
C3359 VDDA.t93 GNDA 0.09806f
C3360 VDDA.t139 GNDA 0.02596f
C3361 VDDA.t95 GNDA 0.02596f
C3362 VDDA.n356 GNDA 0.11364f
C3363 VDDA.t137 GNDA 0.09806f
C3364 VDDA.n357 GNDA 0.10084f
C3365 VDDA.n358 GNDA 0.10575f
C3366 VDDA.t138 GNDA 0.02581f
C3367 VDDA.n359 GNDA 0.11165f
C3368 VDDA.t60 GNDA 0.02581f
C3369 VDDA.n360 GNDA 0.11165f
C3370 VDDA.t243 GNDA 0.02581f
C3371 VDDA.t97 GNDA 0.02581f
C3372 VDDA.n361 GNDA 0.09214f
C3373 VDDA.t205 GNDA 0.02581f
C3374 VDDA.t192 GNDA 0.02581f
C3375 VDDA.n362 GNDA 0.10025f
C3376 VDDA.t198 GNDA 0.02581f
C3377 VDDA.t227 GNDA 0.02581f
C3378 VDDA.n363 GNDA 0.10025f
C3379 VDDA.t184 GNDA 0.02581f
C3380 VDDA.t235 GNDA 0.02581f
C3381 VDDA.n364 GNDA 0.10025f
C3382 VDDA.n365 GNDA 0.21732f
C3383 VDDA.n366 GNDA 0.21732f
C3384 VDDA.n367 GNDA 0.21498f
C3385 VDDA.n368 GNDA 0.15958f
C3386 VDDA.t96 GNDA 0.09806f
C3387 VDDA.n369 GNDA 0.0911f
C3388 VDDA.n370 GNDA 0.08165f
C3389 VDDA.n371 GNDA 0.16935f
C3390 VDDA.t59 GNDA 0.09806f
C3391 VDDA.n372 GNDA 0.05592f
C3392 VDDA.n373 GNDA 0.06697f
C3393 VDDA.n374 GNDA 0.08598f
C3394 VDDA.n375 GNDA 0.0581f
C3395 VDDA.n376 GNDA 0.11797f
C3396 VDDA.n377 GNDA 0.23344f
C3397 VDDA.n378 GNDA 0.12778f
C3398 VDDA.n379 GNDA 0.09249f
C3399 VDDA.n380 GNDA 0.22342f
C3400 VDDA.n381 GNDA 0.11959f
C3401 VDDA.n382 GNDA 0.07141f
C3402 VDDA.n383 GNDA 0.10249f
C3403 VDDA.n384 GNDA 0.16527f
C3404 VDDA.n385 GNDA 0.13087f
C3405 VDDA.t1 GNDA 0.04388f
C3406 VDDA.n386 GNDA 0.14148f
C3407 VDDA.n387 GNDA 0.12923f
C3408 VDDA.n388 GNDA 0.64008f
C3409 VDDA.n389 GNDA 0.69827f
C3410 VDDA.n390 GNDA 0.40891f
C3411 VDDA.n391 GNDA 0.07971f
C3412 VDDA.t266 GNDA 0.06841f
C3413 VDDA.t259 GNDA 0.06841f
C3414 VDDA.n392 GNDA 0.2762f
C3415 VDDA.n393 GNDA 0.07202f
C3416 VDDA.n394 GNDA 0.09082f
C3417 VDDA.n395 GNDA 0.16051f
C3418 VDDA.n396 GNDA 2.08652f
C3419 VDDA.t12 GNDA 1.77021f
C3420 VDDA.t0 GNDA 0.52102f
C3421 VDDA.t28 GNDA 0.52102f
C3422 VDDA.n397 GNDA 3.4094f
C3423 VDDA.n398 GNDA 0.0995f
C3424 VDDA.n399 GNDA 0.05622f
C3425 VDDA.n400 GNDA 0.0461f
C3426 VDDA.n401 GNDA 0.03029f
C3427 VDDA.n402 GNDA 0.01873f
C3428 VDDA.n403 GNDA 0.02759f
C3429 VDDA.n404 GNDA 0.09724f
C3430 VDDA.n405 GNDA 0.05155f
C3431 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t7 GNDA 0.18931f
C3432 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t2 GNDA 0.18931f
C3433 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n0 GNDA 0.73533f
C3434 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t5 GNDA 0.18936f
C3435 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t4 GNDA 0.18936f
C3436 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n1 GNDA 0.95127f
C3437 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n2 GNDA 1.158f
C3438 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t6 GNDA 0.18936f
C3439 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t1 GNDA 0.18936f
C3440 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n3 GNDA 0.86568f
C3441 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t3 GNDA 0.18931f
C3442 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t8 GNDA 0.18931f
C3443 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n4 GNDA 0.85788f
C3444 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n5 GNDA 1.09031f
C3445 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n6 GNDA 0.69922f
C3446 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t13 GNDA 0.21344f
C3447 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t15 GNDA 0.20701f
C3448 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n7 GNDA 1.36507f
C3449 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t10 GNDA 0.21344f
C3450 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t9 GNDA 0.20701f
C3451 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n8 GNDA 1.77158f
C3452 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n9 GNDA 0.47809f
C3453 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t11 GNDA 0.21344f
C3454 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t12 GNDA 0.20701f
C3455 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n10 GNDA 1.58627f
C3456 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t14 GNDA 0.21344f
C3457 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.t0 GNDA 0.20701f
C3458 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n11 GNDA 1.55038f
C3459 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n12 GNDA 0.47475f
C3460 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3.n13 GNDA 0.65091f
C3461 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t48 GNDA 0.5333f
C3462 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t46 GNDA 0.53137f
C3463 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n0 GNDA 0.70204f
C3464 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t86 GNDA 0.53137f
C3465 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n1 GNDA 0.35199f
C3466 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t36 GNDA 0.53137f
C3467 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n2 GNDA 0.35199f
C3468 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t60 GNDA 0.53137f
C3469 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n3 GNDA 0.35199f
C3470 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t67 GNDA 0.53137f
C3471 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n4 GNDA 0.35199f
C3472 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t93 GNDA 0.53137f
C3473 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n5 GNDA 0.35199f
C3474 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t61 GNDA 0.53137f
C3475 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n6 GNDA 0.35199f
C3476 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t72 GNDA 0.53137f
C3477 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n7 GNDA 0.35199f
C3478 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t71 GNDA 0.53137f
C3479 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n8 GNDA 0.35199f
C3480 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t30 GNDA 0.53137f
C3481 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n9 GNDA 0.35199f
C3482 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t53 GNDA 0.53137f
C3483 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n10 GNDA 0.2714f
C3484 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t32 GNDA 0.5333f
C3485 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t82 GNDA 0.53137f
C3486 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n11 GNDA 0.70204f
C3487 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t69 GNDA 0.53137f
C3488 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n12 GNDA 0.35199f
C3489 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t47 GNDA 0.53137f
C3490 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n13 GNDA 0.35199f
C3491 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t77 GNDA 0.53137f
C3492 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n14 GNDA 0.35199f
C3493 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t39 GNDA 0.53137f
C3494 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n15 GNDA 0.35199f
C3495 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t90 GNDA 0.53137f
C3496 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n16 GNDA 0.35199f
C3497 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t98 GNDA 0.53137f
C3498 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n17 GNDA 0.35134f
C3499 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n18 GNDA 0.11998f
C3500 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t96 GNDA 0.5333f
C3501 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t89 GNDA 0.53137f
C3502 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n19 GNDA 0.70204f
C3503 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t68 GNDA 0.53137f
C3504 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n20 GNDA 0.35199f
C3505 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t41 GNDA 0.53137f
C3506 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n21 GNDA 0.35199f
C3507 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t92 GNDA 0.53137f
C3508 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n22 GNDA 0.35199f
C3509 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t91 GNDA 0.53137f
C3510 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n23 GNDA 0.35199f
C3511 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t64 GNDA 0.53137f
C3512 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n24 GNDA 0.35199f
C3513 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t95 GNDA 0.53137f
C3514 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n25 GNDA 0.35199f
C3515 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t94 GNDA 0.53137f
C3516 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n26 GNDA 0.35199f
C3517 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t81 GNDA 0.53137f
C3518 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n27 GNDA 0.35199f
C3519 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t65 GNDA 0.53137f
C3520 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n28 GNDA 0.35199f
C3521 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t38 GNDA 0.53137f
C3522 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n29 GNDA 0.2714f
C3523 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t27 GNDA 0.5333f
C3524 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t56 GNDA 0.53137f
C3525 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n30 GNDA 0.70204f
C3526 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t58 GNDA 0.53137f
C3527 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n31 GNDA 0.35199f
C3528 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t85 GNDA 0.53137f
C3529 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n32 GNDA 0.35199f
C3530 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t88 GNDA 0.53137f
C3531 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n33 GNDA 0.35199f
C3532 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t59 GNDA 0.53137f
C3533 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n34 GNDA 0.35199f
C3534 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t84 GNDA 0.53137f
C3535 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n35 GNDA 0.35199f
C3536 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t66 GNDA 0.53137f
C3537 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n36 GNDA 0.35134f
C3538 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n37 GNDA 0.08124f
C3539 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n38 GNDA 0.46703f
C3540 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t40 GNDA 0.5333f
C3541 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t28 GNDA 0.53137f
C3542 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n39 GNDA 0.70204f
C3543 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t87 GNDA 0.53137f
C3544 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n40 GNDA 0.35199f
C3545 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t62 GNDA 0.53137f
C3546 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n41 GNDA 0.35199f
C3547 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t33 GNDA 0.53137f
C3548 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n42 GNDA 0.35199f
C3549 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t29 GNDA 0.53137f
C3550 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n43 GNDA 0.35199f
C3551 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t78 GNDA 0.53137f
C3552 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n44 GNDA 0.35199f
C3553 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t37 GNDA 0.53137f
C3554 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n45 GNDA 0.35199f
C3555 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t35 GNDA 0.53137f
C3556 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n46 GNDA 0.35199f
C3557 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t101 GNDA 0.53137f
C3558 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n47 GNDA 0.35199f
C3559 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t79 GNDA 0.53137f
C3560 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n48 GNDA 0.35199f
C3561 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t52 GNDA 0.53137f
C3562 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n49 GNDA 0.2714f
C3563 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t42 GNDA 0.5333f
C3564 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t73 GNDA 0.53137f
C3565 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n50 GNDA 0.70204f
C3566 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t74 GNDA 0.53137f
C3567 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n51 GNDA 0.35199f
C3568 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t23 GNDA 0.53137f
C3569 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n52 GNDA 0.35199f
C3570 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t26 GNDA 0.53137f
C3571 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n53 GNDA 0.35199f
C3572 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t75 GNDA 0.53137f
C3573 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n54 GNDA 0.35199f
C3574 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t22 GNDA 0.53137f
C3575 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n55 GNDA 0.35199f
C3576 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t83 GNDA 0.53137f
C3577 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n56 GNDA 0.35134f
C3578 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n57 GNDA 0.08124f
C3579 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n58 GNDA 0.26714f
C3580 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t63 GNDA 0.5333f
C3581 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t50 GNDA 0.53137f
C3582 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n59 GNDA 0.70204f
C3583 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t34 GNDA 0.53137f
C3584 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n60 GNDA 0.35199f
C3585 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t80 GNDA 0.53137f
C3586 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n61 GNDA 0.35199f
C3587 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t54 GNDA 0.53137f
C3588 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n62 GNDA 0.35199f
C3589 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t51 GNDA 0.53137f
C3590 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n63 GNDA 0.35199f
C3591 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t24 GNDA 0.53137f
C3592 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n64 GNDA 0.35199f
C3593 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t57 GNDA 0.53137f
C3594 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n65 GNDA 0.35199f
C3595 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t55 GNDA 0.53137f
C3596 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n66 GNDA 0.35199f
C3597 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t43 GNDA 0.53137f
C3598 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n67 GNDA 0.35199f
C3599 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t25 GNDA 0.53137f
C3600 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n68 GNDA 0.35199f
C3601 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t76 GNDA 0.53137f
C3602 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n69 GNDA 0.2714f
C3603 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t70 GNDA 0.5333f
C3604 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t97 GNDA 0.53137f
C3605 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n70 GNDA 0.70204f
C3606 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t99 GNDA 0.53137f
C3607 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n71 GNDA 0.35199f
C3608 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t45 GNDA 0.53137f
C3609 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n72 GNDA 0.35199f
C3610 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t49 GNDA 0.53137f
C3611 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n73 GNDA 0.35199f
C3612 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t100 GNDA 0.53137f
C3613 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n74 GNDA 0.35199f
C3614 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t44 GNDA 0.53137f
C3615 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n75 GNDA 0.35199f
C3616 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t31 GNDA 0.53137f
C3617 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n76 GNDA 0.35134f
C3618 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n77 GNDA 0.08124f
C3619 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n78 GNDA 0.25098f
C3620 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t7 GNDA 0.13905f
C3621 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t12 GNDA 0.13905f
C3622 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n79 GNDA 0.71322f
C3623 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t16 GNDA 0.13905f
C3624 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t13 GNDA 0.13905f
C3625 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n80 GNDA 0.57542f
C3626 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n81 GNDA 0.85759f
C3627 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t17 GNDA 0.13905f
C3628 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t19 GNDA 0.13905f
C3629 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n82 GNDA 0.57542f
C3630 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n83 GNDA 0.53178f
C3631 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n84 GNDA 0.55633f
C3632 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t9 GNDA 0.13905f
C3633 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t2 GNDA 0.13905f
C3634 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n85 GNDA 0.71439f
C3635 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t10 GNDA 0.13905f
C3636 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t20 GNDA 0.13905f
C3637 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n86 GNDA 0.57542f
C3638 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n87 GNDA 0.85761f
C3639 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t5 GNDA 0.13905f
C3640 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t6 GNDA 0.13905f
C3641 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n88 GNDA 0.57542f
C3642 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n89 GNDA 0.3693f
C3643 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t21 GNDA 0.13952f
C3644 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t8 GNDA 0.36491f
C3645 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n90 GNDA 4.02968f
C3646 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n91 GNDA 0.36665f
C3647 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t3 GNDA 0.13905f
C3648 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t0 GNDA 0.13905f
C3649 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n92 GNDA 0.57542f
C3650 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n93 GNDA 0.44924f
C3651 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t1 GNDA 0.13905f
C3652 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t4 GNDA 0.13905f
C3653 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n94 GNDA 0.57542f
C3654 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n95 GNDA 1.10684f
C3655 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n96 GNDA 2.66466f
C3656 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t15 GNDA 0.13905f
C3657 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t18 GNDA 0.13905f
C3658 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n97 GNDA 0.57427f
C3659 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n98 GNDA 0.72111f
C3660 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t11 GNDA 0.13905f
C3661 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.t14 GNDA 0.13905f
C3662 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n99 GNDA 0.57542f
C3663 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n100 GNDA 0.61172f
C3664 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n101 GNDA 0.32496f
C3665 opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1.n102 GNDA 1.12763f
.ends

