** sch_path: /home/yohanes/10-bit-DAC/xschem/cm_pcell3.sch
.subckt cm_pcell3 VB1 VB2 ROUT VDDA
*.PININFO VDDA:I VB1:O VB2:O ROUT:O
XM1 VB2 net1 VB1 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=20 W=1.8 nf=1 m=2
XM2 net1 net1 VB2 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=20 W=1.8 nf=1 m=2
XM3 net2 ROUT net1 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=20 W=1.8 nf=1 m=2
XM4 ROUT ROUT net2 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=20 W=1.8 nf=1 m=2
XM5 VDDA VDDA VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1.8 nf=1 m=8
.ends
