magic
tech sky130A
magscale 1 2
timestamp 1750867770
<< error_s >>
rect 12930 -1959 12936 -1953
rect 12984 -1959 12990 -1953
rect 12924 -1965 12930 -1959
rect 12990 -1965 12996 -1959
<< metal1 >>
rect 9046 1081 9832 1109
rect 9045 1001 9744 1029
rect 8206 173 9656 201
rect 9056 141 9656 173
rect 9046 85 9304 113
rect 9056 53 9304 85
rect 9046 -3 9062 25
rect 9056 -35 9062 -3
rect 9122 -35 9128 25
rect 9046 -91 9216 -63
rect 9056 -123 9216 -91
rect 9056 -651 9062 -591
rect 9122 -651 9128 -591
rect 9056 -827 9062 -767
rect 9122 -827 9128 -767
rect 9056 -1059 9062 -1027
rect 9028 -1087 9062 -1059
rect 9122 -1087 9128 -1027
rect 9056 -1147 9062 -1115
rect 9027 -1175 9062 -1147
rect 9122 -1175 9128 -1115
rect 9156 -1471 9216 -123
rect 9156 -1537 9216 -1531
rect 9244 -1559 9304 53
rect 9508 25 9568 31
rect 9332 -591 9392 -585
rect 9332 -1295 9392 -651
rect 9332 -1361 9392 -1355
rect 9420 -767 9480 -761
rect 9420 -1383 9480 -827
rect 9508 -1207 9568 -35
rect 9596 -1119 9656 141
rect 9684 -1031 9744 1001
rect 9772 -943 9832 1081
rect 9772 -1009 9832 -1003
rect 9684 -1097 9744 -1091
rect 9596 -1185 9656 -1179
rect 9508 -1273 9568 -1267
rect 9420 -1449 9480 -1443
rect 9028 -1658 9062 -1598
rect 9122 -1658 9128 -1598
rect 9244 -1625 9304 -1619
rect 9028 -1663 9128 -1658
rect 9027 -1719 9062 -1691
rect 9056 -1751 9062 -1719
rect 9122 -1751 9128 -1691
rect 9784 -1779 9845 -1747
rect 9028 -1843 9845 -1779
rect 8865 -1875 9845 -1843
<< via1 >>
rect 9062 -35 9122 25
rect 9062 -651 9122 -591
rect 9062 -827 9122 -767
rect 9062 -1087 9122 -1027
rect 9062 -1175 9122 -1115
rect 9156 -1531 9216 -1471
rect 9508 -35 9568 25
rect 9332 -651 9392 -591
rect 9332 -1355 9392 -1295
rect 9420 -827 9480 -767
rect 9772 -1003 9832 -943
rect 9684 -1091 9744 -1031
rect 9596 -1179 9656 -1119
rect 9508 -1267 9568 -1207
rect 9420 -1443 9480 -1383
rect 9062 -1658 9122 -1598
rect 9244 -1619 9304 -1559
rect 9062 -1751 9122 -1691
<< metal2 >>
rect 9056 -35 9062 25
rect 9122 -35 9508 25
rect 9568 -35 9574 25
rect 9056 -651 9062 -591
rect 9122 -651 9332 -591
rect 9392 -651 9398 -591
rect 9056 -827 9062 -767
rect 9122 -827 9420 -767
rect 9480 -827 9486 -767
rect 9766 -1003 9772 -943
rect 9832 -1003 9845 -943
rect 9056 -1087 9062 -1027
rect 9122 -1032 9156 -1027
rect 9122 -1087 9166 -1032
rect 9156 -1088 9166 -1087
rect 9222 -1088 9232 -1032
rect 9678 -1091 9684 -1031
rect 9744 -1091 9845 -1031
rect 9056 -1175 9062 -1115
rect 9122 -1175 9128 -1115
rect 9068 -1219 9128 -1175
rect 9590 -1179 9596 -1119
rect 9656 -1179 9845 -1119
rect 9068 -1275 9166 -1219
rect 9222 -1275 9232 -1219
rect 9502 -1267 9508 -1207
rect 9568 -1267 9845 -1207
rect 9326 -1355 9332 -1295
rect 9392 -1355 9845 -1295
rect 9414 -1443 9420 -1383
rect 9480 -1443 9845 -1383
rect 9150 -1531 9156 -1471
rect 9216 -1531 9845 -1471
rect 9056 -1658 9062 -1598
rect 9122 -1602 9128 -1598
rect 9165 -1658 9175 -1602
rect 9238 -1619 9244 -1559
rect 9304 -1619 9845 -1559
rect 9056 -1663 9128 -1658
rect 5386 -1959 5542 -1843
rect 5570 -1959 5726 -1843
rect 5754 -1959 5818 -1843
rect 5846 -1959 5910 -1843
rect 5938 -1959 6002 -1843
rect 6030 -1959 6094 -1843
rect 8320 -1959 8384 -1843
rect 8412 -1959 8476 -1843
rect 8504 -1959 8568 -1843
rect 8596 -1959 8660 -1843
rect 8688 -1959 8844 -1731
rect 9056 -1751 9062 -1691
rect 9122 -1728 9128 -1691
rect 9056 -1784 9108 -1751
rect 9164 -1784 9174 -1728
rect 8872 -1959 9028 -1843
rect 12665 -4447 12725 -4387
rect 13309 -4447 13369 -4387
rect 13953 -4447 14013 -4387
rect 14597 -4447 14657 -4387
rect 15241 -4447 15301 -4387
rect 15885 -4447 15945 -4387
rect 16529 -4447 16589 -4387
rect 17173 -4447 17233 -4387
rect 17817 -4447 17877 -4387
rect 18461 -4447 18521 -4387
<< via2 >>
rect 9166 -1088 9222 -1032
rect 9166 -1275 9222 -1219
rect 9109 -1658 9122 -1602
rect 9122 -1658 9165 -1602
rect 9108 -1751 9122 -1728
rect 9122 -1751 9164 -1728
rect 9108 -1784 9164 -1751
<< metal3 >>
rect 9156 -1032 9232 -1027
rect 9156 -1088 9166 -1032
rect 9222 -1088 9232 -1032
rect 9156 -1094 9232 -1088
rect 9156 -1154 9845 -1094
rect 9156 -1219 9845 -1214
rect 9156 -1275 9166 -1219
rect 9222 -1274 9845 -1219
rect 9222 -1275 9232 -1274
rect 9156 -1280 9232 -1275
rect 9099 -1602 9175 -1597
rect 9099 -1658 9109 -1602
rect 9165 -1603 9175 -1602
rect 9165 -1658 9845 -1603
rect 9099 -1663 9845 -1658
rect 9098 -1728 9845 -1723
rect 9098 -1784 9108 -1728
rect 9164 -1783 9845 -1728
rect 9164 -1784 9174 -1783
rect 9098 -1789 9174 -1784
<< comment >>
rect 12575 -4143 12673 -4102
use dcell_buffer_bus  dcell_buffer_bus_0 ~/10-bit-DAC/mag
timestamp 1750863581
transform 1 0 0 0 1 0
box 5366 -4551 25377 -1953
use dcell_lv  dcell_lv_0 ~/10-bit-DAC/mag
timestamp 1750867770
transform 1 0 5395 0 1 -747
box -9 -1096 3665 1886
<< labels >>
flabel metal2 s 18461 -4447 18521 -4387 0 FreeSans 160 180 0 0 DIN0
port 0 nsew
flabel metal2 s 17817 -4447 17877 -4387 0 FreeSans 160 180 0 0 DIN1
port 1 nsew
flabel metal2 s 17173 -4447 17233 -4387 0 FreeSans 160 180 0 0 DIN2
port 2 nsew
flabel metal2 s 16529 -4447 16589 -4387 0 FreeSans 160 180 0 0 DIN3
port 3 nsew
flabel metal2 s 15885 -4447 15945 -4387 0 FreeSans 160 180 0 0 DIN4
port 4 nsew
flabel metal2 s 15241 -4447 15301 -4387 0 FreeSans 160 180 0 0 DIN5
port 5 nsew
flabel metal2 s 14597 -4447 14657 -4387 0 FreeSans 160 180 0 0 DIN6
port 6 nsew
flabel metal2 s 13953 -4447 14013 -4387 0 FreeSans 160 180 0 0 DIN7
port 7 nsew
flabel metal2 s 13309 -4447 13369 -4387 0 FreeSans 160 180 0 0 DIN8
port 8 nsew
flabel metal2 s 12665 -4447 12725 -4387 0 FreeSans 160 180 0 0 DIN9
port 9 nsew
flabel metal2 s 9244 -1619 9304 -1559 0 FreeSans 160 0 0 0 S[1]
port 10 nsew
flabel metal2 s 9420 -1443 9480 -1383 0 FreeSans 160 0 0 0 S[2]
port 11 nsew
flabel metal2 s 9596 -1179 9656 -1119 0 FreeSans 160 0 0 0 S[3]
port 12 nsew
flabel metal2 s 9772 -1003 9832 -943 0 FreeSans 160 0 0 0 S[4]
port 13 nsew
flabel metal2 s 9156 -1531 9216 -1471 0 FreeSans 160 0 0 0 SB[1]
port 14 nsew
flabel metal2 s 9332 -1355 9392 -1295 0 FreeSans 160 0 0 0 SB[2]
port 15 nsew
flabel metal2 s 9508 -1267 9568 -1207 0 FreeSans 160 0 0 0 SB[3]
port 16 nsew
flabel metal2 s 9684 -1091 9744 -1031 0 FreeSans 160 0 0 0 SB[4]
port 17 nsew
flabel metal2 s 9062 -1751 9122 -1691 0 FreeSans 160 0 0 0 DS[8]
port 18 nsew
flabel metal2 s 9062 -1175 9122 -1115 0 FreeSans 160 0 0 0 DS[9]
port 19 nsew
flabel metal2 s 9062 -1658 9122 -1598 0 FreeSans 160 0 0 0 DSB[8]
port 20 nsew
flabel metal2 s 9062 -1087 9122 -1027 0 FreeSans 160 0 0 0 DSB[9]
port 21 nsew
flabel metal1 s 12457 -3840 12457 -3840 0 FreeSans 160 0 0 0 VDD
port 22 nsew
flabel metal1 s 12504 -4447 12504 -4447 0 FreeSans 160 0 0 0 GND
port 23 nsew
<< end >>
