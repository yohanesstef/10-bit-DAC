magic
tech sky130A
magscale 1 2
timestamp 1749007001
<< xpolycontact >>
rect -141 460 141 892
rect -141 -892 141 -460
<< xpolyres >>
rect -141 -460 141 460
<< viali >>
rect -125 477 125 874
rect -125 -874 125 -477
<< metal1 >>
rect -131 874 131 886
rect -131 477 -125 874
rect 125 477 131 874
rect -131 465 131 477
rect -131 -477 131 -465
rect -131 -874 -125 -477
rect 125 -874 131 -477
rect -131 -886 131 -874
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 4.757 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 7.014k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
