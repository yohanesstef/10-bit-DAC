magic
tech sky130A
magscale 1 2
timestamp 1750064919
<< error_s >>
rect -254 1208 798 1274
rect -254 -29 -188 1208
rect -128 1119 672 1148
rect -128 0 -51 1119
rect -15 63 15 1019
rect 529 63 559 1019
rect -15 59 559 63
rect 595 0 672 1119
rect -128 -3 -62 0
rect 606 -3 672 0
rect -128 -7 672 -3
rect -128 -29 -62 -7
rect -254 -95 -62 -29
rect 606 -29 672 -7
rect 732 -29 798 1208
rect 606 -95 798 -29
<< magnet >>
rect 662 1161 719 1195
rect 685 1104 719 1161
<< mvnsubdiff >>
rect -188 1148 732 1208
rect -188 -29 -128 1148
rect 672 -29 732 1148
<< poly >>
rect -90 33 -30 1116
rect 574 33 634 1116
<< locali >>
rect -175 1161 719 1195
rect -175 -29 -141 1161
rect 685 -29 719 1161
<< metal1 >>
rect -198 1138 742 1218
rect -198 -29 -118 1138
rect -9 951 37 1138
rect 218 1060 295 1106
rect 476 1060 553 1106
rect 249 1019 295 1060
rect 507 1019 553 1060
rect 507 31 553 59
rect -9 -29 553 31
rect 662 -29 742 1138
use sky130_fd_pr__pfet_g5v0d10v5_XEEY48  sky130_fd_pr__pfet_g5v0d10v5_XEEY48_0
timestamp 1750064013
transform 1 0 272 0 1 575
box -353 -582 353 544
<< end >>
