magic
tech sky130A
magscale 1 2
timestamp 1750150351
<< metal1 >>
rect 36114 1975 36211 2035
tri 36211 1975 36271 2035 sw
rect 36331 1975 36337 2035
rect 36397 1975 36403 2035
rect 36114 1855 36120 1915
rect 36180 1855 36186 1915
tri 36186 1890 36271 1975 ne
tri 36271 1915 36331 1975 sw
rect 36271 1890 36403 1915
tri 36271 1855 36306 1890 ne
rect 36306 1855 36403 1890
<< via1 >>
rect 36337 1975 36397 2035
rect 36120 1855 36180 1915
<< metal2 >>
tri 36271 2000 36306 2035 se
rect 36306 2000 36337 2035
tri 36186 1915 36271 2000 se
rect 36271 1975 36337 2000
rect 36397 1975 36403 2035
tri 36271 1915 36331 1975 nw
rect 36114 1855 36120 1915
rect 36180 1855 36211 1915
tri 36211 1855 36271 1915 nw
<< end >>
