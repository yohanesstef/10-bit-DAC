magic
tech sky130A
magscale 1 2
timestamp 1750150351
<< pwell >>
rect -45 -846 1585 816
<< mvpsubdiffcont >>
rect 4 -737 38 707
rect 1502 -737 1536 707
rect 64 -797 1476 -763
<< metal1 >>
rect 688 597 734 685
rect 793 625 799 685
rect 859 625 865 685
rect 675 537 681 597
rect 741 537 747 597
rect 806 541 852 625
rect 688 536 734 537
rect 430 75 476 103
rect 1064 75 1110 103
rect 430 15 626 75
rect 915 15 1044 75
rect 1104 15 1110 75
rect 1219 -45 1279 692
rect 430 -105 626 -45
rect 915 -105 1044 -45
rect 1104 -105 1110 -45
rect 430 -133 476 -105
rect 1064 -133 1110 -105
rect 1219 -111 1279 -105
rect 1307 75 1367 692
rect 1307 -111 1367 15
rect 675 -619 681 -559
rect 741 -619 747 -559
rect 688 -707 734 -619
rect 806 -647 852 -526
rect 793 -707 799 -647
rect 859 -707 865 -647
<< via1 >>
rect 261 625 321 685
rect 799 625 859 685
rect 173 537 233 597
rect 681 537 741 597
rect 1044 15 1104 75
rect 1044 -105 1104 -45
rect 1219 -105 1279 -45
rect 1307 15 1367 75
rect 261 -619 321 -559
rect 681 -619 741 -559
rect 173 -707 233 -647
rect 799 -707 859 -647
<< metal2 >>
rect 167 625 261 685
rect 321 625 799 685
rect 859 625 865 685
rect 167 537 173 597
rect 233 537 681 597
rect 741 537 865 597
rect 1038 15 1044 75
rect 1104 15 1307 75
rect 1367 15 1373 75
rect 1038 -105 1044 -45
rect 1104 -105 1219 -45
rect 1279 -105 1373 -45
rect 167 -619 261 -559
rect 321 -619 681 -559
rect 741 -619 865 -559
rect 167 -707 173 -647
rect 233 -707 799 -647
rect 859 -707 865 -647
use cross_pair  cross_pair_0
timestamp 1750150351
transform 1 0 -35488 0 1 -1960
box 36114 1855 36403 2035
use fc_ncell2_2  fc_ncell2_2_0
timestamp 1750017694
transform 1 0 431 0 1 67
box -440 -82 1118 713
use fc_ncell2_2  fc_ncell2_2_1
timestamp 1750017694
transform 1 0 431 0 -1 -97
box -440 -82 1118 713
<< end >>
