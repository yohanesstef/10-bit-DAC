magic
tech sky130A
magscale 1 2
timestamp 1749465145
<< error_s >>
rect 24468 -18552 24474 -18546
rect 24522 -18552 24528 -18546
rect 24462 -18558 24468 -18552
rect 24528 -18558 24534 -18552
<< pwell >>
rect 12802 -21608 26239 -18026
<< psubdiff >>
rect 12838 -18122 13098 -18062
rect 25943 -18122 26203 -18062
rect 12838 -18322 12898 -18122
rect 12838 -21512 12898 -21312
rect 26143 -18322 26203 -18122
rect 26143 -21512 26203 -21312
rect 12838 -21572 13098 -21512
rect 25943 -21572 26203 -21512
<< psubdiffcont >>
rect 13098 -18122 25943 -18062
rect 12838 -21312 12898 -18322
rect 26143 -21312 26203 -18322
rect 13098 -21572 25943 -21512
<< locali >>
rect 12838 -18122 13098 -18062
rect 25943 -18122 26203 -18062
rect 12838 -18322 12898 -18122
rect 13252 -18218 13684 -18122
rect 13762 -18218 14194 -18122
rect 14826 -18218 15258 -18122
rect 15358 -18218 15790 -18122
rect 16334 -18218 16766 -18122
rect 16876 -18218 17308 -18122
rect 17945 -18218 18377 -18122
rect 18507 -18218 18939 -18122
rect 19488 -18218 19920 -18122
rect 20060 -18218 20492 -18122
rect 21124 -18218 21556 -18122
rect 21768 -18218 22200 -18122
rect 22744 -18218 23176 -18122
rect 23398 -18218 23830 -18122
rect 24462 -18218 24894 -18122
rect 25372 -18218 25804 -18122
rect 26143 -18322 26203 -18122
rect 24462 -18542 24894 -18500
rect 25372 -18542 25804 -18500
rect 12838 -21512 12898 -21312
rect 13246 -21512 13678 -21416
rect 13768 -21512 14200 -21416
rect 14831 -21512 15263 -21416
rect 15353 -21512 15785 -21416
rect 16329 -21512 16761 -21416
rect 16881 -21512 17313 -21416
rect 17950 -21512 18382 -21416
rect 18502 -21512 18934 -21416
rect 19472 -21512 19904 -21416
rect 20076 -21512 20508 -21416
rect 21144 -21512 21576 -21416
rect 21748 -21512 22180 -21416
rect 22708 -21512 23140 -21416
rect 23434 -21512 23866 -21416
rect 24544 -21512 24976 -21416
rect 25290 -21512 25722 -21416
rect 26143 -21512 26203 -21312
rect 12838 -21572 13098 -21512
rect 25943 -21572 26203 -21512
<< via1 >>
rect 14122 -18814 14182 -18552
rect 15718 -18814 15778 -18552
rect 17236 -18814 17296 -18552
rect 18867 -18814 18927 -18552
rect 20420 -18814 20480 -18552
rect 22128 -18814 22188 -18552
rect 23758 -18814 23818 -18552
rect 24468 -18814 24528 -18552
rect 14474 -21082 14534 -20820
rect 15713 -21082 15773 -20820
rect 17588 -21082 17648 -20820
rect 18862 -21082 18922 -20820
rect 20772 -21082 20832 -20820
rect 22108 -21082 22168 -20820
rect 24110 -21082 24170 -20820
rect 25650 -21082 25710 -20820
<< metal2 >>
rect 12802 -18814 14122 -18552
rect 14182 -18814 14188 -18552
rect 15712 -18814 15718 -18552
rect 15778 -18814 17236 -18552
rect 17296 -18814 17302 -18552
rect 18861 -18814 18867 -18552
rect 18927 -18814 20420 -18552
rect 20480 -18814 20486 -18552
rect 22122 -18814 22128 -18552
rect 22188 -18814 23758 -18552
rect 23818 -18814 23824 -18552
rect 24462 -18814 24468 -18552
rect 24528 -18814 26239 -18552
rect 14468 -21082 14474 -20820
rect 14534 -21082 15713 -20820
rect 15773 -21082 15779 -20820
rect 17582 -21082 17588 -20820
rect 17648 -21082 18862 -20820
rect 18922 -21082 18928 -20820
rect 20766 -21082 20772 -20820
rect 20832 -21082 22108 -20820
rect 22168 -21082 22174 -20820
rect 24104 -21082 24110 -20820
rect 24170 -21082 25650 -20820
rect 25710 -21082 25716 -20820
use rseg_4_1  rseg_4_1_0
timestamp 1749369846
transform 1 0 11667 0 1 4554
box 1327 -25970 2873 -22772
use rseg_4_2  rseg_4_2_0
timestamp 1749369846
transform 1 0 10449 0 1 4573
box 4119 -25989 5599 -22791
use rseg_4_3  rseg_4_3_0
timestamp 1749369846
transform 1 0 8582 0 1 4696
box 7494 -26112 9072 -22914
use rseg_4_4  rseg_4_4_0
timestamp 1749369846
transform 1 0 6286 0 1 4832
box 11396 -26248 12911 -23050
use rseg_4_5  rseg_4_5_0
timestamp 1749369846
transform 1 0 4494 0 1 4812
box 14731 -26228 16344 -23030
use rseg_4_6  rseg_4_6_0
timestamp 1749369846
transform 1 0 3186 0 1 4844
box 17680 -26260 19272 -23062
use rseg_4_7  rseg_4_7_0
timestamp 1749369846
transform 1 0 1778 0 1 4879
box 20708 -26295 22398 -23097
use rseg_4_8  rseg_4_8_0
timestamp 1749369846
transform 1 0 400 0 1 4877
box 23804 -26293 25647 -23095
<< labels >>
flabel metal1 s 13258 -18552 13258 -18552 2 FreeSans 240 0 0 0 v1
port 1 ne
flabel metal1 s 14216 -18552 14216 -18552 2 FreeSans 240 0 0 0 v2
port 2 ne
flabel metal1 s 13170 -18552 13170 -18552 2 FreeSans 240 0 0 0 v3
port 3 ne
flabel metal1 s 14304 -18552 14304 -18552 2 FreeSans 240 0 0 0 v4
port 4 ne
flabel metal1 s 13082 -18552 13082 -18552 2 FreeSans 240 0 0 0 v5
port 5 ne
flabel metal1 s 14392 -18552 14392 -18552 2 FreeSans 240 0 0 0 v6
port 6 ne
flabel metal1 s 12994 -18552 12994 -18552 2 FreeSans 240 0 0 0 v7
port 7 ne
flabel metal1 s 14480 -18552 14480 -18552 2 FreeSans 240 0 0 0 v8
port 8 ne
flabel metal1 s 14568 -18552 14568 -18552 2 FreeSans 240 0 0 0 v9
port 9 ne
flabel metal1 s 15988 -18552 15988 -18552 2 FreeSans 240 0 0 0 v10
port 10 ne
flabel metal1 s 14656 -18552 14656 -18552 2 FreeSans 240 0 0 0 v11
port 11 ne
flabel metal1 s 15900 -18552 15900 -18552 2 FreeSans 240 0 0 0 v12
port 12 ne
flabel metal1 s 14744 -18552 14744 -18552 2 FreeSans 240 0 0 0 v13
port 13 ne
flabel metal1 s 15812 -18552 15812 -18552 2 FreeSans 240 0 0 0 v14
port 14 ne
flabel metal1 s 14832 -18552 14832 -18552 2 FreeSans 240 0 0 0 v15
port 15 ne
flabel metal1 s 15724 -18552 15724 -18552 2 FreeSans 240 0 0 0 v16
port 16 ne
flabel metal1 s 16340 -18552 16340 -18552 2 FreeSans 240 0 0 0 v17
port 17 ne
flabel metal1 s 17330 -18552 17330 -18552 2 FreeSans 240 0 0 0 v18
port 18 ne
flabel metal1 s 16252 -18552 16252 -18552 2 FreeSans 240 0 0 0 v19
port 19 ne
flabel metal1 s 17418 -18552 17418 -18552 2 FreeSans 240 0 0 0 v20
port 20 ne
flabel metal1 s 16164 -18552 16164 -18552 2 FreeSans 240 0 0 0 v21
port 21 ne
flabel metal1 s 17506 -18552 17506 -18552 2 FreeSans 240 0 0 0 v22
port 22 ne
flabel metal1 s 16076 -18552 16076 -18552 2 FreeSans 240 0 0 0 v23
port 23 ne
flabel metal1 s 17594 -18552 17594 -18552 2 FreeSans 240 0 0 0 v24
port 24 ne
flabel metal1 s 17682 -18552 17682 -18552 2 FreeSans 240 0 0 0 v25
port 25 ne
flabel metal1 s 19137 -18552 19137 -18552 2 FreeSans 240 0 0 0 v26
port 26 ne
flabel metal1 s 17770 -18552 17770 -18552 2 FreeSans 240 0 0 0 v27
port 27 ne
flabel metal1 s 19049 -18552 19049 -18552 2 FreeSans 240 0 0 0 v28
port 28 ne
flabel metal1 s 17858 -18552 17858 -18552 2 FreeSans 240 0 0 0 v29
port 29 ne
flabel metal1 s 18961 -18552 18961 -18552 2 FreeSans 240 0 0 0 v30
port 30 ne
flabel metal1 s 18873 -18552 18873 -18552 2 FreeSans 240 0 0 0 v32
port 32 ne
flabel metal1 s 20514 -18552 20514 -18552 2 FreeSans 240 0 0 0 v34
port 34 ne
flabel metal1 s 19401 -18552 19401 -18552 2 FreeSans 240 0 0 0 v35
port 35 ne
flabel metal1 s 20602 -18552 20602 -18552 2 FreeSans 240 0 0 0 v36
port 36 ne
flabel metal1 s 19313 -18552 19313 -18552 2 FreeSans 240 0 0 0 v37
port 37 ne
flabel metal1 s 20690 -18552 20690 -18552 2 FreeSans 240 0 0 0 v38
port 38 ne
flabel metal1 s 19225 -18552 19225 -18552 2 FreeSans 240 0 0 0 v39
port 39 ne
flabel metal1 s 20778 -18552 20778 -18552 2 FreeSans 240 0 0 0 v40
port 40 ne
flabel metal1 s 20866 -18552 20866 -18552 2 FreeSans 240 0 0 0 v41
port 41 ne
flabel metal1 s 22398 -18552 22398 -18552 2 FreeSans 240 0 0 0 v42
port 42 ne
flabel metal1 s 20954 -18552 20954 -18552 2 FreeSans 240 0 0 0 v43
port 43 ne
flabel metal1 s 22310 -18552 22310 -18552 2 FreeSans 240 0 0 0 v44
port 44 ne
flabel metal1 s 21042 -18552 21042 -18552 2 FreeSans 240 0 0 0 v45
port 45 ne
flabel metal1 s 22222 -18552 22222 -18552 2 FreeSans 240 0 0 0 v46
port 46 ne
flabel metal1 s 21130 -18552 21130 -18552 2 FreeSans 240 0 0 0 v47
port 47 ne
flabel metal1 s 22134 -18552 22134 -18552 2 FreeSans 240 0 0 0 v48
port 48 ne
flabel metal1 s 22750 -18552 22750 -18552 2 FreeSans 240 0 0 0 v49
port 49 ne
flabel metal1 s 23852 -18552 23852 -18552 2 FreeSans 240 0 0 0 v50
port 50 ne
flabel metal1 s 22662 -18552 22662 -18552 2 FreeSans 240 0 0 0 v51
port 51 ne
flabel metal1 s 23940 -18552 23940 -18552 2 FreeSans 240 0 0 0 v52
port 52 ne
flabel metal1 s 22574 -18552 22574 -18552 2 FreeSans 240 0 0 0 v53
port 53 ne
flabel metal1 s 24028 -18552 24028 -18552 2 FreeSans 240 0 0 0 v54
port 54 ne
flabel metal1 s 22486 -18552 22486 -18552 2 FreeSans 240 0 0 0 v55
port 55 ne
flabel metal1 s 24116 -18552 24116 -18552 2 FreeSans 240 0 0 0 v56
port 56 ne
flabel metal1 s 24204 -18552 24204 -18552 2 FreeSans 240 0 0 0 v57
port 57 ne
flabel metal1 s 25987 -18552 25987 -18552 2 FreeSans 240 0 0 0 v58
port 58 ne
flabel metal1 s 24292 -18552 24292 -18552 2 FreeSans 240 0 0 0 v59
port 59 ne
flabel metal1 s 25899 -18552 25899 -18552 2 FreeSans 240 0 0 0 v60
port 60 ne
flabel metal1 s 24380 -18552 24380 -18552 2 FreeSans 240 0 0 0 v61
port 61 ne
flabel metal1 s 25811 -18552 25811 -18552 2 FreeSans 240 0 0 0 v62
port 62 ne
flabel metal1 s 19494 -18552 19494 -18552 2 FreeSans 240 0 0 0 v33
port 33 ne
flabel metal1 s 17951 -18552 17951 -18552 2 FreeSans 240 0 0 0 v31
port 31 ne
<< end >>
