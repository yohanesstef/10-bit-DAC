magic
tech sky130A
magscale 1 2
timestamp 1748966771
<< xpolycontact >>
rect -141 171 141 603
rect -141 -603 141 -171
<< xpolyres >>
rect -141 -171 141 171
<< viali >>
rect -125 188 125 585
rect -125 -585 125 -188
<< metal1 >>
rect -131 585 131 597
rect -131 188 -125 585
rect 125 188 131 585
rect -131 176 131 188
rect -131 -188 131 -176
rect -131 -585 -125 -188
rect 125 -585 131 -188
rect -131 -597 131 -585
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.8655599999 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 2.913k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
