magic
tech sky130A
magscale 1 2
timestamp 1750079478
<< error_s >>
rect 1019 1476 1025 1482
rect 1073 1476 1079 1482
rect 1137 1476 1143 1482
rect 1191 1476 1197 1482
rect 2523 1476 2529 1482
rect 2577 1476 2583 1482
rect 2641 1476 2647 1482
rect 2695 1476 2701 1482
rect 1013 1470 1019 1476
rect 1079 1470 1085 1476
rect 1131 1470 1137 1476
rect 1197 1470 1203 1476
rect 2517 1470 2523 1476
rect 2583 1470 2589 1476
rect 2635 1470 2641 1476
rect 2701 1470 2707 1476
rect 1013 1416 1019 1422
rect 1079 1416 1085 1422
rect 1131 1416 1137 1422
rect 1197 1416 1203 1422
rect 2517 1416 2523 1422
rect 2583 1416 2589 1422
rect 2635 1416 2641 1422
rect 2701 1416 2707 1422
rect 1019 1410 1025 1416
rect 1073 1410 1079 1416
rect 1137 1410 1143 1416
rect 1191 1410 1197 1416
rect 2523 1410 2529 1416
rect 2577 1410 2583 1416
rect 2641 1410 2647 1416
rect 2695 1410 2701 1416
rect 267 1388 273 1394
rect 321 1388 327 1394
rect 385 1388 391 1394
rect 439 1388 445 1394
rect 1771 1388 1777 1394
rect 1825 1388 1831 1394
rect 1889 1388 1895 1394
rect 1943 1388 1949 1394
rect 261 1382 267 1388
rect 327 1382 333 1388
rect 379 1382 385 1388
rect 445 1382 451 1388
rect 1765 1382 1771 1388
rect 1831 1382 1837 1388
rect 1883 1382 1889 1388
rect 1949 1382 1955 1388
rect 261 1328 267 1334
rect 327 1328 333 1334
rect 379 1328 385 1334
rect 445 1328 451 1334
rect 1765 1328 1771 1334
rect 1831 1328 1837 1334
rect 1883 1328 1889 1334
rect 1949 1328 1955 1334
rect 267 1322 273 1328
rect 321 1322 327 1328
rect 385 1322 391 1328
rect 439 1322 445 1328
rect 1771 1322 1777 1328
rect 1825 1322 1831 1328
rect 1889 1322 1895 1328
rect 1943 1322 1949 1328
rect 761 1300 767 1306
rect 815 1300 821 1306
rect 1395 1300 1401 1306
rect 1449 1300 1455 1306
rect 2265 1300 2271 1306
rect 2319 1300 2325 1306
rect 2899 1300 2905 1306
rect 2953 1300 2959 1306
rect 755 1294 761 1300
rect 821 1294 827 1300
rect 1389 1294 1395 1300
rect 1455 1294 1461 1300
rect 2259 1294 2265 1300
rect 2325 1294 2331 1300
rect 2893 1294 2899 1300
rect 2959 1294 2965 1300
rect 755 1240 761 1246
rect 821 1240 827 1246
rect 1389 1240 1395 1246
rect 1455 1240 1461 1246
rect 2259 1240 2265 1246
rect 2325 1240 2331 1246
rect 2893 1240 2899 1246
rect 2959 1240 2965 1246
rect 761 1234 767 1240
rect 815 1234 821 1240
rect 1395 1234 1401 1240
rect 1449 1234 1455 1240
rect 2265 1234 2271 1240
rect 2319 1234 2325 1240
rect 2899 1234 2905 1240
rect 2953 1234 2959 1240
rect 9 1212 15 1218
rect 63 1212 69 1218
rect 643 1212 649 1218
rect 697 1212 703 1218
rect 1513 1212 1519 1218
rect 1567 1212 1573 1218
rect 2147 1212 2153 1218
rect 2201 1212 2207 1218
rect 3 1206 9 1212
rect 69 1206 75 1212
rect 637 1206 643 1212
rect 703 1206 709 1212
rect 1507 1206 1513 1212
rect 1573 1206 1579 1212
rect 2141 1206 2147 1212
rect 2207 1206 2213 1212
rect 3 1152 9 1158
rect 69 1152 75 1158
rect 637 1152 643 1158
rect 703 1152 709 1158
rect 1507 1152 1513 1158
rect 1573 1152 1579 1158
rect 2141 1152 2147 1158
rect 2207 1152 2213 1158
rect 9 1146 15 1152
rect 63 1146 69 1152
rect 643 1146 649 1152
rect 697 1146 703 1152
rect 1513 1146 1519 1152
rect 1567 1146 1573 1152
rect 2147 1146 2153 1152
rect 2201 1146 2207 1152
rect 643 860 649 866
rect 697 860 703 866
rect 761 860 767 866
rect 815 860 821 866
rect 637 854 643 860
rect 703 854 709 860
rect 755 854 761 860
rect 821 854 827 860
rect 637 800 643 806
rect 703 800 709 806
rect 755 800 761 806
rect 821 800 827 806
rect 643 794 649 800
rect 697 794 703 800
rect 761 794 767 800
rect 815 794 821 800
rect 1395 772 1401 778
rect 1449 772 1455 778
rect 1513 772 1519 778
rect 1567 772 1573 778
rect 1389 766 1395 772
rect 1455 766 1461 772
rect 1507 766 1513 772
rect 1573 766 1579 772
rect 1389 712 1395 718
rect 1455 712 1461 718
rect 1507 712 1513 718
rect 1573 712 1579 718
rect 1395 706 1401 712
rect 1449 706 1455 712
rect 1513 706 1519 712
rect 1567 706 1573 712
rect 385 684 391 690
rect 439 684 445 690
rect 1019 684 1025 690
rect 1073 684 1079 690
rect 379 678 385 684
rect 445 678 451 684
rect 1013 678 1019 684
rect 1079 678 1085 684
rect 379 624 385 630
rect 445 624 451 630
rect 1013 624 1019 630
rect 1079 624 1085 630
rect 385 618 391 624
rect 439 618 445 624
rect 1019 618 1025 624
rect 1073 618 1079 624
rect 1137 596 1143 602
rect 1191 596 1197 602
rect 1771 596 1777 602
rect 1825 596 1831 602
rect 1131 590 1137 596
rect 1197 590 1203 596
rect 1765 590 1771 596
rect 1831 590 1837 596
rect 1131 536 1137 542
rect 1197 536 1203 542
rect 1765 536 1771 542
rect 1831 536 1837 542
rect 1137 530 1143 536
rect 1191 530 1197 536
rect 1771 530 1777 536
rect 1825 530 1831 536
rect 9 156 15 162
rect 63 156 69 162
rect 3 150 9 156
rect 69 150 75 156
rect 3 96 9 102
rect 69 96 75 102
rect 9 90 15 96
rect 63 90 69 96
<< metal1 >>
rect 1013 1416 1019 1476
rect 1079 1416 1085 1476
rect 1131 1416 1137 1476
rect 1197 1416 1203 1476
rect 2517 1416 2523 1476
rect 2583 1416 2589 1476
rect 2635 1416 2641 1476
rect 2701 1416 2707 1476
rect 261 1328 267 1388
rect 327 1328 333 1388
rect 379 1328 385 1388
rect 445 1328 451 1388
rect 3 1152 9 1212
rect 69 1152 75 1212
rect 16 1034 62 1152
rect 274 1046 320 1328
rect 392 926 438 1328
rect 755 1240 761 1300
rect 821 1240 827 1300
rect 637 1152 643 1212
rect 703 1152 709 1212
rect 650 1046 696 1152
rect 768 1046 814 1240
rect 1026 926 1072 1416
rect 1144 926 1190 1416
rect 1765 1328 1771 1388
rect 1831 1328 1837 1388
rect 1883 1328 1889 1388
rect 1949 1328 1955 1388
rect 1389 1240 1395 1300
rect 1455 1240 1461 1300
rect 1402 1034 1448 1240
rect 1507 1152 1513 1212
rect 1573 1152 1579 1212
rect 1520 1034 1566 1152
rect 1778 927 1824 1328
rect 1896 927 1942 1328
rect 2259 1240 2265 1300
rect 2325 1240 2331 1300
rect 2141 1152 2147 1212
rect 2207 1152 2213 1212
rect 2154 1034 2200 1152
rect 2272 1034 2318 1240
rect 2530 986 2576 1416
rect 2648 986 2694 1416
rect 2893 1240 2899 1300
rect 2959 1240 2965 1300
rect 2906 1034 2952 1240
rect 637 800 643 860
rect 703 800 709 860
rect 755 800 761 860
rect 821 800 827 860
rect 379 624 385 684
rect 445 624 451 684
rect 650 646 696 800
rect 16 156 62 526
rect 274 332 320 533
rect 768 526 814 800
rect 1389 712 1395 772
rect 1455 712 1461 772
rect 1507 712 1513 772
rect 1573 712 1579 772
rect 2272 734 2318 938
rect 1013 624 1019 684
rect 1079 624 1085 684
rect 1402 646 1448 712
rect 1026 583 1072 624
rect 1131 536 1137 596
rect 1197 536 1203 596
rect 1520 526 1566 712
rect 1896 674 2318 734
rect 2394 926 2694 986
rect 1896 634 1942 674
rect 2394 646 2454 926
rect 1765 536 1771 596
rect 1831 536 1837 596
rect 2154 586 2454 646
rect 1896 420 1942 538
rect 2530 420 2576 616
rect 1896 360 2576 420
rect 261 272 267 332
rect 327 272 333 332
rect 3 96 9 156
rect 69 96 75 156
<< via1 >>
rect 1019 1416 1079 1476
rect 1137 1416 1197 1476
rect 2523 1416 2583 1476
rect 2641 1416 2701 1476
rect 267 1328 327 1388
rect 385 1328 445 1388
rect 9 1152 69 1212
rect 761 1240 821 1300
rect 643 1152 703 1212
rect 1771 1328 1831 1388
rect 1889 1328 1949 1388
rect 1395 1240 1455 1300
rect 1513 1152 1573 1212
rect 2265 1240 2325 1300
rect 2147 1152 2207 1212
rect 2899 1240 2959 1300
rect 643 800 703 860
rect 761 800 821 860
rect 385 624 445 684
rect 1395 712 1455 772
rect 1513 712 1573 772
rect 1019 624 1079 684
rect 1137 536 1197 596
rect 1771 536 1831 596
rect 267 272 327 332
rect 9 96 69 156
<< metal2 >>
rect 261 272 267 332
rect 327 272 333 332
use cm_ncell2_cell  cm_ncell2_cell_0
timestamp 1750079478
transform 1 0 -16 0 1 -4
box -4 -8 3506 1588
<< end >>
