magic
tech sky130A
magscale 1 2
timestamp 1749538868
<< metal1 >>
rect 15177 -23125 15237 -21181
rect 15265 -22477 15325 -21181
rect 15353 -21829 15413 -21181
rect 15454 -21505 15862 -21443
rect 16493 -21505 16553 -21181
rect 16465 -21767 16553 -21505
rect 16044 -21829 16465 -21767
rect 15353 -22091 15441 -21829
rect 15454 -22131 15862 -22091
rect 15447 -22153 15862 -22131
rect 16581 -22153 16641 -21181
rect 16459 -22414 16641 -22153
rect 16459 -22415 16605 -22414
rect 16038 -22477 16454 -22415
rect 15265 -22739 15452 -22477
rect 15452 -22801 15868 -22739
rect 16669 -22801 16729 -21181
rect 16459 -23063 16729 -22801
rect 16038 -23125 16454 -23063
rect 15177 -23387 15452 -23125
rect 15457 -23449 15873 -23387
rect 16757 -23449 16817 -21181
rect 16449 -23711 16817 -23449
use sky130_fd_pr__res_xhigh_po_1p41_6E4UWG  sky130_fd_pr__res_xhigh_po_1p41_6E4UWG_0
timestamp 1749204500
transform 0 -1 15953 1 0 -23904
box -141 -502 141 502
use sky130_fd_pr__res_xhigh_po_1p41_355JL6  sky130_fd_pr__res_xhigh_po_1p41_355JL6_0
timestamp 1748944356
transform 0 -1 15953 1 0 -21960
box -141 -518 141 518
use sky130_fd_pr__res_xhigh_po_1p41_355LL6  sky130_fd_pr__res_xhigh_po_1p41_355LL6_0
timestamp 1749204500
transform 0 -1 15953 1 0 -20988
box -141 -518 141 518
use sky130_fd_pr__res_xhigh_po_1p41_VXMCTQ  sky130_fd_pr__res_xhigh_po_1p41_VXMCTQ_0
timestamp 1748944356
transform 0 -1 15953 1 0 -22932
box -141 -512 141 512
use sky130_fd_pr__res_xhigh_po_1p41_355JL6  XR33
timestamp 1748944356
transform 0 -1 15953 1 0 -21312
box -141 -518 141 518
use sky130_fd_pr__res_xhigh_po_1p41_355JL6  XR34
timestamp 1748944356
transform 0 -1 15953 1 0 -21636
box -141 -518 141 518
use sky130_fd_pr__res_xhigh_po_1p41_VXMCTQ  XR36
timestamp 1748944356
transform 0 -1 15953 1 0 -22284
box -141 -512 141 512
use sky130_fd_pr__res_xhigh_po_1p41_9JVM35  XR37
timestamp 1748944356
transform 0 -1 15953 1 0 -22608
box -141 -507 141 507
use sky130_fd_pr__res_xhigh_po_1p41_9JVM35  XR39
timestamp 1748944356
transform 0 -1 15953 1 0 -23256
box -141 -507 141 507
use sky130_fd_pr__res_xhigh_po_1p41_6E4SWG  XR40
timestamp 1748944356
transform 0 -1 15953 1 0 -23580
box -141 -502 141 502
<< end >>
