magic
tech sky130A
magscale 1 2
timestamp 1748941537
<< xpolycontact >>
rect -141 152 141 584
rect -141 -584 141 -152
<< xpolyres >>
rect -141 -152 141 152
<< viali >>
rect -125 169 125 566
rect -125 -566 125 -169
<< metal1 >>
rect -131 566 131 578
rect -131 169 -125 566
rect 125 169 131 566
rect -131 157 131 169
rect -131 -169 131 -157
rect -131 -566 -125 -169
rect 125 -566 131 -169
rect -131 -578 131 -566
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.681 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 2.651k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
