* PEX produced on Thu Jun 12 20:23:40 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from seg_selector_logic.ext - technology: sky130A

.subckt seg_selector_logic_posim b[6] b[7] b[8] b[9] bb[6] bb[7] bb[8] bb[9] S[1] S[2] S[3]
+ S[4] SB[1] SB[2] SB[3] SB[4] VDD GND
X0 x4/x3.B.t0 b[7].t0 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 SB[4].t0 S[4].t3 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2 a_1793_n4793.t1 x3/x3.B.t5 GND.t48 GND.t47 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VDD.t54 b[8].t0 x3/x3.B.t3 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VDD.t73 bb[8].t0 x2/x4.A.t0 VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 x2/x4.A.t1 bb[8].t1 a_781_n5657.t0 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_1497_n4793.t1 b[6].t0 a_1413_n4793.t1 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 x3/x3.B.t4 b[9].t0 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 x2/x5.Y.t1 bb[6].t0 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X9 x2/x5.Y.t2 bb[6].t1 a_1781_n5657.t1 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X10 S[3].t1 x3/x3.B.t6 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 SB[1].t0 S[1].t3 VDD.t44 VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 x1/x3.B.t0 bb[9].t0 a_2253_n4569.t0 GND.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 VDD.t3 bb[9].t1 x1/x3.B.t1 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 x3/x3.B.t0 bb[7].t0 a_1497_n4793.t0 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X15 S[3].t0 x3/x3.A.t5 a_1793_n4793.t0 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 x3/x3.B.t2 b[6].t1 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X17 VDD.t50 bb[9].t2 x2/x4.B.t1 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X18 x2/x4.B.t0 bb[9].t3 a_1057_n5657.t0 GND.t29 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_1057_n5657.t1 b[7].t1 GND.t46 GND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X20 x2/x4.B.t2 b[7].t2 VDD.t58 VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VDD.t19 x4/x3.A.t3 a_1329_n4319.t1 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X22 a_861_n4793.t0 bb[6].t2 a_777_n4793.t0 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 VDD.t13 bb[7].t1 x3/x3.B.t1 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X24 VDD.t71 x3/x3.A.t6 S[3].t2 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 a_777_n4793.t1 b[7].t3 GND.t44 GND.t43 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X26 GND.t19 x4/x3.A.t4 S[4].t2 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 x3/x3.A.t1 b[9].t1 a_945_n4793.t0 GND.t55 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X28 SB[3].t1 S[3].t3 GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X29 VDD.t43 bb[6].t3 x3/x3.A.t2 VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_1329_n4319.t0 x4/x3.B.t3 S[4].t1 VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X31 a_2525_n4319.t1 x1/x3.B.t3 S[1].t1 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X32 a_781_n4569.t0 b[9].t2 GND.t54 GND.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X33 S[4].t0 x4/x3.B.t4 GND.t18 GND.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X34 x1/x3.A.t1 bb[7].t2 a_1977_n4569.t0 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 S[1].t0 x1/x3.B.t4 GND.t22 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 x3/x3.A.t4 b[7].t4 VDD.t56 VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X37 x4/x3.A.t0 b[9].t3 VDD.t68 VDD.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VDD.t11 bb[7].t3 x1/x3.A.t0 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X39 VDD.t35 x1/x3.A.t3 a_2525_n4319.t0 VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X40 a_945_n4793.t1 b[8].t1 a_861_n4793.t1 GND.t38 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X41 VDD.t21 b[6].t2 x2/x4.C.t1 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 x2/x4.C.t2 b[6].t3 a_1333_n5657.t1 GND.t50 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X43 VDD.t66 b[9].t4 x3/x3.A.t0 VDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X44 SB[3].t0 S[3].t4 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X45 S[2].t4 x2/x5.Y.t4 VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X46 a_2065_n5657.t1 x2/x5.Y.t5 GND.t33 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X47 x3/x3.A.t3 b[8].t2 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X48 x1/x3.A.t2 bb[6].t4 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X49 a_1977_n4569.t1 bb[6].t5 GND.t8 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X50 GND.t37 x1/x3.A.t4 S[1].t2 GND.t36 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X51 x2/x4.C.t0 bb[9].t4 VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X52 a_1333_n5657.t0 bb[9].t5 GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X53 a_1781_n5657.t0 bb[7].t4 a_1697_n5657.t0 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X54 VDD.t9 b[8].t3 x4/x3.A.t1 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X55 x4/x3.A.t2 b[8].t4 a_781_n4569.t1 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X56 VDD.t1 bb[7].t5 x2/x5.Y.t0 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X57 x2/x5.Y.t3 b[8].t5 VDD.t52 VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X58 S[2].t1 x2/x4.B.t3 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X59 a_1697_n5657.t1 b[8].t6 GND.t4 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 a_2233_n5657.t0 x2/x4.B.t4 a_2149_n5657.t1 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X61 S[2].t3 x2/x4.A.t3 a_2233_n5657.t1 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X62 VDD.t7 x2/x4.A.t4 S[2].t2 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X63 a_781_n5657.t1 b[9].t5 GND.t52 GND.t51 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X64 a_2149_n5657.t0 x2/x4.C.t3 a_2065_n5657.t0 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X65 x2/x4.A.t2 b[9].t6 VDD.t64 VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X66 VDD.t46 x2/x4.C.t4 S[2].t0 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X67 SB[2].t0 S[2].t5 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X68 SB[2].t1 S[2].t6 GND.t2 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X69 a_1413_n4793.t0 b[8].t7 a_1329_n4793.t1 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X70 VDD.t62 b[6].t4 x4/x3.B.t2 VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X71 x4/x3.B.t1 b[6].t5 a_1057_n4569.t0 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X72 a_1329_n4793.t0 b[9].t7 GND.t56 GND.t17 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X73 x1/x3.B.t2 bb[8].t2 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X74 a_1057_n4569.t1 b[7].t5 GND.t42 GND.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X75 SB[4].t1 S[4].t4 GND.t40 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X76 a_2253_n4569.t1 bb[8].t3 GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X77 SB[1].t1 S[1].t4 GND.t26 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R0 b[7].n3 b[7].t4 231.017
R1 b[7].n0 b[7].t0 229.369
R2 b[7].n6 b[7].t2 229.369
R3 b[7].n3 b[7].t3 158.716
R4 b[7].n0 b[7].t5 157.07
R5 b[7].n6 b[7].t1 157.07
R6 b[7].n1 b[7].n0 152.475
R7 b[7].n4 b[7].n3 152
R8 b[7].n7 b[7].n6 152
R9 b[7].n7 b[7].n5 20.9232
R10 b[7].n2 b[7].n1 17.1938
R11 b[7].n5 b[7].n4 15.9118
R12 b[7].n1 b[7] 5.45235
R13 b[7].n4 b[7] 4.26717
R14 b[7] b[7].n7 2.10199
R15 b[7].n5 b[7].n2 1.30714
R16 b[7].n2 b[7] 0.424328
R17 VDD.n74 VDD.t34 674.802
R18 VDD.t38 VDD.n112 553.428
R19 VDD.n113 VDD 432.123
R20 VDD.n71 VDD.t25 420.43
R21 VDD.t18 VDD 411.372
R22 VDD VDD.t2 366.978
R23 VDD.t61 VDD 366.978
R24 VDD VDD.t10 361.06
R25 VDD.t8 VDD 361.06
R26 VDD.n17 VDD.t66 340.301
R27 VDD.n46 VDD.t13 340.301
R28 VDD.n10 VDD.t7 336.416
R29 VDD.n37 VDD.n35 320.976
R30 VDD.n51 VDD.n19 320.976
R31 VDD.n61 VDD.n16 320.976
R32 VDD.n44 VDD.n23 318.305
R33 VDD VDD.t38 313.707
R34 VDD.n29 VDD.t26 255.905
R35 VDD.n106 VDD.t39 255.905
R36 VDD.n29 VDD.t44 255.904
R37 VDD.n25 VDD.t30 250.722
R38 VDD.n46 VDD.t52 249.52
R39 VDD.n94 VDD.t9 249.363
R40 VDD.n99 VDD.t62 249.363
R41 VDD.n83 VDD.t11 249.363
R42 VDD.n5 VDD.t3 249.363
R43 VDD.n43 VDD.t71 249.362
R44 VDD.n53 VDD.t70 249.062
R45 VDD.n14 VDD.t56 249.062
R46 VDD.n13 VDD.t50 248.929
R47 VDD.t2 VDD.t4 248.599
R48 VDD.t10 VDD.t14 248.599
R49 VDD.t59 VDD.t61 248.599
R50 VDD.t67 VDD.t8 248.599
R51 VDD.n53 VDD.t48 247.394
R52 VDD.n58 VDD.t58 247.394
R53 VDD.n14 VDD.t64 247.394
R54 VDD.n95 VDD.t60 247.394
R55 VDD.n2 VDD.t15 247.394
R56 VDD.n82 VDD.t5 247.394
R57 VDD.n45 VDD.t17 247.394
R58 VDD.n0 VDD.t68 247.393
R59 VDD.n20 VDD.t21 245.178
R60 VDD.n59 VDD.t73 245.178
R61 VDD.n42 VDD.t28 245.178
R62 VDD.n104 VDD.t19 243.512
R63 VDD.n75 VDD.t35 243.512
R64 VDD VDD.n66 230.766
R65 VDD.n112 VDD 219.004
R66 VDD.n69 VDD.n11 213.119
R67 VDD.n67 VDD.n13 213.119
R68 VDD.n68 VDD.n12 213.119
R69 VDD.n112 VDD.n111 213.119
R70 VDD.t34 VDD.t31 213.084
R71 VDD.t24 VDD.t18 213.084
R72 VDD.n70 VDD.n9 209.368
R73 VDD.t4 VDD 207.166
R74 VDD.t14 VDD 207.166
R75 VDD VDD.t59 207.166
R76 VDD VDD.t67 207.166
R77 VDD VDD.t40 206.45
R78 VDD.t31 VDD 189.409
R79 VDD VDD.t24 189.409
R80 VDD.t25 VDD 177.916
R81 VDD.t32 VDD.t45 140.989
R82 VDD.t40 VDD.t16 140.989
R83 VDD.t49 VDD.t57 140.989
R84 VDD.t22 VDD.t20 134.276
R85 VDD.t53 VDD.t47 134.276
R86 VDD.t36 VDD.t72 134.276
R87 VDD.t42 VDD.t63 134.276
R88 VDD VDD.n70 125.883
R89 VDD VDD.n67 124.206
R90 VDD.t27 VDD 107.421
R91 VDD.t51 VDD 107.421
R92 VDD.t69 VDD 107.421
R93 VDD.t55 VDD 107.421
R94 VDD.n69 VDD.t32 100.707
R95 VDD.n68 VDD.t22 100.707
R96 VDD.t0 VDD 97.3503
R97 VDD.n70 VDD.t6 93.9934
R98 VDD.t65 VDD 90.6365
R99 VDD.n67 VDD.t49 80.5659
R100 VDD.t45 VDD.t29 72.1736
R101 VDD VDD.t36 70.4952
R102 VDD.t29 VDD.t27 68.8168
R103 VDD VDD.t12 67.1383
R104 VDD.t6 VDD.n69 60.4245
R105 VDD.t12 VDD.n68 60.4245
R106 VDD VDD.t51 43.6401
R107 VDD.n23 VDD.t41 38.4155
R108 VDD.n28 VDD.n8 34.6358
R109 VDD.n30 VDD.n9 34.6358
R110 VDD.n100 VDD.n88 34.6358
R111 VDD.n107 VDD.n1 34.6358
R112 VDD.n77 VDD.n76 34.6358
R113 VDD.n52 VDD.n51 30.8711
R114 VDD.n62 VDD.n61 30.8711
R115 VDD.n38 VDD.n37 30.8711
R116 VDD.t57 VDD.t65 26.8556
R117 VDD.n19 VDD.t23 26.5955
R118 VDD.n19 VDD.t54 26.5955
R119 VDD.n16 VDD.t37 26.5955
R120 VDD.n16 VDD.t43 26.5955
R121 VDD.n23 VDD.t1 26.5955
R122 VDD.n35 VDD.t33 26.5955
R123 VDD.n35 VDD.t46 26.5955
R124 VDD.n94 VDD.n90 25.977
R125 VDD.n99 VDD.n89 25.977
R126 VDD.n84 VDD.n83 25.977
R127 VDD.n81 VDD.n5 25.977
R128 VDD.n53 VDD.n52 24.4711
R129 VDD.n62 VDD.n14 24.4711
R130 VDD.n90 VDD.n0 24.4711
R131 VDD.n95 VDD.n89 24.4711
R132 VDD.n105 VDD.n104 24.4711
R133 VDD.n84 VDD.n2 24.4711
R134 VDD.n82 VDD.n81 24.4711
R135 VDD.n36 VDD.n11 23.7181
R136 VDD.n71 VDD.n8 23.7181
R137 VDD.n100 VDD.n99 23.7181
R138 VDD.n111 VDD.n1 23.7181
R139 VDD.n77 VDD.n5 23.7181
R140 VDD.n20 VDD.n12 22.5887
R141 VDD.n59 VDD.n58 22.5887
R142 VDD.n43 VDD.n42 22.5887
R143 VDD.n11 VDD.n10 22.5887
R144 VDD.t16 VDD.t0 20.1418
R145 VDD.n104 VDD.n88 19.9534
R146 VDD.n76 VDD.n75 19.9534
R147 VDD.n44 VDD.n43 18.824
R148 VDD.n38 VDD.n25 18.4476
R149 VDD.n41 VDD.n25 16.1887
R150 VDD.n17 VDD.n13 14.3064
R151 VDD.n46 VDD.n45 14.3064
R152 VDD.n45 VDD.n44 14.3064
R153 VDD.n75 VDD.n74 13.5534
R154 VDD.n53 VDD.n13 12.8005
R155 VDD.n58 VDD.n17 12.8005
R156 VDD.n66 VDD.n14 12.8005
R157 VDD.n113 VDD.n0 12.8005
R158 VDD.n95 VDD.n94 12.8005
R159 VDD.n111 VDD.n2 12.8005
R160 VDD.n83 VDD.n82 12.8005
R161 VDD.n46 VDD.n12 12.0476
R162 VDD.n29 VDD.n28 10.5417
R163 VDD.n107 VDD.n106 10.5417
R164 VDD.n74 VDD.n73 9.3005
R165 VDD.n75 VDD.n7 9.3005
R166 VDD.n76 VDD.n6 9.3005
R167 VDD.n78 VDD.n77 9.3005
R168 VDD.n79 VDD.n5 9.3005
R169 VDD.n81 VDD.n80 9.3005
R170 VDD.n82 VDD.n4 9.3005
R171 VDD.n83 VDD.n3 9.3005
R172 VDD.n85 VDD.n84 9.3005
R173 VDD.n86 VDD.n2 9.3005
R174 VDD.n111 VDD.n110 9.3005
R175 VDD.n109 VDD.n1 9.3005
R176 VDD.n108 VDD.n107 9.3005
R177 VDD.n105 VDD.n87 9.3005
R178 VDD.n104 VDD.n103 9.3005
R179 VDD.n102 VDD.n88 9.3005
R180 VDD.n101 VDD.n100 9.3005
R181 VDD.n99 VDD.n98 9.3005
R182 VDD.n97 VDD.n89 9.3005
R183 VDD.n96 VDD.n95 9.3005
R184 VDD.n94 VDD.n93 9.3005
R185 VDD.n92 VDD.n90 9.3005
R186 VDD.n91 VDD.n0 9.3005
R187 VDD.n114 VDD.n113 9.3005
R188 VDD.n66 VDD.n65 9.3005
R189 VDD.n72 VDD.n71 9.3005
R190 VDD.n26 VDD.n8 9.3005
R191 VDD.n28 VDD.n27 9.3005
R192 VDD.n31 VDD.n30 9.3005
R193 VDD.n32 VDD.n9 9.3005
R194 VDD.n33 VDD.n11 9.3005
R195 VDD.n36 VDD.n34 9.3005
R196 VDD.n39 VDD.n38 9.3005
R197 VDD.n41 VDD.n40 9.3005
R198 VDD.n43 VDD.n24 9.3005
R199 VDD.n44 VDD.n22 9.3005
R200 VDD.n45 VDD.n21 9.3005
R201 VDD.n47 VDD.n46 9.3005
R202 VDD.n48 VDD.n12 9.3005
R203 VDD.n50 VDD.n49 9.3005
R204 VDD.n52 VDD.n18 9.3005
R205 VDD.n54 VDD.n53 9.3005
R206 VDD.n55 VDD.n13 9.3005
R207 VDD.n56 VDD.n17 9.3005
R208 VDD.n58 VDD.n57 9.3005
R209 VDD.n60 VDD.n15 9.3005
R210 VDD.n63 VDD.n62 9.3005
R211 VDD.n64 VDD.n14 9.3005
R212 VDD.n30 VDD.n29 8.28285
R213 VDD.n106 VDD.n105 8.28285
R214 VDD.t20 VDD.t53 6.71428
R215 VDD.t47 VDD.t69 6.71428
R216 VDD.t72 VDD.t42 6.71428
R217 VDD.t63 VDD.t55 6.71428
R218 VDD.n73 VDD.n72 6.66136
R219 VDD VDD.n115 3.96214
R220 VDD.n51 VDD.n50 3.76521
R221 VDD.n61 VDD.n60 3.76521
R222 VDD.n37 VDD.n36 3.76521
R223 VDD.n115 VDD 3.09034
R224 VDD.n50 VDD.n20 1.12991
R225 VDD.n60 VDD.n59 1.12991
R226 VDD.n42 VDD.n41 1.12991
R227 VDD.n10 VDD.n9 1.12991
R228 VDD.n7 VDD.n6 0.120292
R229 VDD.n78 VDD.n6 0.120292
R230 VDD.n80 VDD.n79 0.120292
R231 VDD.n80 VDD.n4 0.120292
R232 VDD.n85 VDD.n3 0.120292
R233 VDD.n86 VDD.n85 0.120292
R234 VDD.n109 VDD.n108 0.120292
R235 VDD.n108 VDD.n87 0.120292
R236 VDD.n103 VDD.n102 0.120292
R237 VDD.n102 VDD.n101 0.120292
R238 VDD.n98 VDD.n97 0.120292
R239 VDD.n97 VDD.n96 0.120292
R240 VDD.n93 VDD.n92 0.120292
R241 VDD.n92 VDD.n91 0.120292
R242 VDD.n27 VDD.n26 0.120292
R243 VDD.n31 VDD.n27 0.120292
R244 VDD.n39 VDD.n34 0.120292
R245 VDD.n40 VDD.n39 0.120292
R246 VDD.n24 VDD.n22 0.120292
R247 VDD.n22 VDD.n21 0.120292
R248 VDD.n49 VDD.n18 0.120292
R249 VDD.n54 VDD.n18 0.120292
R250 VDD.n57 VDD.n56 0.120292
R251 VDD.n63 VDD.n15 0.120292
R252 VDD.n64 VDD.n63 0.120292
R253 VDD VDD.n7 0.0603958
R254 VDD.n79 VDD 0.0603958
R255 VDD VDD.n3 0.0603958
R256 VDD.n110 VDD 0.0603958
R257 VDD VDD.n109 0.0603958
R258 VDD.n103 VDD 0.0603958
R259 VDD.n98 VDD 0.0603958
R260 VDD.n93 VDD 0.0603958
R261 VDD.n114 VDD 0.0603958
R262 VDD.n26 VDD 0.0603958
R263 VDD.n32 VDD 0.0603958
R264 VDD.n33 VDD 0.0603958
R265 VDD.n34 VDD 0.0603958
R266 VDD VDD.n24 0.0603958
R267 VDD.n47 VDD 0.0603958
R268 VDD.n48 VDD 0.0603958
R269 VDD.n49 VDD 0.0603958
R270 VDD.n55 VDD 0.0603958
R271 VDD.n56 VDD 0.0603958
R272 VDD VDD.n15 0.0603958
R273 VDD.n65 VDD 0.0603958
R274 VDD.n110 VDD 0.0382604
R275 VDD.n115 VDD 0.0365577
R276 VDD.n73 VDD 0.03175
R277 VDD VDD.n114 0.03175
R278 VDD.n72 VDD 0.03175
R279 VDD VDD.n32 0.03175
R280 VDD VDD.n33 0.03175
R281 VDD VDD.n48 0.03175
R282 VDD VDD.n55 0.03175
R283 VDD.n65 VDD 0.03175
R284 VDD.n4 VDD 0.0239375
R285 VDD VDD.n86 0.0239375
R286 VDD.n96 VDD 0.0239375
R287 VDD.n91 VDD 0.0239375
R288 VDD.n21 VDD 0.0239375
R289 VDD.n57 VDD 0.0239375
R290 VDD VDD.n87 0.0226354
R291 VDD VDD.n31 0.0226354
R292 VDD VDD.n78 0.0213333
R293 VDD.n101 VDD 0.0213333
R294 VDD.n40 VDD 0.0213333
R295 VDD VDD.n47 0.0213333
R296 VDD VDD.n54 0.0213333
R297 VDD VDD.n64 0.0213333
R298 x4/x3.B.n0 x4/x3.B.t3 230.363
R299 x4/x3.B.n3 x4/x3.B.n2 201.161
R300 x4/x3.B.n0 x4/x3.B.t4 158.064
R301 x4/x3.B.n1 x4/x3.B.n0 155.328
R302 x4/x3.B.n4 x4/x3.B.t1 140.53
R303 x4/x3.B x4/x3.B.n3 36.416
R304 x4/x3.B.n3 x4/x3.B.n1 29.1319
R305 x4/x3.B.n2 x4/x3.B.t2 26.5955
R306 x4/x3.B.n2 x4/x3.B.t0 26.5955
R307 x4/x3.B.n4 x4/x3.B 16.5652
R308 x4/x3.B x4/x3.B.n4 9.03579
R309 x4/x3.B.n1 x4/x3.B 3.0725
R310 x4/x3.B.n4 x4/x3.B 1.72748
R311 S[4].n1 S[4] 593.34
R312 S[4].n2 S[4].n1 289.24
R313 S[4].n4 S[4].t3 230.576
R314 S[4].n4 S[4].t4 158.275
R315 S[4].n5 S[4].n4 152
R316 S[4].n3 S[4].n0 147.262
R317 S[4].n3 S[4].n2 29.5774
R318 S[4].n1 S[4].t1 26.5955
R319 S[4].n0 S[4].t2 24.9236
R320 S[4].n0 S[4].t0 24.9236
R321 S[4].n2 S[4] 11.3699
R322 S[4].n5 S[4] 11.2025
R323 S[4] S[4].n3 9.78711
R324 S[4] S[4].n5 6.66717
R325 SB[4].n0 SB[4].t0 235.56
R326 SB[4] SB[4].t1 152.889
R327 SB[4] SB[4].n0 2.22659
R328 SB[4].n0 SB[4] 1.55202
R329 x3/x3.B.n2 x3/x3.B.n1 258.363
R330 x3/x3.B.n6 x3/x3.B.t0 257
R331 x3/x3.B.n6 x3/x3.B.t0 249
R332 x3/x3.B.n3 x3/x3.B.t6 229.369
R333 x3/x3.B.n2 x3/x3.B.n0 202.094
R334 x3/x3.B.n3 x3/x3.B.t5 157.07
R335 x3/x3.B.n4 x3/x3.B.n3 152
R336 x3/x3.B.n7 x3/x3.B.n5 61.3652
R337 x3/x3.B.n0 x3/x3.B.t1 32.5055
R338 x3/x3.B.n0 x3/x3.B.t2 32.5055
R339 x3/x3.B.n1 x3/x3.B.t3 26.5955
R340 x3/x3.B.n1 x3/x3.B.t4 26.5955
R341 x3/x3.B.n5 x3/x3.B.n4 19.8407
R342 x3/x3.B.n7 x3/x3.B.n6 6.51278
R343 x3/x3.B.n4 x3/x3.B 5.92643
R344 x3/x3.B x3/x3.B.n7 4.04261
R345 x3/x3.B.n5 x3/x3.B.n2 1.12991
R346 GND.n110 GND.n1 1.01257e+06
R347 GND.n13 GND.n1 7616.32
R348 GND.n110 GND.n109 7503.85
R349 GND.n13 GND.t1 2662.78
R350 GND.n7 GND.t50 1993.53
R351 GND GND.t14 1865.37
R352 GND GND.t31 1765.7
R353 GND GND.t29 1737.22
R354 GND GND.t12 1737.22
R355 GND.t1 GND 1509.39
R356 GND.t14 GND.t16 1366.99
R357 GND.t31 GND.t23 1366.99
R358 GND.n68 GND.t36 1213.79
R359 GND.n30 GND.n25 1198.25
R360 GND.n43 GND.n31 1198.25
R361 GND.n29 GND.n16 1198.25
R362 GND.n67 GND.n66 1198.25
R363 GND.n109 GND.n108 1198.25
R364 GND.n92 GND.n7 1198.25
R365 GND.n14 GND.n13 1198.25
R366 GND.t16 GND.t24 1196.12
R367 GND.t24 GND.t32 1196.12
R368 GND.t23 GND.t3 1196.12
R369 GND.t50 GND.t34 1196.12
R370 GND.t29 GND.t45 1196.12
R371 GND.t12 GND.t51 1196.12
R372 GND GND.n7 1082.2
R373 GND.n109 GND 1053.72
R374 GND.t34 GND 996.764
R375 GND.t45 GND 996.764
R376 GND.t51 GND 996.764
R377 GND.t32 GND 911.327
R378 GND.t3 GND 911.327
R379 GND.n68 GND.n1 708.047
R380 GND.t5 GND.t20 708.047
R381 GND.t17 GND.t5 708.047
R382 GND.t49 GND.t41 708.047
R383 GND.n111 GND.n110 708.047
R384 GND.t38 GND.t15 674.331
R385 GND.t9 GND.t53 674.331
R386 GND.t27 GND 649.043
R387 GND.t39 GND 649.043
R388 GND.n31 GND 640.614
R389 GND GND.n67 632.184
R390 GND.n111 GND 623.755
R391 GND.n69 GND.n68 599.125
R392 GND.n112 GND.n111 599.125
R393 GND GND.t10 590.038
R394 GND GND.t7 590.038
R395 GND GND.t47 590.038
R396 GND.t21 GND 539.465
R397 GND GND.t17 539.465
R398 GND.t43 GND 539.465
R399 GND GND.t30 514.177
R400 GND.t55 GND 455.173
R401 GND.t0 GND.t39 446.743
R402 GND GND.t0 446.743
R403 GND.n67 GND.t13 404.599
R404 GND.n31 GND.t49 404.599
R405 GND.t30 GND.t27 379.31
R406 GND.n29 GND.t13 370.882
R407 GND.n30 GND.t6 370.882
R408 GND.t36 GND.t25 362.452
R409 GND.t20 GND 362.452
R410 GND GND.t38 354.024
R411 GND.t25 GND.t21 345.594
R412 GND.t10 GND.n29 337.166
R413 GND.t47 GND.n30 337.166
R414 GND.n6 GND.t4 274.812
R415 GND.t6 GND 252.875
R416 GND.t7 GND 193.87
R417 GND.n75 GND.t2 158.361
R418 GND.n26 GND.t40 158.361
R419 GND.n24 GND.t28 158.361
R420 GND.n44 GND.t18 155.63
R421 GND.n48 GND.t19 154.131
R422 GND.n15 GND.t37 154.131
R423 GND.n21 GND.t26 153.631
R424 GND.n17 GND.t22 152.381
R425 GND.n97 GND.t35 150.922
R426 GND.n102 GND.t46 150.922
R427 GND.n2 GND.t52 150.922
R428 GND.n53 GND.t48 150.922
R429 GND.n57 GND.t8 150.922
R430 GND.n62 GND.t11 150.922
R431 GND.n39 GND.t42 150.922
R432 GND.n44 GND.t56 149.493
R433 GND.n9 GND.t33 149.493
R434 GND.n32 GND.t54 147.411
R435 GND.n33 GND.t44 146.245
R436 GND.t41 GND.t55 134.867
R437 GND.n87 GND.n86 34.6358
R438 GND.n88 GND.n87 34.6358
R439 GND.n76 GND.n11 34.6358
R440 GND.n80 GND.n11 34.6358
R441 GND.n81 GND.n80 34.6358
R442 GND.n82 GND.n81 34.6358
R443 GND.n74 GND.n73 34.6358
R444 GND.n93 GND.n5 34.6358
R445 GND.n98 GND.n4 34.6358
R446 GND.n104 GND.n103 34.6358
R447 GND.n38 GND.n34 34.6358
R448 GND.t15 GND.t9 33.717
R449 GND.t53 GND.t43 33.717
R450 GND.n34 GND.n33 32.7534
R451 GND.n88 GND.n6 25.977
R452 GND.n48 GND.n27 24.4711
R453 GND.n49 GND.n48 24.4711
R454 GND.n20 GND.n15 24.4711
R455 GND.n86 GND.n9 24.0946
R456 GND.n112 GND.n0 23.7181
R457 GND.n73 GND.n14 23.7181
R458 GND.n93 GND.n92 23.7181
R459 GND.n98 GND.n97 23.7181
R460 GND.n103 GND.n102 23.7181
R461 GND.n53 GND.n52 23.7181
R462 GND.n62 GND.n61 23.7181
R463 GND.n43 GND.n28 23.7181
R464 GND.n39 GND.n38 23.7181
R465 GND.n66 GND.n17 23.3417
R466 GND.n97 GND.n5 22.2123
R467 GND.n102 GND.n4 22.2123
R468 GND.n104 GND.n2 22.2123
R469 GND.n58 GND.n57 22.2123
R470 GND.n39 GND.n28 22.2123
R471 GND.n82 GND.n9 19.9534
R472 GND.n44 GND.n27 19.9534
R473 GND.n21 GND.n20 19.2005
R474 GND.n22 GND.n21 15.4358
R475 GND.n69 GND.n15 13.5534
R476 GND.n92 GND.n6 13.177
R477 GND.n44 GND.n43 13.177
R478 GND.n108 GND.n2 12.8005
R479 GND.n57 GND.n25 12.8005
R480 GND.n66 GND.n16 12.8005
R481 GND.n53 GND.n25 11.2946
R482 GND.n62 GND.n16 11.2946
R483 GND.n75 GND.n74 10.5417
R484 GND.n52 GND.n26 10.5417
R485 GND.n61 GND.n24 10.5417
R486 GND.n113 GND.n112 9.3005
R487 GND.n70 GND.n69 9.3005
R488 GND.n18 GND.n15 9.3005
R489 GND.n20 GND.n19 9.3005
R490 GND.n23 GND.n22 9.3005
R491 GND.n66 GND.n65 9.3005
R492 GND.n64 GND.n16 9.3005
R493 GND.n63 GND.n62 9.3005
R494 GND.n61 GND.n60 9.3005
R495 GND.n59 GND.n58 9.3005
R496 GND.n57 GND.n56 9.3005
R497 GND.n55 GND.n25 9.3005
R498 GND.n54 GND.n53 9.3005
R499 GND.n52 GND.n51 9.3005
R500 GND.n50 GND.n49 9.3005
R501 GND.n48 GND.n47 9.3005
R502 GND.n46 GND.n27 9.3005
R503 GND.n45 GND.n44 9.3005
R504 GND.n43 GND.n42 9.3005
R505 GND.n41 GND.n28 9.3005
R506 GND.n40 GND.n39 9.3005
R507 GND.n38 GND.n37 9.3005
R508 GND.n36 GND.n34 9.3005
R509 GND.n35 GND.n0 9.3005
R510 GND.n108 GND.n107 9.3005
R511 GND.n71 GND.n14 9.3005
R512 GND.n73 GND.n72 9.3005
R513 GND.n74 GND.n12 9.3005
R514 GND.n77 GND.n76 9.3005
R515 GND.n78 GND.n11 9.3005
R516 GND.n80 GND.n79 9.3005
R517 GND.n81 GND.n10 9.3005
R518 GND.n83 GND.n82 9.3005
R519 GND.n84 GND.n9 9.3005
R520 GND.n86 GND.n85 9.3005
R521 GND.n87 GND.n8 9.3005
R522 GND.n89 GND.n88 9.3005
R523 GND.n90 GND.n6 9.3005
R524 GND.n92 GND.n91 9.3005
R525 GND.n94 GND.n93 9.3005
R526 GND.n95 GND.n5 9.3005
R527 GND.n97 GND.n96 9.3005
R528 GND.n99 GND.n98 9.3005
R529 GND.n100 GND.n4 9.3005
R530 GND.n102 GND.n101 9.3005
R531 GND.n103 GND.n3 9.3005
R532 GND.n105 GND.n104 9.3005
R533 GND.n106 GND.n2 9.3005
R534 GND.n71 GND.n70 7.14052
R535 GND.n76 GND.n75 6.77697
R536 GND.n49 GND.n26 6.77697
R537 GND.n58 GND.n24 6.77697
R538 GND GND.n114 3.72256
R539 GND.n114 GND 2.85076
R540 GND.n33 GND.n32 1.12991
R541 GND.n32 GND.n0 0.753441
R542 GND.n114 GND 0.473256
R543 GND.n22 GND.n17 0.376971
R544 GND.n19 GND.n18 0.120292
R545 GND.n23 GND.n19 0.120292
R546 GND.n60 GND.n59 0.120292
R547 GND.n51 GND.n50 0.120292
R548 GND.n47 GND.n46 0.120292
R549 GND.n46 GND.n45 0.120292
R550 GND.n41 GND.n40 0.120292
R551 GND.n37 GND.n36 0.120292
R552 GND.n36 GND.n35 0.120292
R553 GND.n72 GND.n12 0.120292
R554 GND.n77 GND.n12 0.120292
R555 GND.n79 GND.n78 0.120292
R556 GND.n79 GND.n10 0.120292
R557 GND.n83 GND.n10 0.120292
R558 GND.n84 GND.n83 0.120292
R559 GND.n85 GND.n8 0.120292
R560 GND.n89 GND.n8 0.120292
R561 GND.n90 GND.n89 0.120292
R562 GND.n95 GND.n94 0.120292
R563 GND.n96 GND.n95 0.120292
R564 GND.n100 GND.n99 0.120292
R565 GND.n101 GND.n100 0.120292
R566 GND.n105 GND.n3 0.120292
R567 GND.n106 GND.n105 0.120292
R568 GND.n18 GND 0.0603958
R569 GND.n65 GND 0.0603958
R570 GND GND.n64 0.0603958
R571 GND GND.n63 0.0603958
R572 GND.n60 GND 0.0603958
R573 GND.n56 GND 0.0603958
R574 GND GND.n55 0.0603958
R575 GND GND.n54 0.0603958
R576 GND.n51 GND 0.0603958
R577 GND.n47 GND 0.0603958
R578 GND.n42 GND 0.0603958
R579 GND GND.n41 0.0603958
R580 GND.n37 GND 0.0603958
R581 GND.n113 GND 0.0603958
R582 GND.n72 GND 0.0603958
R583 GND.n78 GND 0.0603958
R584 GND.n85 GND 0.0603958
R585 GND.n91 GND 0.0603958
R586 GND.n94 GND 0.0603958
R587 GND.n99 GND 0.0603958
R588 GND GND.n3 0.0603958
R589 GND.n107 GND 0.0603958
R590 GND.n55 GND 0.0343542
R591 GND.n70 GND 0.0330521
R592 GND.n65 GND 0.0330521
R593 GND.n64 GND 0.0330521
R594 GND.n42 GND 0.0330521
R595 GND GND.n113 0.0330521
R596 GND GND.n71 0.0330521
R597 GND.n91 GND 0.0330521
R598 GND.n107 GND 0.0330521
R599 GND.n63 GND 0.0239375
R600 GND.n56 GND 0.0239375
R601 GND.n54 GND 0.0239375
R602 GND.n40 GND 0.0239375
R603 GND.n96 GND 0.0239375
R604 GND.n101 GND 0.0239375
R605 GND GND.n106 0.0239375
R606 GND.n59 GND 0.0226354
R607 GND.n50 GND 0.0226354
R608 GND GND.n77 0.0226354
R609 GND GND.n23 0.0213333
R610 GND.n45 GND 0.0213333
R611 GND.n35 GND 0.0213333
R612 GND GND.n84 0.0213333
R613 GND GND.n90 0.0213333
R614 a_1793_n4793.t0 a_1793_n4793.t1 49.8467
R615 b[8].n5 b[8].t2 241.536
R616 b[8].n3 b[8].t0 241.536
R617 b[8].n8 b[8].t5 230.363
R618 b[8].n0 b[8].t3 230.155
R619 b[8] b[8].n5 177.839
R620 b[8].n5 b[8].t1 169.237
R621 b[8].n3 b[8].t7 169.237
R622 b[8].n4 b[8].n3 159.37
R623 b[8].n8 b[8].t6 158.064
R624 b[8].n0 b[8].t4 157.856
R625 b[8].n1 b[8].n0 152
R626 b[8].n9 b[8].n8 152
R627 b[8].n6 b[8].n4 40.9264
R628 b[8].n9 b[8].n7 35.3808
R629 b[8].n2 b[8].n1 17.557
R630 b[8].n6 b[8] 12.9576
R631 b[8].n7 b[8].n6 6.5302
R632 b[8].n4 b[8] 3.49141
R633 b[8] b[8].n9 3.2005
R634 b[8].n1 b[8] 2.10199
R635 b[8].n7 b[8].n2 0.852062
R636 b[8].n2 b[8] 0.533703
R637 bb[8].n3 bb[8].t0 230.155
R638 bb[8].n0 bb[8].t2 229.369
R639 bb[8].n3 bb[8].t1 157.856
R640 bb[8].n0 bb[8].t3 157.07
R641 bb[8].n1 bb[8].n0 152
R642 bb[8].n4 bb[8].n3 152
R643 bb[8].n4 bb[8].n2 38.4791
R644 bb[8].n2 bb[8].n1 20.0252
R645 bb[8].n1 bb[8] 5.92643
R646 bb[8] bb[8].n4 2.10199
R647 bb[8].n2 bb[8] 0.619641
R648 x2/x4.A x2/x4.A.n3 237.577
R649 x2/x4.A.n0 x2/x4.A.t4 228.649
R650 x2/x4.A.n0 x2/x4.A.t3 156.35
R651 x2/x4.A.n1 x2/x4.A.n0 152
R652 x2/x4.A.n2 x2/x4.A.t1 131.691
R653 x2/x4.A.n2 x2/x4.A.n1 35.0201
R654 x2/x4.A.n3 x2/x4.A.t0 26.5955
R655 x2/x4.A.n3 x2/x4.A.t2 26.5955
R656 x2/x4.A.n4 x2/x4.A 16.5652
R657 x2/x4.A x2/x4.A.n4 9.03579
R658 x2/x4.A.n4 x2/x4.A.n2 8.8386
R659 x2/x4.A.n4 x2/x4.A 1.72748
R660 x2/x4.A.n1 x2/x4.A 1.43334
R661 a_781_n5657.t0 a_781_n5657.t1 49.8467
R662 b[6].n3 b[6].t1 241.536
R663 b[6].n0 b[6].t4 230.155
R664 b[6].n5 b[6].t2 230.155
R665 b[6] b[6].n3 177.839
R666 b[6].n3 b[6].t0 169.237
R667 b[6].n0 b[6].t5 157.856
R668 b[6].n5 b[6].t3 157.856
R669 b[6].n1 b[6].n0 152
R670 b[6].n6 b[6].n5 152
R671 b[6].n6 b[6].n4 23.3603
R672 b[6].n4 b[6] 22.9626
R673 b[6].n2 b[6].n1 19.8793
R674 b[6].n1 b[6] 2.10199
R675 b[6] b[6].n6 2.10199
R676 b[6].n4 b[6].n2 1.23683
R677 b[6].n2 b[6] 0.314953
R678 a_1413_n4793.t0 a_1413_n4793.t1 49.8467
R679 a_1497_n4793.t0 a_1497_n4793.t1 60.9236
R680 b[9].n0 b[9].t0 231.017
R681 b[9].n2 b[9].t3 229.369
R682 b[9].n5 b[9].t6 229.369
R683 b[9].n1 b[9].t4 228.649
R684 b[9].n0 b[9].t7 158.716
R685 b[9].n2 b[9].t2 157.07
R686 b[9].n5 b[9].t5 157.07
R687 b[9].n1 b[9].t1 156.35
R688 b[9] b[9].n0 156.268
R689 b[9].n3 b[9].n2 153.423
R690 b[9].n6 b[9].n5 152
R691 b[9].n8 b[9].n1 152
R692 b[9].n8 b[9] 53.8309
R693 b[9].n7 b[9].n6 19.5676
R694 b[9].n8 b[9].n7 16.4183
R695 b[9].n4 b[9].n3 14.4998
R696 b[9].n6 b[9] 5.92643
R697 b[9].n3 b[9] 4.5042
R698 b[9] b[9].n8 1.43334
R699 b[9].n7 b[9].n4 1.10597
R700 b[9].n4 b[9] 0.725109
R701 bb[6].n2 bb[6].t3 241.536
R702 bb[6].n0 bb[6].t0 232.214
R703 bb[6].n6 bb[6].t4 229.369
R704 bb[6].n2 bb[6].t2 169.237
R705 bb[6].n0 bb[6].t1 159.915
R706 bb[6].n6 bb[6].t5 157.07
R707 bb[6].n3 bb[6].n2 155.88
R708 bb[6].n1 bb[6].n0 152
R709 bb[6].n7 bb[6].n6 152
R710 bb[6].n4 bb[6].n3 23.417
R711 bb[6].n4 bb[6].n1 22.0085
R712 bb[6].n7 bb[6].n5 18.2158
R713 bb[6].n3 bb[6] 6.98232
R714 bb[6] bb[6].n7 5.92643
R715 bb[6].n1 bb[6] 2.27147
R716 bb[6].n5 bb[6].n4 1.42823
R717 bb[6].n5 bb[6] 0.580578
R718 x2/x5.Y.n4 x2/x5.Y.t1 274.793
R719 x2/x5.Y.n0 x2/x5.Y.t4 231.017
R720 x2/x5.Y.n4 x2/x5.Y.n3 205.28
R721 x2/x5.Y.n0 x2/x5.Y.t5 158.716
R722 x2/x5.Y.n1 x2/x5.Y.n0 152.583
R723 x2/x5.Y.n2 x2/x5.Y.t2 130.49
R724 x2/x5.Y x2/x5.Y.n4 67.4857
R725 x2/x5.Y x2/x5.Y.n2 38.9629
R726 x2/x5.Y.n3 x2/x5.Y.t0 26.5955
R727 x2/x5.Y.n3 x2/x5.Y.t3 26.5955
R728 x2/x5.Y.n2 x2/x5.Y.n1 22.1046
R729 x2/x5.Y.n1 x2/x5.Y 3.68535
R730 a_1781_n5657.t0 a_1781_n5657.t1 60.9236
R731 S[3].n0 S[3].t4 230.576
R732 S[3] S[3].n2 224.778
R733 S[3].n3 S[3] 217.601
R734 S[3].n0 S[3].t3 158.275
R735 S[3].n6 S[3].n0 152.8
R736 S[3].n1 S[3].t0 132.067
R737 S[3].n4 S[3].n3 64.0005
R738 S[3].n2 S[3].t2 26.5955
R739 S[3].n2 S[3].t1 26.5955
R740 S[3].n6 S[3] 9.9183
R741 S[3] S[3].n5 9.79142
R742 S[3] S[3].n6 5.86717
R743 S[3].n3 S[3] 3.38874
R744 S[3].n5 S[3].n1 2.6841
R745 S[3].n5 S[3].n4 1.47388
R746 S[3].n1 S[3] 1.17559
R747 S[3].n4 S[3] 0.921363
R748 S[1].n0 S[1].t3 230.576
R749 S[1].n1 S[1].t1 218.572
R750 S[1].n0 S[1].t4 158.275
R751 S[1].n4 S[1].n0 152
R752 S[1].n3 S[1].n2 94.1864
R753 S[1].n3 S[1].n1 86.3316
R754 S[1].n2 S[1].t2 24.9236
R755 S[1].n2 S[1].t0 24.9236
R756 S[1] S[1].n3 16.7298
R757 S[1].n4 S[1] 13.9107
R758 S[1].n1 S[1] 7.54721
R759 S[1] S[1].n4 6.66717
R760 SB[1] SB[1].t0 230.518
R761 SB[1] SB[1].t1 162.351
R762 SB[1].n0 SB[1] 10.5744
R763 SB[1] SB[1].n0 7.23528
R764 SB[1].n0 SB[1] 5.04292
R765 bb[9].n1 bb[9].t1 230.155
R766 bb[9].n5 bb[9].t2 230.155
R767 bb[9].n0 bb[9].t4 229.369
R768 bb[9] bb[9].n0 157.927
R769 bb[9].n1 bb[9].t0 157.856
R770 bb[9].n5 bb[9].t3 157.856
R771 bb[9].n0 bb[9].t5 157.07
R772 bb[9].n2 bb[9].n1 152
R773 bb[9].n6 bb[9].n5 152
R774 bb[9].n4 bb[9].n3 33.573
R775 bb[9].n3 bb[9].n2 19.1764
R776 bb[9].n4 bb[9] 11.0938
R777 bb[9].n6 bb[9].n4 9.9845
R778 bb[9] bb[9].n6 2.3045
R779 bb[9].n2 bb[9] 2.10199
R780 bb[9].n3 bb[9] 0.729016
R781 a_2253_n4569.t0 a_2253_n4569.t1 49.8467
R782 x1/x3.B.n1 x1/x3.B.t0 268.077
R783 x1/x3.B.n1 x1/x3.B.t0 258.846
R784 x1/x3.B x1/x3.B.n0 237.577
R785 x1/x3.B.n2 x1/x3.B.t3 230.363
R786 x1/x3.B.n2 x1/x3.B.t4 158.064
R787 x1/x3.B.n3 x1/x3.B.n2 153.28
R788 x1/x3.B.n0 x1/x3.B.t1 26.5955
R789 x1/x3.B.n0 x1/x3.B.t2 26.5955
R790 x1/x3.B.n4 x1/x3.B.n3 19.4367
R791 x1/x3.B.n5 x1/x3.B 16.5652
R792 x1/x3.B.n5 x1/x3.B 9.03579
R793 x1/x3.B.n5 x1/x3.B.n4 7.72113
R794 x1/x3.B.n3 x1/x3.B 5.1205
R795 x1/x3.B x1/x3.B.n5 1.72748
R796 x1/x3.B.n4 x1/x3.B.n1 1.11796
R797 bb[7].n6 bb[7].t5 241.536
R798 bb[7].n0 bb[7].t3 230.155
R799 bb[7].n3 bb[7].t1 228.649
R800 bb[7].n6 bb[7].t4 169.237
R801 bb[7].n0 bb[7].t2 157.856
R802 bb[7].n3 bb[7].t0 156.35
R803 bb[7] bb[7].n6 154.744
R804 bb[7].n1 bb[7].n0 152
R805 bb[7].n4 bb[7].n3 152
R806 bb[7].n5 bb[7].n4 24.2462
R807 bb[7] bb[7].n5 20.7968
R808 bb[7].n2 bb[7].n1 19.5604
R809 bb[7].n4 bb[7] 6.13383
R810 bb[7].n1 bb[7] 2.10199
R811 bb[7].n5 bb[7].n2 1.1548
R812 bb[7].n2 bb[7] 0.314953
R813 x3/x3.A.n5 x3/x3.A.n0 258.363
R814 x3/x3.A.n1 x3/x3.A.t6 230.155
R815 x3/x3.A.n4 x3/x3.A.n3 196.889
R816 x3/x3.A.n1 x3/x3.A.t5 157.856
R817 x3/x3.A.n2 x3/x3.A.n1 152
R818 x3/x3.A.n6 x3/x3.A.t1 132.982
R819 x3/x3.A.n6 x3/x3.A.n5 62.4946
R820 x3/x3.A.n3 x3/x3.A.t0 32.5055
R821 x3/x3.A.n3 x3/x3.A.t3 32.5055
R822 x3/x3.A.n4 x3/x3.A.n2 30.2423
R823 x3/x3.A.n0 x3/x3.A.t2 26.5955
R824 x3/x3.A.n0 x3/x3.A.t4 26.5955
R825 x3/x3.A.n5 x3/x3.A.n4 5.2056
R826 x3/x3.A x3/x3.A.n6 4.04261
R827 x3/x3.A.n2 x3/x3.A 2.3045
R828 x2/x4.B.n3 x2/x4.B.t0 268.077
R829 x2/x4.B.n3 x2/x4.B.t0 258.846
R830 x2/x4.B.n1 x2/x4.B.t3 241.536
R831 x2/x4.B x2/x4.B.n0 237.577
R832 x2/x4.B.n1 x2/x4.B.t4 169.237
R833 x2/x4.B.n2 x2/x4.B.n1 153.032
R834 x2/x4.B.n3 x2/x4.B.n2 32.8186
R835 x2/x4.B.n2 x2/x4.B 31.0244
R836 x2/x4.B.n0 x2/x4.B.t1 26.5955
R837 x2/x4.B.n0 x2/x4.B.t2 26.5955
R838 x2/x4.B.n4 x2/x4.B 16.5652
R839 x2/x4.B.n4 x2/x4.B 9.03579
R840 x2/x4.B.n4 x2/x4.B.n3 8.8386
R841 x2/x4.B x2/x4.B.n4 1.72748
R842 a_1057_n5657.t0 a_1057_n5657.t1 49.8467
R843 x4/x3.A x4/x3.A.n3 237.577
R844 x4/x3.A.n0 x4/x3.A.t3 231.835
R845 x4/x3.A.n0 x4/x3.A.t4 157.07
R846 x4/x3.A.n1 x4/x3.A.n0 152
R847 x4/x3.A.n2 x4/x3.A.t2 132.505
R848 x4/x3.A.n3 x4/x3.A.t1 26.5955
R849 x4/x3.A.n3 x4/x3.A.t0 26.5955
R850 x4/x3.A.n2 x4/x3.A.n1 22.6473
R851 x4/x3.A.n4 x4/x3.A 16.5652
R852 x4/x3.A x4/x3.A.n4 9.03579
R853 x4/x3.A.n4 x4/x3.A.n2 8.0259
R854 x4/x3.A.n1 x4/x3.A 2.01193
R855 x4/x3.A.n4 x4/x3.A 1.72748
R856 a_1329_n4319.t0 a_1329_n4319.t1 41.3705
R857 a_777_n4793.t0 a_777_n4793.t1 49.8467
R858 a_861_n4793.t0 a_861_n4793.t1 49.8467
R859 a_945_n4793.t0 a_945_n4793.t1 60.9236
R860 SB[3] SB[3].t0 230.518
R861 SB[3] SB[3].t1 148.715
R862 SB[3].n0 SB[3] 11.6875
R863 SB[3] SB[3].n0 7.23528
R864 SB[3].n0 SB[3] 5.04292
R865 a_2525_n4319.t0 a_2525_n4319.t1 41.3705
R866 a_781_n4569.t0 a_781_n4569.t1 49.8467
R867 a_1977_n4569.t0 a_1977_n4569.t1 49.8467
R868 x1/x3.A x1/x3.A.n0 237.577
R869 x1/x3.A.n2 x1/x3.A.t3 231.835
R870 x1/x3.A.n2 x1/x3.A.t4 157.07
R871 x1/x3.A x1/x3.A.n2 154.304
R872 x1/x3.A.n1 x1/x3.A.t1 140.53
R873 x1/x3.A.n3 x1/x3.A 32.1479
R874 x1/x3.A.n0 x1/x3.A.t0 26.5955
R875 x1/x3.A.n0 x1/x3.A.t2 26.5955
R876 x1/x3.A x1/x3.A.n3 14.3064
R877 x1/x3.A.n1 x1/x3.A 9.03579
R878 x1/x3.A.n3 x1/x3.A.n1 2.25932
R879 x1/x3.A.n1 x1/x3.A 1.72748
R880 x2/x4.C.n1 x2/x4.C.t4 241.536
R881 x2/x4.C.n3 x2/x4.C.n0 227.412
R882 x2/x4.C.n1 x2/x4.C.t3 169.237
R883 x2/x4.C.n2 x2/x4.C.n1 155.103
R884 x2/x4.C.n4 x2/x4.C.t2 140.53
R885 x2/x4.C.n3 x2/x4.C.n2 30.9223
R886 x2/x4.C.n0 x2/x4.C.t1 26.5955
R887 x2/x4.C.n0 x2/x4.C.t0 26.5955
R888 x2/x4.C x2/x4.C.n4 16.5652
R889 x2/x4.C x2/x4.C.n3 10.1652
R890 x2/x4.C.n4 x2/x4.C 9.03579
R891 x2/x4.C.n2 x2/x4.C 7.75808
R892 x2/x4.C.n4 x2/x4.C 1.72748
R893 a_1333_n5657.t0 a_1333_n5657.t1 49.8467
R894 S[2].n2 S[2].n1 258.363
R895 S[2].n3 S[2].t5 230.576
R896 S[2].n2 S[2].n0 202.095
R897 S[2].n3 S[2].t6 158.275
R898 S[2].n4 S[2].n3 152
R899 S[2].n6 S[2].t3 126.469
R900 S[2].n7 S[2].n2 62.4946
R901 S[2].n0 S[2].t2 32.5055
R902 S[2].n0 S[2].t1 32.5055
R903 S[2].n1 S[2].t0 26.5955
R904 S[2].n1 S[2].t4 26.5955
R905 S[2].n5 S[2].n4 11.7269
R906 S[2].n6 S[2].n5 10.2876
R907 S[2].n4 S[2] 6.66717
R908 S[2].n7 S[2].n6 6.51278
R909 S[2] S[2].n7 4.04261
R910 S[2].n5 S[2] 0.0496071
R911 a_2065_n5657.t0 a_2065_n5657.t1 49.8467
R912 a_1697_n5657.t0 a_1697_n5657.t1 49.8467
R913 a_2149_n5657.t0 a_2149_n5657.t1 49.8467
R914 a_2233_n5657.t0 a_2233_n5657.t1 60.9236
R915 SB[2].n0 SB[2].t0 235.56
R916 SB[2] SB[2].t1 162.351
R917 SB[2] SB[2].n0 2.22659
R918 SB[2].n0 SB[2] 1.55202
R919 a_1329_n4793.t0 a_1329_n4793.t1 49.8467
R920 a_1057_n4569.t0 a_1057_n4569.t1 49.8467
C0 bb[7] SB[2] 0.02239f
C1 bb[6] b[8] 0.19889f
C2 bb[6] S[1] 0.10327f
C3 b[6] x2/x4.A 0.02251f
C4 VDD bb[9] 1.50788f
C5 bb[6] x3/x3.A 0.63473f
C6 b[8] x2/x5.Y 0.10245f
C7 b[6] b[9] 0.19231f
C8 bb[6] x1/x3.A 0.48789f
C9 bb[6] x1/x3.B 0.01836f
C10 SB[1] S[1] 0.05837f
C11 x2/x4.A VDD 0.31708f
C12 x4/x3.B S[4] 0.11239f
C13 x2/x4.B bb[8] 0.02487f
C14 x4/x3.A S[4] 0.17548f
C15 b[8] x3/x3.B 0.06214f
C16 bb[6] bb[8] 0.39479f
C17 b[9] VDD 0.67375f
C18 b[6] bb[7] 0.0823f
C19 VDD SB[4] 0.19141f
C20 x3/x3.A x3/x3.B 0.28615f
C21 x2/x5.Y bb[8] 0.02389f
C22 S[2] VDD 0.45155f
C23 x2/x4.C bb[9] 0.56698f
C24 bb[6] x2/x4.B 0.02952f
C25 VDD SB[2] 0.18329f
C26 VDD bb[7] 1.52111f
C27 x2/x4.B x2/x5.Y 0.04842f
C28 b[8] x4/x3.B 0.0151f
C29 b[8] x4/x3.A 0.15683f
C30 x2/x4.A x2/x4.C 0.01642f
C31 bb[6] x2/x5.Y 0.26143f
C32 bb[6] SB[1] 0.03872f
C33 b[7] b[8] 1.604f
C34 SB[4] S[4] 0.0648f
C35 bb[6] x3/x3.B 0.04268f
C36 b[7] x3/x3.A 0.01426f
C37 b[6] VDD 1.58049f
C38 S[2] x2/x4.C 0.05364f
C39 b[8] bb[9] 0.02535f
C40 bb[9] S[1] 0.0499f
C41 bb[7] S[3] 0.21691f
C42 x2/x4.C bb[7] 0.02737f
C43 x1/x3.A bb[9] 0.10418f
C44 bb[7] SB[3] 0.02755f
C45 b[8] x2/x4.A 0.01733f
C46 b[7] bb[8] 0.17431f
C47 x1/x3.B bb[9] 0.24146f
C48 b[8] b[9] 1.73039f
C49 bb[8] bb[9] 2.47438f
C50 x2/x4.B b[7] 0.05963f
C51 b[6] x2/x4.C 0.20013f
C52 x3/x3.A b[9] 0.18934f
C53 bb[6] b[7] 0.12948f
C54 b[6] S[4] 0.02557f
C55 S[2] S[1] 0.01308f
C56 x2/x4.B bb[9] 0.22399f
C57 b[8] bb[7] 0.11379f
C58 x2/x4.A bb[8] 0.18555f
C59 bb[7] S[1] 0.06935f
C60 VDD S[3] 0.30353f
C61 bb[6] bb[9] 0.28516f
C62 VDD x2/x4.C 0.25864f
C63 b[9] bb[8] 0.06634f
C64 VDD S[4] 0.4088f
C65 x2/x4.B x2/x4.A 0.77374f
C66 x1/x3.A bb[7] 0.14095f
C67 x2/x5.Y bb[9] 0.01838f
C68 VDD SB[3] 0.17952f
C69 x1/x3.B bb[7] 0.02024f
C70 S[2] bb[8] 0.03119f
C71 bb[6] x2/x4.A 0.04063f
C72 x2/x4.B b[9] 0.01203f
C73 bb[8] SB[2] 0.01815f
C74 bb[7] bb[8] 1.71241f
C75 b[6] b[8] 0.94458f
C76 x2/x4.A x2/x5.Y 0.0249f
C77 bb[6] b[9] 0.06734f
C78 S[2] x2/x4.B 0.14478f
C79 bb[6] SB[4] 0.01172f
C80 x4/x3.A x4/x3.B 0.18203f
C81 b[6] x3/x3.A 0.12678f
C82 x2/x4.B bb[7] 0.01119f
C83 S[2] bb[6] 0.11507f
C84 b[8] VDD 0.82193f
C85 bb[6] SB[2] 0.03033f
C86 VDD S[1] 0.26736f
C87 b[7] x4/x3.B 0.0979f
C88 b[7] x4/x3.A 0.05552f
C89 bb[6] bb[7] 1.98066f
C90 S[3] SB[3] 0.06166f
C91 S[2] x2/x5.Y 0.02252f
C92 x3/x3.A VDD 0.59342f
C93 b[6] bb[8] 0.06793f
C94 b[9] x3/x3.B 0.01904f
C95 x1/x3.A VDD 0.33716f
C96 x2/x5.Y bb[7] 0.22293f
C97 VDD x1/x3.B 0.25876f
C98 bb[7] SB[1] 0.02914f
C99 b[6] x2/x4.B 0.04129f
C100 b[7] bb[9] 0.07544f
C101 VDD bb[8] 0.7778f
C102 x3/x3.B bb[7] 0.3076f
C103 b[6] bb[6] 0.06741f
C104 S[3] S[1] 0.01483f
C105 b[8] x2/x4.C 0.0386f
C106 b[9] x4/x3.B 0.04039f
C107 x2/x4.B VDD 0.25711f
C108 b[9] x4/x3.A 0.06751f
C109 x3/x3.A S[3] 0.21439f
C110 b[7] x2/x4.A 0.03671f
C111 bb[6] VDD 2.03244f
C112 b[7] b[9] 0.21615f
C113 x2/x4.A bb[9] 0.09901f
C114 b[6] x3/x3.B 0.15193f
C115 x2/x5.Y VDD 0.49397f
C116 x2/x4.C bb[8] 0.01032f
C117 b[9] bb[9] 0.01319f
C118 VDD SB[1] 0.18056f
C119 VDD x3/x3.B 0.4727f
C120 S[2] bb[9] 0.05784f
C121 x2/x4.B x2/x4.C 0.60657f
C122 bb[9] SB[2] 0.02527f
C123 b[9] x2/x4.A 0.07319f
C124 bb[7] bb[9] 0.10932f
C125 bb[6] S[3] 0.04467f
C126 x3/x3.A b[8] 0.19756f
C127 bb[6] x2/x4.C 0.04624f
C128 b[6] x4/x3.B 0.29967f
C129 b[6] x4/x3.A 0.04884f
C130 bb[6] S[4] 0.02711f
C131 S[2] x2/x4.A 0.24608f
C132 x1/x3.A S[1] 0.09198f
C133 bb[6] SB[3] 0.02906f
C134 x2/x5.Y x2/x4.C 0.15447f
C135 x1/x3.B S[1] 0.14368f
C136 b[6] b[7] 2.22369f
C137 VDD x4/x3.B 0.29439f
C138 b[8] bb[8] 0.3493f
C139 VDD x4/x3.A 0.32055f
C140 bb[8] S[1] 0.03303f
C141 x1/x3.A x1/x3.B 0.13753f
C142 x3/x3.B S[3] 0.0651f
C143 b[6] bb[9] 0.1254f
C144 S[2] SB[2] 0.05715f
C145 b[7] VDD 0.64562f
C146 x2/x4.B b[8] 0.01469f
C147 x1/x3.A bb[8] 0.06718f
C148 S[2] bb[7] 0.04673f
C149 x1/x3.B bb[8] 0.09248f
C150 SB[2] GND 0.1621f
C151 S[2] GND 0.41125f
C152 SB[1] GND 0.15239f
C153 SB[3] GND 0.13905f
C154 S[3] GND 0.35805f
C155 S[1] GND 0.53545f
C156 SB[4] GND 0.1485f
C157 bb[9] GND 1.22111f
C158 bb[8] GND 0.7447f
C159 bb[7] GND 1.53581f
C160 bb[6] GND 1.06674f
C161 S[4] GND 0.36132f
C162 b[6] GND 2.12314f
C163 b[7] GND 0.94529f
C164 b[8] GND 1.54472f
C165 b[9] GND 1.27579f
C166 VDD GND 11.76536f
C167 x2/x4.A GND 0.89795f
C168 x2/x4.B GND 0.43129f
C169 x2/x4.C GND 0.41895f
C170 x2/x5.Y GND 0.45514f
C171 x3/x3.A GND 0.26387f
C172 x3/x3.B GND 0.32651f
C173 x1/x3.A GND 0.5014f
C174 x1/x3.B GND 0.44412f
C175 x4/x3.A GND 0.68096f
C176 x4/x3.B GND 0.40117f
C177 bb[9].t4 GND 0.04041f
C178 bb[9].t5 GND 0.02522f
C179 bb[9].n0 GND 0.08034f
C180 bb[9].t1 GND 0.04046f
C181 bb[9].t0 GND 0.02526f
C182 bb[9].n1 GND 0.07702f
C183 bb[9].n2 GND 0.1206f
C184 bb[9].n3 GND 1.43173f
C185 bb[9].n4 GND 0.33953f
C186 bb[9].t2 GND 0.04046f
C187 bb[9].t3 GND 0.02526f
C188 bb[9].n5 GND 0.07702f
C189 bb[9].n6 GND 0.01086f
C190 bb[6].t0 GND 0.0304f
C191 bb[6].t1 GND 0.019f
C192 bb[6].n0 GND 0.05344f
C193 bb[6].n1 GND 0.0951f
C194 bb[6].t2 GND 0.01937f
C195 bb[6].t3 GND 0.03084f
C196 bb[6].n2 GND 0.04176f
C197 bb[6].n3 GND 0.18254f
C198 bb[6].n4 GND 0.88317f
C199 bb[6].n5 GND 0.40624f
C200 bb[6].t4 GND 0.03026f
C201 bb[6].t5 GND 0.01888f
C202 bb[6].n6 GND 0.05953f
C203 bb[6].n7 GND 0.05649f
C204 b[6].t4 GND 0.03325f
C205 b[6].t5 GND 0.02076f
C206 b[6].n0 GND 0.06328f
C207 b[6].n1 GND 0.11027f
C208 b[6].n2 GND 0.36709f
C209 b[6].t0 GND 0.02125f
C210 b[6].t1 GND 0.03384f
C211 b[6].n3 GND 0.05099f
C212 b[6].n4 GND 1.00668f
C213 b[6].t2 GND 0.03325f
C214 b[6].t3 GND 0.02076f
C215 b[6].n5 GND 0.06328f
C216 b[6].n6 GND 0.14263f
C217 bb[8].t2 GND 0.04117f
C218 bb[8].t3 GND 0.02569f
C219 bb[8].n0 GND 0.081f
C220 bb[8].n1 GND 0.13128f
C221 bb[8].n2 GND 1.58778f
C222 bb[8].t0 GND 0.04122f
C223 bb[8].t1 GND 0.02574f
C224 bb[8].n3 GND 0.07846f
C225 bb[8].n4 GND 0.37631f
C226 VDD.t14 GND 0.01149f
C227 VDD.t10 GND 0.01536f
C228 VDD.t4 GND 0.01149f
C229 VDD.t2 GND 0.01551f
C230 VDD.t31 GND 0.01014f
C231 VDD.t34 GND 0.02535f
C232 VDD.n13 GND 0.01361f
C233 VDD.n14 GND 0.01277f
C234 VDD.n46 GND 0.01096f
C235 VDD.n53 GND 0.01277f
C236 VDD.n66 GND 0.03404f
C237 VDD.t63 GND 0.01105f
C238 VDD.t42 GND 0.01105f
C239 VDD.t72 GND 0.01105f
C240 VDD.t36 GND 0.01604f
C241 VDD.t57 GND 0.01315f
C242 VDD.t49 GND 0.01736f
C243 VDD.n67 GND 0.01831f
C244 VDD.t47 GND 0.01105f
C245 VDD.t53 GND 0.01105f
C246 VDD.t20 GND 0.01105f
C247 VDD.t22 GND 0.01841f
C248 VDD.n68 GND 0.01489f
C249 VDD.t51 GND 0.01184f
C250 VDD.t16 GND 0.01263f
C251 VDD.t40 GND 0.02722f
C252 VDD.t27 GND 0.01381f
C253 VDD.t29 GND 0.01105f
C254 VDD.t45 GND 0.0167f
C255 VDD.t32 GND 0.01894f
C256 VDD.n69 GND 0.01489f
C257 VDD.t6 GND 0.0121f
C258 VDD.n70 GND 0.01937f
C259 VDD.t25 GND 0.05152f
C260 VDD.n71 GND 0.05294f
C261 VDD.n72 GND 0.09131f
C262 VDD.n73 GND 0.08615f
C263 VDD.n74 GND 0.0258f
C264 VDD.n112 GND 0.02173f
C265 VDD.t38 GND 0.02185f
C266 VDD.t18 GND 0.01574f
C267 VDD.t24 GND 0.01014f
C268 VDD.t61 GND 0.01551f
C269 VDD.t59 GND 0.01149f
C270 VDD.t8 GND 0.01536f
C271 VDD.t67 GND 0.01149f
C272 VDD.n113 GND 0.01799f
C273 VDD.n115 GND 0.11394f
C274 b[7].t0 GND 0.04098f
C275 b[7].t5 GND 0.02558f
C276 b[7].n0 GND 0.08068f
C277 b[7].n1 GND 0.1138f
C278 b[7].n2 GND 0.42412f
C279 b[7].t3 GND 0.02567f
C280 b[7].t4 GND 0.04109f
C281 b[7].n3 GND 0.07558f
C282 b[7].n4 GND 0.07213f
C283 b[7].n5 GND 0.94143f
C284 b[7].t2 GND 0.04098f
C285 b[7].t1 GND 0.02558f
C286 b[7].n6 GND 0.08063f
C287 b[7].n7 GND 0.11679f
.ends

