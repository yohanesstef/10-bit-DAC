magic
tech sky130A
magscale 1 2
timestamp 1749908815
<< error_p >>
rect -224 -398 -194 330
rect -158 -332 -128 264
rect 128 -332 158 264
rect -158 -336 158 -332
rect 194 -398 224 330
rect -224 -402 224 -398
<< nwell >>
rect -194 -398 194 364
<< mvpmos >>
rect -100 -336 100 264
<< mvpdiff >>
rect -158 252 -100 264
rect -158 -324 -146 252
rect -112 -324 -100 252
rect -158 -336 -100 -324
rect 100 252 158 264
rect 100 -324 112 252
rect 146 -324 158 252
rect 100 -336 158 -324
<< mvpdiffc >>
rect -146 -324 -112 252
rect 112 -324 146 252
<< poly >>
rect -100 345 100 361
rect -100 311 -84 345
rect 84 311 100 345
rect -100 264 100 311
rect -100 -362 100 -336
<< polycont >>
rect -84 311 84 345
<< locali >>
rect -100 311 -84 345
rect 84 311 100 345
rect -146 252 -112 268
rect -146 -340 -112 -324
rect 112 252 146 268
rect 112 -340 146 -324
<< viali >>
rect -63 311 63 345
rect -146 -252 -112 180
rect 112 -252 146 180
<< metal1 >>
rect -75 345 75 351
rect -75 311 -63 345
rect 63 311 75 345
rect -75 305 75 311
rect -152 180 -106 192
rect -152 -252 -146 180
rect -112 -252 -106 180
rect -152 -264 -106 -252
rect 106 180 152 192
rect 106 -252 112 180
rect 146 -252 152 180
rect 106 -264 152 -252
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 75 viadrn 75 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
