magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1114 307 1114
<< psubdiff >>
rect -271 1044 -175 1078
rect 175 1044 271 1078
rect -271 982 -237 1044
rect 237 982 271 1044
rect -271 -1044 -237 -982
rect 237 -1044 271 -982
rect -271 -1078 -175 -1044
rect 175 -1078 271 -1044
<< psubdiffcont >>
rect -175 1044 175 1078
rect -271 -982 -237 982
rect 237 -982 271 982
rect -175 -1078 175 -1044
<< xpolycontact >>
rect -141 516 141 948
rect -141 -948 141 -516
<< xpolyres >>
rect -141 -516 141 516
<< locali >>
rect -271 1044 -175 1078
rect 175 1044 271 1078
rect -271 982 -237 1044
rect 237 982 271 1044
rect -271 -1044 -237 -982
rect 237 -1044 271 -982
rect -271 -1078 -175 -1044
rect 175 -1078 271 -1044
<< viali >>
rect -125 533 125 930
rect -125 -930 125 -533
<< metal1 >>
rect -131 930 131 942
rect -131 533 -125 930
rect 125 533 131 930
rect -131 521 131 533
rect -131 -533 131 -521
rect -131 -930 -125 -533
rect 125 -930 131 -533
rect -131 -942 131 -930
<< properties >>
string FIXED_BBOX -254 -1061 254 1061
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 5.32 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 7.813k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
