magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -791 307 791
<< psubdiff >>
rect -271 721 -175 755
rect 175 721 271 755
rect -271 659 -237 721
rect 237 659 271 721
rect -271 -721 -237 -659
rect 237 -721 271 -659
rect -271 -755 -175 -721
rect 175 -755 271 -721
<< psubdiffcont >>
rect -175 721 175 755
rect -271 -659 -237 659
rect 237 -659 271 659
rect -175 -755 175 -721
<< xpolycontact >>
rect -141 193 141 625
rect -141 -625 141 -193
<< xpolyres >>
rect -141 -193 141 193
<< locali >>
rect -271 721 -175 755
rect 175 721 271 755
rect -271 659 -237 721
rect 237 659 271 721
rect -271 -721 -237 -659
rect 237 -721 271 -659
rect -271 -755 -175 -721
rect 175 -755 271 -721
<< viali >>
rect -125 210 125 607
rect -125 -607 125 -210
<< metal1 >>
rect -131 607 131 619
rect -131 210 -125 607
rect 125 210 131 607
rect -131 198 131 210
rect -131 -210 131 -198
rect -131 -607 -125 -210
rect 125 -607 131 -210
rect -131 -619 131 -607
<< properties >>
string FIXED_BBOX -254 -738 254 738
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 2.091 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 3.232k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
