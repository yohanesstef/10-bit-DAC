magic
tech sky130A
magscale 1 2
timestamp 1749552768
<< locali >>
rect 5445 5062 5479 5814
rect 8079 5051 8113 5780
rect 10713 5028 10747 5814
<< metal1 >>
rect 6549 6630 6609 6636
rect 5389 6454 5449 6460
rect 5200 6278 5260 6284
rect 5200 6130 5260 6218
rect 5201 6022 5241 6130
rect 5201 5928 5261 6022
rect 5389 5928 5449 6394
rect 6361 6454 6421 6460
rect 5665 6366 5725 6372
rect 5477 6190 5537 6196
rect 5537 6130 5543 6190
rect 5477 6022 5517 6130
rect 5477 5928 5537 6022
rect 5665 5928 5725 6306
rect 5969 6366 6029 6372
rect 5781 6278 5841 6284
rect 5781 6130 5841 6218
rect 5781 6022 5821 6130
rect 5781 5928 5841 6022
rect 5969 5928 6029 6306
rect 6245 6278 6305 6284
rect 6057 6190 6117 6196
rect 6117 6130 6123 6190
rect 6057 6022 6097 6130
rect 6057 5928 6117 6022
rect 6245 5928 6305 6218
rect 6361 6190 6421 6394
rect 6355 6130 6361 6190
rect 6421 6130 6427 6190
rect 6361 6022 6401 6130
rect 6361 5928 6421 6022
rect 6549 5928 6609 6570
rect 6825 6542 6885 6548
rect 6637 6366 6697 6373
rect 6637 6130 6697 6306
rect 6637 6022 6677 6130
rect 6637 5928 6697 6022
rect 6825 5928 6885 6482
rect 7101 6454 7161 6460
rect 6913 6278 6973 6284
rect 6913 6130 6973 6218
rect 6913 6022 6953 6130
rect 6913 5928 6973 6022
rect 7101 5928 7161 6394
rect 7405 6454 7465 6460
rect 7189 6190 7249 6196
rect 7189 5928 7249 6130
rect 7405 5928 7465 6394
rect 7493 6366 7553 6372
rect 7493 6130 7553 6306
rect 7681 6366 7741 6372
rect 7493 6022 7533 6130
rect 7493 5928 7553 6022
rect 7681 5928 7741 6306
rect 7769 6278 7829 6284
rect 7769 6130 7829 6218
rect 7957 6278 8017 6284
rect 7769 6022 7809 6130
rect 7769 5928 7829 6022
rect 7957 5928 8017 6218
rect 8351 5108 8411 6012
rect 8627 5196 8687 6012
rect 8903 5284 8963 6012
rect 9179 5372 9239 6012
rect 9455 5460 9515 6012
rect 9723 5812 9783 6012
rect 10003 5900 10059 6012
rect 10279 5900 10335 6012
rect 10555 5900 10611 6012
rect 10831 5900 10887 6012
rect 9723 5746 9783 5752
rect 9999 5724 10059 5900
rect 9999 5658 10059 5664
rect 10275 5636 10335 5900
rect 10275 5570 10335 5576
rect 10551 5548 10611 5900
rect 10551 5482 10611 5488
rect 9455 5394 9515 5400
rect 10827 5460 10887 5900
rect 10827 5394 10887 5400
rect 9179 5306 9239 5312
rect 8903 5218 8963 5224
rect 8627 5130 8687 5136
rect 8351 5042 8411 5048
rect 5730 4554 5790 4842
rect 6006 4642 6066 4842
rect 6282 4730 6342 4842
rect 6558 4730 6618 4842
rect 6282 4670 6414 4730
rect 6006 4582 6326 4642
rect 5730 4494 6238 4554
rect 6178 4026 6238 4494
rect 6266 4026 6326 4582
rect 6354 4026 6414 4670
rect 6442 4670 6618 4730
rect 6442 4026 6502 4670
rect 6821 4642 6881 4842
rect 6530 4582 6881 4642
rect 6530 4026 6590 4582
rect 7097 4554 7157 4842
rect 6618 4494 7157 4554
rect 6618 4026 6678 4494
rect 7373 4466 7433 4842
rect 6706 4406 7433 4466
rect 6706 4026 6766 4406
rect 7649 4378 7709 4842
rect 6794 4318 7709 4378
rect 6794 4026 6854 4318
rect 7925 4290 7985 4842
rect 8346 4730 8406 4842
rect 6882 4230 7985 4290
rect 8286 4670 8406 4730
rect 6882 4026 6942 4230
rect 8286 4010 8346 4670
rect 8627 4642 8687 4841
rect 8374 4582 8687 4642
rect 8374 4026 8434 4582
rect 8903 4554 8963 4842
rect 8568 4553 8963 4554
rect 8462 4494 8963 4553
rect 8462 4026 8522 4494
rect 9179 4466 9239 4842
rect 8550 4406 9239 4466
rect 8550 4026 8610 4406
rect 9455 4378 9515 4842
rect 8638 4318 9515 4378
rect 8638 4026 8698 4318
rect 9731 4290 9791 4842
rect 8726 4230 9791 4290
rect 8726 4026 8786 4230
rect 10007 4202 10067 4842
rect 8814 4142 10067 4202
rect 8814 4026 8874 4142
rect 10283 4114 10343 4842
rect 8902 4054 10343 4114
rect 8902 4026 8962 4054
rect 10559 4026 10619 4842
rect 8990 3966 10619 4026
<< via1 >>
rect 6549 6570 6609 6630
rect 5389 6394 5449 6454
rect 5200 6218 5260 6278
rect 6361 6394 6421 6454
rect 5665 6306 5725 6366
rect 5477 6130 5537 6190
rect 5969 6306 6029 6366
rect 5781 6218 5841 6278
rect 6245 6218 6305 6278
rect 6057 6130 6117 6190
rect 6361 6130 6421 6190
rect 6825 6482 6885 6542
rect 6637 6306 6697 6366
rect 7101 6394 7161 6454
rect 6913 6218 6973 6278
rect 7405 6394 7465 6454
rect 7189 6130 7249 6190
rect 7493 6306 7553 6366
rect 7681 6306 7741 6366
rect 7769 6218 7829 6278
rect 7957 6218 8017 6278
rect 9723 5752 9783 5812
rect 9999 5664 10059 5724
rect 10275 5576 10335 5636
rect 10551 5488 10611 5548
rect 9455 5400 9515 5460
rect 10827 5400 10887 5460
rect 9179 5312 9239 5372
rect 8903 5224 8963 5284
rect 8627 5136 8687 5196
rect 8351 5048 8411 5108
<< metal2 >>
rect 6543 6570 6549 6630
rect 6609 6570 9981 6630
rect 6819 6482 6825 6542
rect 6885 6482 10257 6542
rect 5383 6394 5389 6454
rect 5449 6394 6361 6454
rect 6421 6394 6427 6454
rect 7095 6394 7101 6454
rect 7161 6394 7405 6454
rect 7465 6394 10533 6454
rect 5659 6306 5665 6366
rect 5725 6306 5969 6366
rect 6029 6306 6637 6366
rect 6697 6306 7493 6366
rect 7553 6306 7559 6366
rect 7675 6306 7681 6366
rect 7741 6306 10809 6366
rect 5194 6218 5200 6278
rect 5260 6218 5781 6278
rect 5841 6218 5847 6278
rect 6219 6218 6245 6278
rect 6305 6218 6913 6278
rect 6973 6218 7769 6278
rect 7829 6218 7835 6278
rect 7951 6218 7957 6278
rect 8017 6218 11085 6278
rect 5471 6130 5477 6190
rect 5537 6130 6057 6190
rect 6117 6130 6123 6190
rect 6355 6130 6361 6190
rect 6421 6130 7189 6190
rect 7249 6130 7255 6190
rect 7744 5752 9723 5812
rect 9783 5752 10450 5812
rect 7468 5664 9999 5724
rect 10059 5664 10174 5724
rect 7192 5576 10275 5636
rect 10335 5576 10341 5636
rect 6916 5488 10551 5548
rect 10611 5488 10617 5548
rect 6640 5400 9455 5460
rect 9515 5400 10827 5460
rect 10887 5400 10893 5460
rect 6364 5312 9179 5372
rect 9239 5312 9245 5372
rect 6088 5224 8903 5284
rect 8963 5224 8969 5284
rect 5812 5136 8627 5196
rect 8687 5136 8693 5196
rect 5602 5048 8351 5108
rect 8411 5048 8417 5108
use hpmos_9  hpmos_9_0 ~/10-bit-DAC/mag
timestamp 1749528210
transform 1 0 3159 0 1 3796
box 2208 736 5032 2022
use hpmos_9  hpmos_9_1
timestamp 1749528210
transform 1 0 5793 0 1 3796
box 2208 736 5032 2022
use rseg_3_v3  rseg_3_v3_0 ~/10-bit-DAC/mag
timestamp 1749552768
transform 1 0 -6844 0 1 5644
box 12478 -5378 17402 -1618
use tps3_switch_10  tps3_switch_10_0 ~/10-bit-DAC/mag
timestamp 1749525104
transform 1 0 8035 0 1 5711
box -34 -9 3216 925
use tps3_switch_final_stage  tps3_switch_final_stage_0 ~/10-bit-DAC/mag
timestamp 1749520983
transform 1 0 6315 0 1 5868
box -1308 -166 1876 442
<< labels >>
flabel metal2 s 5634 3322 5634 3322 4 FreeSans 800 0 0 0 V0
port 0 se
flabel metal2 s 10558 3322 10558 3322 6 FreeSans 800 0 0 0 V16
port 1 sw
flabel metal2 s 5761 6098 5761 6098 4 FreeSans 320 0 0 0 b[3]
port 2 se
flabel metal2 s 7199 6100 7199 6100 4 FreeSans 320 0 0 0 b[4]
port 3 se
flabel metal2 s 8174 6097 8174 6097 4 FreeSans 320 0 0 0 b[5]
port 4 se
flabel metal2 s 8177 4929 8177 4929 4 FreeSans 320 0 0 0 b[6]
port 5 se
flabel metal2 s 5186 6099 5186 6099 4 FreeSans 320 0 0 0 bb[3]
port 6 se
flabel metal2 s 6362 6090 6362 6090 4 FreeSans 320 0 0 0 bb[4]
port 7 se
flabel metal2 s 9755 6084 9755 6084 4 FreeSans 320 0 0 0 bb[5]
port 8 se
flabel metal2 s 5602 4912 5602 4912 4 FreeSans 320 0 0 0 bb[6]
port 9 se
flabel metal2 s 5202 6266 5202 6266 4 FreeSans 320 0 0 0 VH
port 10 se
flabel metal2 s 5501 6178 5501 6178 4 FreeSans 320 0 0 0 VL
port 11 se
flabel locali s 5706 3778 5706 3778 4 FreeSans 320 0 0 0 GND
port 12 se
flabel locali s 5477 4636 5477 4636 4 FreeSans 320 0 0 0 VPB
port 13 se
<< end >>
