magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -894 307 894
<< psubdiff >>
rect -271 824 -175 858
rect 175 824 271 858
rect -271 762 -237 824
rect 237 762 271 824
rect -271 -824 -237 -762
rect 237 -824 271 -762
rect -271 -858 -175 -824
rect 175 -858 271 -824
<< psubdiffcont >>
rect -175 824 175 858
rect -271 -762 -237 762
rect 237 -762 271 762
rect -175 -858 175 -824
<< xpolycontact >>
rect -141 296 141 728
rect -141 -728 141 -296
<< xpolyres >>
rect -141 -296 141 296
<< locali >>
rect -271 824 -175 858
rect 175 824 271 858
rect -271 762 -237 824
rect 237 762 271 824
rect -271 -824 -237 -762
rect 237 -824 271 -762
rect -271 -858 -175 -824
rect 175 -858 271 -824
<< viali >>
rect -125 313 125 710
rect -125 -710 125 -313
<< metal1 >>
rect -131 710 131 722
rect -131 313 -125 710
rect 125 313 131 710
rect -131 301 131 313
rect -131 -313 131 -301
rect -131 -710 -125 -313
rect 125 -710 131 -313
rect -131 -722 131 -710
<< properties >>
string FIXED_BBOX -254 -841 254 841
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 3.116 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 4.686k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
