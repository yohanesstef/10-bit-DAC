.subckt rseg_4_v3 v0 v1 v2 v3 v4 v5 v6 v7 v8 v9 v10 v11 v12 v13 v14 v15 v16 v17 v18 v19 v20 v21 v22 v23 v24 v25 v26 v27 v28 v29 v30 v31 v32 v33 v34 v35 v36 v37 v38 v39 v40 v41 v42 v43 v44 v45 v46 v47 v48 v49 v50 v51 v52 v53 v54 v55 v56 v57 v58 v59 v60 v61 v62 v63 gnd
XRD1 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.5538 mult=1 m=1
XRD8 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6050 mult=1 m=1
XRD9 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6050 mult=1 m=1
XRD16 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6563 mult=1 m=1
XRD17 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7074 mult=1 m=1
XRD24 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7587 mult=1 m=1
XRD25 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7587 mult=1 m=1
XRD32 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.8100 mult=1 m=1
XRD33 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.8612 mult=1 m=1
XRD40 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.0150 mult=1 m=1
XRD41 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.0150 mult=1 m=1
XRD48 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.2200 mult=1 m=1
XRD49 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.2713 mult=1 m=1
XRD56 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.6300 mult=1 m=1
XRD57 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.7326 mult=1 m=1
XRD63 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=2.5526 mult=1 m=1
XRD64 gnd gnd gnd sky130_fd_pr__res_xhigh_po_1p41 L=2.5526 mult=1 m=1

XR1 v0 v1 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.5538 mult=1 m=1
XR2 v1 v2 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.5537 mult=1 m=1
XR3 v2 v3 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6050 mult=1 m=1
XR4 v3 v4 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.5537 mult=1 m=1
XR5 v4 v5 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6050 mult=1 m=1
XR6 v5 v6 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.5537 mult=1 m=1
XR7 v6 v7 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6050 mult=1 m=1
XR8 v7 v8 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6050 mult=1 m=1
XR9 v8 v9 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6050 mult=1 m=1
XR10 v9 v10 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6563 mult=1 m=1
XR11 v10 v11 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6050 mult=1 m=1
XR12 v11 v12 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6563 mult=1 m=1
XR13 v12 v13 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6050 mult=1 m=1
XR14 v13 v14 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6563 mult=1 m=1
XR15 v14 v15 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6563 mult=1 m=1
XR16 v15 v16 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6563 mult=1 m=1
XR17 v16 v17 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7074 mult=1 m=1
XR18 v17 v18 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.6563 mult=1 m=1
XR19 v18 v19 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7074 mult=1 m=1
XR20 v19 v20 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7074 mult=1 m=1
XR21 v20 v21 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7074 mult=1 m=1
XR22 v21 v22 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7074 mult=1 m=1
XR23 v22 v23 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7587 mult=1 m=1
XR24 v23 v24 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7587 mult=1 m=1
XR25 v24 v25 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7587 mult=1 m=1
XR26 v25 v26 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7587 mult=1 m=1
XR27 v26 v27 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.7587 mult=1 m=1
XR28 v27 v28 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.8100 mult=1 m=1
XR29 v28 v29 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.8100 mult=1 m=1
XR30 v29 v30 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.8100 mult=1 m=1
XR31 v30 v31 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.8612 mult=1 m=1
XR32 v31 v32 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.8100 mult=1 m=1
XR33 v32 v33 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.8612 mult=1 m=1
XR34 v33 v34 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.9125 mult=1 m=1
XR35 v34 v35 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.8612 mult=1 m=1
XR36 v35 v36 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.9638 mult=1 m=1
XR37 v36 v37 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.9125 mult=1 m=1
XR38 v37 v38 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.9638 mult=1 m=1
XR39 v38 v39 gnd sky130_fd_pr__res_xhigh_po_1p41 L=0.9638 mult=1 m=1
XR40 v39 v40 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.0150 mult=1 m=1
XR41 v40 v41 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.0150 mult=1 m=1
XR42 v41 v42 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.0150 mult=1 m=1
XR43 v42 v43 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.0663 mult=1 m=1
XR44 v43 v44 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.1175 mult=1 m=1
XR45 v44 v45 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.1175 mult=1 m=1
XR46 v45 v46 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.1687 mult=1 m=1
XR47 v46 v47 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.1687 mult=1 m=1
XR48 v47 v48 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.2200 mult=1 m=1
XR49 v48 v49 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.2713 mult=1 m=1
XR50 v49 v50 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.2713 mult=1 m=1
XR51 v50 v51 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.3738 mult=1 m=1
XR52 v51 v52 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.3738 mult=1 m=1
XR53 v52 v53 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.4763 mult=1 m=1
XR54 v53 v54 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.4763 mult=1 m=1
XR55 v54 v55 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.5788 mult=1 m=1
XR56 v55 v56 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.6300 mult=1 m=1
XR57 v56 v57 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.7326 mult=1 m=1
XR58 v57 v58 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.7838 mult=1 m=1
XR59 v58 v59 gnd sky130_fd_pr__res_xhigh_po_1p41 L=1.9375 mult=1 m=1
XR60 v59 v60 gnd sky130_fd_pr__res_xhigh_po_1p41 L=2.0401 mult=1 m=1
XR61 v60 v61 gnd sky130_fd_pr__res_xhigh_po_1p41 L=2.1426 mult=1 m=1
XR62 v61 v62 gnd sky130_fd_pr__res_xhigh_po_1p41 L=2.3988 mult=1 m=1
XR63 v62 v63 gnd sky130_fd_pr__res_xhigh_po_1p41 L=2.5526 mult=1 m=1
.ends