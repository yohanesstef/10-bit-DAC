magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1170 307 1170
<< psubdiff >>
rect -271 1100 -175 1134
rect 175 1100 271 1134
rect -271 1038 -237 1100
rect 237 1038 271 1100
rect -271 -1100 -237 -1038
rect 237 -1100 271 -1038
rect -271 -1134 -175 -1100
rect 175 -1134 271 -1100
<< psubdiffcont >>
rect -175 1100 175 1134
rect -271 -1038 -237 1038
rect 237 -1038 271 1038
rect -175 -1134 175 -1100
<< xpolycontact >>
rect -141 572 141 1004
rect -141 -1004 141 -572
<< xpolyres >>
rect -141 -572 141 572
<< locali >>
rect -271 1100 -175 1134
rect 175 1100 271 1134
rect -271 1038 -237 1100
rect 237 1038 271 1100
rect -271 -1100 -237 -1038
rect 237 -1100 271 -1038
rect -271 -1134 -175 -1100
rect 175 -1134 271 -1100
<< viali >>
rect -125 589 125 986
rect -125 -986 125 -589
<< metal1 >>
rect -131 986 131 998
rect -131 589 -125 986
rect 125 589 131 986
rect -131 577 131 589
rect -131 -589 131 -577
rect -131 -986 -125 -589
rect 125 -986 131 -589
rect -131 -998 131 -986
<< properties >>
string FIXED_BBOX -254 -1117 254 1117
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 5.884 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 8.613k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
