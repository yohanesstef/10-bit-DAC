magic
tech sky130A
timestamp 1749229935
<< error_p >>
rect -87 52 87 54
rect -87 -52 -72 52
rect -54 19 54 21
rect -54 -19 -39 19
rect 39 -19 54 19
rect -54 -21 54 -19
rect 72 -52 87 52
rect -87 -54 87 -52
<< nwell >>
rect -72 -52 72 52
<< mvpmos >>
rect -25 -21 25 21
<< mvpdiff >>
rect -54 15 -25 21
rect -54 -15 -48 15
rect -31 -15 -25 15
rect -54 -21 -25 -15
rect 25 15 54 21
rect 25 -15 31 15
rect 48 -15 54 15
rect 25 -21 54 -15
<< mvpdiffc >>
rect -48 -15 -31 15
rect 31 -15 48 15
<< poly >>
rect -25 21 25 34
rect -25 -34 25 -21
<< locali >>
rect -48 15 -31 23
rect -48 -23 -31 -15
rect 31 15 48 23
rect 31 -23 48 -15
<< viali >>
rect -48 -15 -31 15
rect 31 -15 48 15
<< metal1 >>
rect -51 15 -28 21
rect -51 -15 -48 15
rect -31 -15 -28 15
rect -51 -21 -28 -15
rect 28 15 51 21
rect 28 -15 31 15
rect 48 -15 51 15
rect 28 -21 51 -15
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 0.50 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
