magic
tech sky130A
magscale 1 2
timestamp 1743275510
<< pwell >>
rect -201 -667 201 667
<< psubdiff >>
rect -165 597 -69 631
rect 69 597 165 631
rect -165 535 -131 597
rect 131 535 165 597
rect -165 -597 -131 -535
rect 131 -597 165 -535
rect -165 -631 -69 -597
rect 69 -631 165 -597
<< psubdiffcont >>
rect -69 597 69 631
rect -165 -535 -131 535
rect 131 -535 165 535
rect -69 -631 69 -597
<< xpolycontact >>
rect -35 69 35 501
rect -35 -501 35 -69
<< xpolyres >>
rect -35 -69 35 69
<< locali >>
rect -165 597 -69 631
rect 69 597 165 631
rect -165 535 -131 597
rect 131 535 165 597
rect -165 -597 -131 -535
rect 131 -597 165 -535
rect -165 -631 -69 -597
rect 69 -631 165 -597
<< viali >>
rect -19 86 19 483
rect -19 -483 19 -86
<< metal1 >>
rect -25 483 25 495
rect -25 86 -19 483
rect 19 86 25 483
rect -25 74 25 86
rect -25 -86 25 -74
rect -25 -483 -19 -86
rect 19 -483 25 -86
rect -25 -495 25 -483
<< properties >>
string FIXED_BBOX -148 -614 148 614
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.846 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 5.909k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
