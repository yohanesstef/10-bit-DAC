magic
tech sky130A
magscale 1 2
timestamp 1749738669
<< nwell >>
rect 602 -1802 729 -1481
rect 2093 -1802 2158 -1481
<< pwell >>
rect 602 -1423 2158 -37
<< locali >>
rect 784 -1273 842 -1237
rect 1980 -1273 2038 -1237
rect 1047 -1485 1156 -1431
rect 1599 -1485 1773 -1431
rect 784 -1747 842 -1711
rect 1980 -1747 2038 -1711
<< viali >>
rect 893 -1478 927 -1444
rect 979 -1487 1013 -1427
rect 1255 -1487 1289 -1427
rect 1346 -1478 1380 -1444
rect 1444 -1480 1478 -1446
rect 1531 -1487 1565 -1427
rect 1807 -1487 1841 -1427
rect 1895 -1477 1929 -1443
<< metal1 >>
rect 668 1344 2092 1440
rect 914 1036 1034 1042
rect 914 976 920 1036
rect 1028 976 1034 1036
rect 914 973 1034 976
rect 1256 1036 1376 1042
rect 1256 976 1262 1036
rect 1370 976 1376 1036
rect 914 252 974 973
rect 1256 959 1376 976
rect 1598 1036 1718 1042
rect 1598 976 1604 1036
rect 1712 976 1718 1036
rect 1598 959 1718 976
rect 1940 1036 2060 1042
rect 1940 976 1946 1036
rect 2054 976 2060 1036
rect 1940 959 2060 976
rect 1256 252 1316 959
rect 1598 252 1658 959
rect 1940 252 2000 959
rect 821 200 1034 252
rect 1177 200 1376 252
rect 1533 200 1718 252
rect 1876 200 2060 252
rect 821 -68 933 200
rect 1177 -68 1289 200
rect 1533 -78 1645 200
rect 1889 -79 2001 200
rect 821 -552 933 -312
rect 1177 -552 1289 -312
rect 821 -952 950 -552
rect 930 -990 990 -984
rect 930 -1056 990 -1050
rect 668 -1268 767 -1172
rect 1025 -1199 1085 -755
rect 1166 -952 1289 -552
rect 1533 -552 1645 -312
rect 1889 -552 2001 -312
rect 1533 -952 1662 -552
rect 1120 -990 1180 -984
rect 1120 -1056 1180 -1050
rect 1642 -990 1702 -984
rect 1642 -1056 1702 -1050
rect 1737 -1180 1797 -736
rect 1872 -952 2001 -552
rect 1832 -990 1892 -984
rect 1832 -1056 1892 -1050
rect 2055 -1268 2092 -1172
rect 1332 -1393 1942 -1333
rect 968 -1427 1028 -1421
rect 1244 -1427 1304 -1421
rect 879 -1444 939 -1433
rect 879 -1478 893 -1444
rect 927 -1478 939 -1444
rect 879 -1521 939 -1478
rect 967 -1487 968 -1427
rect 1243 -1487 1244 -1427
rect 968 -1493 1028 -1487
rect 1244 -1493 1304 -1487
rect 1332 -1444 1392 -1393
rect 1520 -1427 1580 -1421
rect 1332 -1478 1346 -1444
rect 1380 -1478 1392 -1444
rect 1332 -1493 1392 -1478
rect 1431 -1446 1491 -1433
rect 1431 -1480 1444 -1446
rect 1478 -1480 1491 -1446
rect 1431 -1521 1491 -1480
rect 1519 -1487 1520 -1427
rect 1520 -1493 1580 -1487
rect 1794 -1427 1854 -1421
rect 1794 -1493 1854 -1487
rect 1882 -1443 1942 -1393
rect 1882 -1477 1895 -1443
rect 1929 -1477 1942 -1443
rect 1882 -1493 1942 -1477
rect 879 -1581 1491 -1521
rect 668 -1812 767 -1716
rect 2055 -1812 2092 -1716
<< via1 >>
rect 920 976 1028 1036
rect 1262 976 1370 1036
rect 1604 976 1712 1036
rect 1946 976 2054 1036
rect 930 -1050 990 -990
rect 1120 -1050 1180 -990
rect 1642 -1050 1702 -990
rect 1832 -1050 1892 -990
rect 968 -1487 979 -1427
rect 979 -1487 1013 -1427
rect 1013 -1487 1028 -1427
rect 1244 -1487 1255 -1427
rect 1255 -1487 1289 -1427
rect 1289 -1487 1304 -1427
rect 1520 -1487 1531 -1427
rect 1531 -1487 1565 -1427
rect 1565 -1487 1580 -1427
rect 1794 -1487 1807 -1427
rect 1807 -1487 1841 -1427
rect 1841 -1487 1854 -1427
<< metal2 >>
rect 914 1036 1034 1470
rect 914 976 920 1036
rect 1028 976 1034 1036
rect 1256 1036 1376 1470
rect 1256 976 1262 1036
rect 1370 976 1376 1036
rect 1598 1036 1718 1470
rect 1598 976 1604 1036
rect 1712 976 1718 1036
rect 1940 1036 2060 1470
rect 1940 976 1946 1036
rect 2054 976 2060 1036
rect 930 -990 990 -984
rect 930 -1427 990 -1050
rect 1120 -990 1180 -984
rect 1120 -1427 1180 -1050
rect 1642 -990 1702 -984
rect 1642 -1427 1702 -1050
rect 1832 -990 1892 -984
rect 1832 -1427 1892 -1050
rect 930 -1487 968 -1427
rect 1028 -1487 1034 -1427
rect 1120 -1487 1244 -1427
rect 1304 -1487 1310 -1427
rect 1514 -1487 1520 -1427
rect 1580 -1487 1702 -1427
rect 1788 -1487 1794 -1427
rect 1854 -1487 1892 -1427
use dec_logic  dec_logic_0
timestamp 1749645942
transform 1 0 341 0 -1 -1218
box 480 -46 1660 594
use dec_ncell_h  dec_ncell_h_0
timestamp 1749656061
transform 1 0 -21 0 1 -207
box 689 -291 2113 159
use dec_ncell_l_1  dec_ncell_l_0
timestamp 1749652636
transform 1 0 -504 0 1 851
box 1434 -1904 1684 -1377
use dec_ncell_l_1  dec_ncell_l_1_0
timestamp 1749652636
transform 1 0 208 0 1 851
box 1434 -1904 1684 -1377
use dec_pcell  dec_pcell_0
timestamp 1749654170
transform 1 0 1203 0 1 -479
box -601 499 955 1949
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 767 0 -1 -1220
box -38 -48 130 592
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_1
timestamp 1704896540
transform 1 0 1963 0 -1 -1220
box -38 -48 130 592
<< labels >>
flabel metal1 s 683 1133 683 1133 3 FreeSans 480 0 0 0 VPBIAS
port 0 e
flabel metal1 s 679 -208 679 -208 3 FreeSans 480 0 0 0 VNBIAS
port 1 e
flabel locali s 1343 -1456 1343 -1456 3 FreeSans 240 0 0 0 b[0]
port 2 e
flabel locali s 1623 -1460 1623 -1460 3 FreeSans 240 0 0 0 b[1]
port 3 e
flabel locali s 918 -1460 918 -1460 3 FreeSans 240 0 0 0 bb[0]
port 4 e
flabel locali s 1062 -1465 1062 -1465 3 FreeSans 240 0 0 0 bb[1]
port 5 e
flabel metal2 s 921 1436 921 1436 3 FreeSans 320 0 0 0 VOUT[0]
port 6 e
flabel metal2 s 1268 1433 1268 1433 3 FreeSans 320 0 0 0 VOUT[1]
port 7 e
flabel metal2 s 1607 1424 1607 1424 3 FreeSans 320 0 0 0 VOUT[2]
port 8 e
flabel metal2 s 1946 1429 1946 1429 3 FreeSans 320 0 0 0 VOUT[3]
port 9 e
flabel metal1 s 676 -1772 676 -1772 3 FreeSans 320 0 0 0 VDD
port 10 e
flabel metal1 s 670 1373 670 1373 3 FreeSans 320 0 0 0 VDDH
port 11 e
flabel metal1 s 671 -1227 671 -1227 3 FreeSans 320 0 0 0 GND
port 12 e
<< end >>
