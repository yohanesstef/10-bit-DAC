magic
tech sky130A
magscale 1 2
timestamp 1750845438
<< nwell >>
rect -308 -802 308 802
<< mvpmos >>
rect -50 420 50 504
rect -50 171 50 255
rect -50 -78 50 6
rect -50 -327 50 -243
rect -50 -576 50 -492
<< mvpdiff >>
rect -108 492 -50 504
rect -108 432 -96 492
rect -62 432 -50 492
rect -108 420 -50 432
rect 50 492 108 504
rect 50 432 62 492
rect 96 432 108 492
rect 50 420 108 432
rect -108 243 -50 255
rect -108 183 -96 243
rect -62 183 -50 243
rect -108 171 -50 183
rect 50 243 108 255
rect 50 183 62 243
rect 96 183 108 243
rect 50 171 108 183
rect -108 -6 -50 6
rect -108 -66 -96 -6
rect -62 -66 -50 -6
rect -108 -78 -50 -66
rect 50 -6 108 6
rect 50 -66 62 -6
rect 96 -66 108 -6
rect 50 -78 108 -66
rect -108 -255 -50 -243
rect -108 -315 -96 -255
rect -62 -315 -50 -255
rect -108 -327 -50 -315
rect 50 -255 108 -243
rect 50 -315 62 -255
rect 96 -315 108 -255
rect 50 -327 108 -315
rect -108 -504 -50 -492
rect -108 -564 -96 -504
rect -62 -564 -50 -504
rect -108 -576 -50 -564
rect 50 -504 108 -492
rect 50 -564 62 -504
rect 96 -564 108 -504
rect 50 -576 108 -564
<< mvpdiffc >>
rect -96 432 -62 492
rect 62 432 96 492
rect -96 183 -62 243
rect 62 183 96 243
rect -96 -66 -62 -6
rect 62 -66 96 -6
rect -96 -315 -62 -255
rect 62 -315 96 -255
rect -96 -564 -62 -504
rect 62 -564 96 -504
<< mvnsubdiff >>
rect -242 724 242 736
rect -242 690 -134 724
rect 134 690 242 724
rect -242 678 242 690
rect -242 628 -184 678
rect -242 -628 -230 628
rect -196 -628 -184 628
rect 184 628 242 678
rect -242 -678 -184 -628
rect 184 -628 196 628
rect 230 -628 242 628
rect 184 -678 242 -628
rect -242 -690 242 -678
rect -242 -724 -134 -690
rect 134 -724 242 -690
rect -242 -736 242 -724
<< mvnsubdiffcont >>
rect -134 690 134 724
rect -230 -628 -196 628
rect 196 -628 230 628
rect -134 -724 134 -690
<< poly >>
rect -50 585 50 601
rect -50 551 -34 585
rect 34 551 50 585
rect -50 504 50 551
rect -50 394 50 420
rect -50 336 50 352
rect -50 302 -34 336
rect 34 302 50 336
rect -50 255 50 302
rect -50 145 50 171
rect -50 87 50 103
rect -50 53 -34 87
rect 34 53 50 87
rect -50 6 50 53
rect -50 -104 50 -78
rect -50 -162 50 -146
rect -50 -196 -34 -162
rect 34 -196 50 -162
rect -50 -243 50 -196
rect -50 -353 50 -327
rect -50 -411 50 -395
rect -50 -445 -34 -411
rect 34 -445 50 -411
rect -50 -492 50 -445
rect -50 -602 50 -576
<< polycont >>
rect -34 551 34 585
rect -34 302 34 336
rect -34 53 34 87
rect -34 -196 34 -162
rect -34 -445 34 -411
<< locali >>
rect -230 690 -134 724
rect 134 690 230 724
rect -230 628 -196 690
rect 196 628 230 690
rect -50 551 -34 585
rect 34 551 50 585
rect -96 492 -62 508
rect -96 416 -62 432
rect 62 492 96 508
rect 62 416 96 432
rect -50 302 -34 336
rect 34 302 50 336
rect -96 243 -62 259
rect -96 167 -62 183
rect 62 243 96 259
rect 62 167 96 183
rect -50 53 -34 87
rect 34 53 50 87
rect -96 -6 -62 10
rect -96 -82 -62 -66
rect 62 -6 96 10
rect 62 -82 96 -66
rect -50 -196 -34 -162
rect 34 -196 50 -162
rect -96 -255 -62 -239
rect -96 -331 -62 -315
rect 62 -255 96 -239
rect 62 -331 96 -315
rect -50 -445 -34 -411
rect 34 -445 50 -411
rect -96 -504 -62 -488
rect -96 -580 -62 -564
rect 62 -504 96 -488
rect 62 -580 96 -564
rect -230 -690 -196 -628
rect 196 -690 230 -628
rect -230 -724 -134 -690
rect 134 -724 230 -690
<< viali >>
rect -26 551 26 585
rect -96 432 -62 492
rect 62 432 96 492
rect -26 302 26 336
rect -96 183 -62 243
rect 62 183 96 243
rect -26 53 26 87
rect -96 -66 -62 -6
rect 62 -66 96 -6
rect -26 -196 26 -162
rect -96 -315 -62 -255
rect 62 -315 96 -255
rect -26 -445 26 -411
rect -96 -564 -62 -504
rect 62 -564 96 -504
<< metal1 >>
rect -38 585 38 591
rect -38 551 -26 585
rect 26 551 38 585
rect -38 545 38 551
rect -102 492 -56 504
rect -102 432 -96 492
rect -62 432 -56 492
rect -102 420 -56 432
rect 56 492 102 504
rect 56 432 62 492
rect 96 432 102 492
rect 56 420 102 432
rect -38 336 38 342
rect -38 302 -26 336
rect 26 302 38 336
rect -38 296 38 302
rect -102 243 -56 255
rect -102 183 -96 243
rect -62 183 -56 243
rect -102 171 -56 183
rect 56 243 102 255
rect 56 183 62 243
rect 96 183 102 243
rect 56 171 102 183
rect -38 87 38 93
rect -38 53 -26 87
rect 26 53 38 87
rect -38 47 38 53
rect -102 -6 -56 6
rect -102 -66 -96 -6
rect -62 -66 -56 -6
rect -102 -78 -56 -66
rect 56 -6 102 6
rect 56 -66 62 -6
rect 96 -66 102 -6
rect 56 -78 102 -66
rect -38 -162 38 -156
rect -38 -196 -26 -162
rect 26 -196 38 -162
rect -38 -202 38 -196
rect -102 -255 -56 -243
rect -102 -315 -96 -255
rect -62 -315 -56 -255
rect -102 -327 -56 -315
rect 56 -255 102 -243
rect 56 -315 62 -255
rect 96 -315 102 -255
rect 56 -327 102 -315
rect -38 -411 38 -405
rect -38 -445 -26 -411
rect 26 -445 38 -411
rect -38 -451 38 -445
rect -102 -504 -56 -492
rect -102 -564 -96 -504
rect -62 -564 -56 -504
rect -102 -576 -56 -564
rect 56 -504 102 -492
rect 56 -564 62 -504
rect 96 -564 102 -504
rect 56 -576 102 -564
<< properties >>
string FIXED_BBOX -213 -707 213 707
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 0.50 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
