magic
tech sky130A
magscale 1 2
timestamp 1750075212
<< metal1 >>
rect -54 -65 43 -5
tri 43 -65 103 -5 sw
rect -54 -185 -48 -125
rect 12 -185 18 -125
tri 18 -150 103 -65 ne
tri 103 -76 114 -65 sw
rect 103 -125 114 -76
tri 114 -125 163 -76 sw
rect 103 -150 169 -125
tri 103 -185 138 -150 ne
rect 138 -185 169 -150
rect 229 -185 235 -125
<< via1 >>
rect -48 -185 12 -125
rect 169 -185 229 -125
<< metal2 >>
tri 103 -40 138 -5 se
rect 138 -40 235 -5
tri 18 -125 103 -40 se
rect 103 -65 235 -40
tri 103 -125 163 -65 nw
rect -54 -185 -48 -125
rect 12 -185 43 -125
tri 43 -185 103 -125 nw
rect 163 -185 169 -125
rect 229 -185 235 -125
<< end >>
