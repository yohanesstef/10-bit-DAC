magic
tech sky130A
magscale 1 2
timestamp 1750148716
<< metal3 >>
rect 2838 164 3132 260
rect 3319 -2276 7463 -2260
rect 3319 -2340 3336 -2276
rect 3400 -2340 4348 -2276
rect 4412 -2340 5360 -2276
rect 5424 -2340 6372 -2276
rect 6436 -2340 7384 -2276
rect 7448 -2340 7463 -2276
rect 3319 -2356 7463 -2340
<< via3 >>
rect 3336 -2340 3400 -2276
rect 4348 -2340 4412 -2276
rect 5360 -2340 5424 -2276
rect 6372 -2340 6436 -2276
rect 7384 -2340 7448 -2276
<< metal4 >>
rect 1827 164 8474 260
rect 1827 -3340 1923 164
rect 2307 -3160 2403 -12
rect 2839 -2668 2935 -347
rect 3319 -2276 3415 -736
rect 3319 -2340 3336 -2276
rect 3400 -2340 3415 -2276
rect 3319 -2440 3415 -2340
rect 3851 -2668 3947 -347
rect 4331 -2276 4427 -736
rect 4331 -2340 4348 -2276
rect 4412 -2340 4427 -2276
rect 4331 -2440 4427 -2340
rect 4863 -2668 4959 -347
rect 5343 -2276 5439 -736
rect 5343 -2340 5360 -2276
rect 5424 -2340 5439 -2276
rect 5343 -2440 5439 -2340
rect 5875 -2668 5971 -347
rect 6355 -2276 6451 -736
rect 6355 -2340 6372 -2276
rect 6436 -2340 6451 -2276
rect 6355 -2440 6451 -2340
rect 6887 -2668 6983 -347
rect 7367 -2276 7463 -736
rect 7367 -2340 7384 -2276
rect 7448 -2340 7463 -2276
rect 7367 -2440 7463 -2340
rect 7899 -3340 7995 164
rect 8379 -3236 8475 -88
rect 1827 -3388 8475 -3340
rect 1875 -3436 8475 -3388
use sky130_fd_pr__cap_mim_m3_1_UWHR8Z  sky130_fd_pr__cap_mim_m3_1_UWHR8Z_0
timestamp 1750148716
transform 1 0 5057 0 1 -1588
box -3422 -2040 3422 2040
<< end >>
