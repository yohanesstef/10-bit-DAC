magic
tech sky130A
magscale 1 2
timestamp 1749652636
<< error_s >>
rect 1438 -1854 1496 -1848
rect 1622 -1854 1680 -1848
rect 1438 -1888 1450 -1854
rect 1622 -1888 1634 -1854
rect 1438 -1894 1496 -1888
rect 1622 -1894 1680 -1888
<< poly >>
rect 1500 -1838 1530 -1829
rect 1434 -1854 1530 -1838
rect 1434 -1888 1450 -1854
rect 1484 -1888 1530 -1854
rect 1434 -1904 1530 -1888
rect 1588 -1838 1618 -1829
rect 1588 -1854 1684 -1838
rect 1588 -1888 1634 -1854
rect 1668 -1888 1684 -1854
rect 1588 -1904 1684 -1888
<< polycont >>
rect 1450 -1888 1484 -1854
rect 1634 -1888 1668 -1854
<< locali >>
rect 1434 -1888 1450 -1854
rect 1484 -1888 1500 -1854
rect 1618 -1888 1634 -1854
rect 1668 -1888 1684 -1854
<< viali >>
rect 1450 -1888 1484 -1854
rect 1634 -1888 1668 -1854
<< metal1 >>
rect 1529 -1847 1589 -1403
rect 1438 -1854 1496 -1848
rect 1438 -1888 1450 -1854
rect 1484 -1888 1496 -1854
rect 1438 -1894 1496 -1888
rect 1622 -1854 1680 -1848
rect 1622 -1888 1634 -1854
rect 1668 -1888 1680 -1854
rect 1622 -1894 1680 -1888
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_2
timestamp 1749643209
transform 1 0 1515 0 1 -1603
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_3
timestamp 1749643209
transform 1 0 1603 0 1 -1603
box -73 -226 73 226
<< end >>
