magic
tech sky130A
timestamp 1746772676
<< checkpaint >>
rect -649 -298 787 -274
rect -649 -322 944 -298
rect -649 -1854 1101 -322
rect -492 -1878 1101 -1854
rect -335 -1902 1101 -1878
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
use sky130_fd_sc_hd__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 0 0 1 -1200
box -19 -24 157 296
use sky130_fd_sc_hd__nand2_1  x2
timestamp 1704896540
transform 1 0 314 0 1 -1248
box -19 -24 157 296
use sky130_fd_sc_hd__nor2_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 157 0 1 -1224
box -19 -24 157 296
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 {bb\[6\]}
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 {bb\[7\]}
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 {bb\[8\]}
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 {bb\[9\]}
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 S
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 VDD
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 128 0 0 0 GND
port 6 nsew
<< end >>
