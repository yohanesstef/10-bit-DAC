magic
tech sky130A
magscale 1 2
timestamp 1750900893
<< error_p >>
rect 1105 -1290 1111 -1284
rect 1171 -1290 1177 -1284
rect 1409 -1290 1415 -1284
rect 1475 -1290 1481 -1284
rect 1111 -1296 1117 -1290
rect 1165 -1296 1171 -1290
rect 1415 -1296 1421 -1290
rect 1469 -1296 1475 -1290
rect 835 -1318 841 -1312
rect 889 -1318 895 -1312
rect 829 -1324 835 -1318
rect 895 -1324 901 -1318
rect 829 -1378 835 -1372
rect 895 -1378 901 -1372
rect 835 -1384 841 -1378
rect 889 -1384 895 -1378
rect 559 -1406 565 -1400
rect 613 -1406 619 -1400
rect 553 -1412 559 -1406
rect 619 -1412 625 -1406
rect 553 -1466 559 -1460
rect 619 -1466 625 -1460
rect 559 -1472 565 -1466
rect 613 -1472 619 -1466
rect 283 -1494 289 -1488
rect 337 -1494 343 -1488
rect 277 -1500 283 -1494
rect 343 -1500 349 -1494
rect 277 -1554 283 -1548
rect 343 -1554 349 -1548
rect 283 -1560 289 -1554
rect 337 -1560 343 -1554
rect 7 -1582 13 -1576
rect 61 -1582 67 -1576
rect 1 -1588 7 -1582
rect 67 -1588 73 -1582
rect 1 -1642 7 -1636
rect 67 -1642 73 -1636
rect 7 -1648 13 -1642
rect 61 -1648 67 -1642
<< error_s >>
rect 5335 -174 5341 -168
rect 5389 -174 5395 -168
rect 5329 -180 5335 -174
rect 5395 -180 5401 -174
rect 5329 -234 5335 -228
rect 5395 -234 5401 -228
rect 5335 -240 5341 -234
rect 5389 -240 5395 -234
rect 5059 -262 5065 -256
rect 5113 -262 5119 -256
rect 5053 -268 5059 -262
rect 5119 -268 5125 -262
rect 5053 -322 5059 -316
rect 5119 -322 5125 -316
rect 5059 -328 5065 -322
rect 5113 -328 5119 -322
rect 4783 -350 4789 -344
rect 4837 -350 4843 -344
rect 4777 -356 4783 -350
rect 4843 -356 4849 -350
rect 4777 -410 4783 -404
rect 4843 -410 4849 -404
rect 4783 -416 4789 -410
rect 4837 -416 4843 -410
rect 4507 -438 4513 -432
rect 4561 -438 4567 -432
rect 4501 -444 4507 -438
rect 4567 -444 4573 -438
rect 4501 -498 4507 -492
rect 4567 -498 4573 -492
rect 4507 -504 4513 -498
rect 4561 -504 4567 -498
rect 3927 -526 3933 -520
rect 3981 -526 3987 -520
rect 4231 -526 4237 -520
rect 4285 -526 4291 -520
rect 3921 -532 3927 -526
rect 3987 -532 3993 -526
rect 4225 -532 4231 -526
rect 4291 -532 4297 -526
rect 3921 -586 3927 -580
rect 3987 -586 3993 -580
rect 4225 -586 4231 -580
rect 4291 -586 4297 -580
rect 3927 -592 3933 -586
rect 3981 -592 3987 -586
rect 4231 -592 4237 -586
rect 4285 -592 4291 -586
rect 3651 -614 3657 -608
rect 3705 -614 3711 -608
rect 3645 -620 3651 -614
rect 3711 -620 3717 -614
rect 3645 -674 3651 -668
rect 3711 -674 3717 -668
rect 3651 -680 3657 -674
rect 3705 -680 3711 -674
rect 3375 -702 3381 -696
rect 3429 -702 3435 -696
rect 3369 -708 3375 -702
rect 3435 -708 3441 -702
rect 3369 -762 3375 -756
rect 3435 -762 3441 -756
rect 3375 -768 3381 -762
rect 3429 -768 3435 -762
rect 3099 -790 3105 -784
rect 3153 -790 3159 -784
rect 3093 -796 3099 -790
rect 3159 -796 3165 -790
rect 3093 -850 3099 -844
rect 3159 -850 3165 -844
rect 3099 -856 3105 -850
rect 3153 -856 3159 -850
rect 2519 -878 2525 -872
rect 2573 -878 2579 -872
rect 2823 -878 2829 -872
rect 2877 -878 2883 -872
rect 2513 -884 2519 -878
rect 2579 -884 2585 -878
rect 2817 -884 2823 -878
rect 2883 -884 2889 -878
rect 2513 -938 2519 -932
rect 2579 -938 2585 -932
rect 2817 -938 2823 -932
rect 2883 -938 2889 -932
rect 2519 -944 2525 -938
rect 2573 -944 2579 -938
rect 2823 -944 2829 -938
rect 2877 -944 2883 -938
rect 2243 -966 2249 -960
rect 2297 -966 2303 -960
rect 2237 -972 2243 -966
rect 2303 -972 2309 -966
rect 2237 -1026 2243 -1020
rect 2303 -1026 2309 -1020
rect 2243 -1032 2249 -1026
rect 2297 -1032 2303 -1026
rect 1967 -1054 1973 -1048
rect 2021 -1054 2027 -1048
rect 1961 -1060 1967 -1054
rect 2027 -1060 2033 -1054
rect 1961 -1114 1967 -1108
rect 2027 -1114 2033 -1108
rect 1967 -1120 1973 -1114
rect 2021 -1120 2027 -1114
rect 1691 -1142 1697 -1136
rect 1745 -1142 1751 -1136
rect 1685 -1148 1691 -1142
rect 1751 -1148 1757 -1142
rect 1685 -1202 1691 -1196
rect 1751 -1202 1757 -1196
rect 1691 -1208 1697 -1202
rect 1745 -1208 1751 -1202
rect 1111 -1230 1117 -1224
rect 1165 -1230 1171 -1224
rect 1415 -1230 1421 -1224
rect 1469 -1230 1475 -1224
rect 1105 -1236 1111 -1230
rect 1171 -1236 1177 -1230
rect 1409 -1236 1415 -1230
rect 1475 -1236 1481 -1230
<< pwell >>
rect -162 -166 5722 372
<< mvpsubdiff >>
rect -126 324 5686 336
rect -126 290 -18 324
rect 5578 290 5686 324
rect -126 278 5686 290
rect -126 228 -68 278
rect -126 -22 -114 228
rect -80 -22 -68 228
rect -126 -72 -68 -22
rect 5628 228 5686 278
rect 5628 -22 5640 228
rect 5674 -22 5686 228
rect 5628 -72 5686 -22
rect -126 -84 5686 -72
rect -126 -118 -18 -84
rect 5578 -118 5686 -84
rect -126 -130 5686 -118
<< mvpsubdiffcont >>
rect -18 290 5578 324
rect -114 -22 -80 228
rect 5640 -22 5674 228
rect -18 -118 5578 -84
<< locali >>
rect -114 290 -18 324
rect 5578 290 5674 324
rect -114 228 -80 290
rect -114 -84 -80 -22
rect 5640 228 5674 290
rect 5640 -84 5674 -22
rect -114 -118 -18 -84
rect 5578 -118 5674 -84
<< metal1 >>
rect 1294 811 1354 817
rect 1018 723 1078 729
rect 742 635 802 641
rect 466 547 526 553
rect 190 459 250 465
rect 7 -1582 67 114
rect 190 30 250 399
rect 283 -1494 343 114
rect 466 30 526 487
rect 559 -1406 619 114
rect 742 30 802 575
rect 835 -1318 895 114
rect 1018 30 1078 663
rect 1111 -1230 1171 114
rect 1294 30 1354 751
rect 2702 811 2762 817
rect 2426 723 2486 729
rect 2150 635 2210 641
rect 1874 547 1934 553
rect 1598 459 1658 465
rect 1111 -1296 1171 -1290
rect 1415 -1230 1475 114
rect 1598 30 1658 399
rect 1691 -1142 1751 114
rect 1874 30 1934 487
rect 1967 -1054 2027 114
rect 2150 30 2210 575
rect 2243 -966 2303 114
rect 2426 30 2486 663
rect 2519 -878 2579 114
rect 2702 30 2762 751
rect 4110 811 4170 817
rect 3834 723 3894 729
rect 3558 635 3618 641
rect 3282 547 3342 553
rect 3006 459 3066 465
rect 2519 -944 2579 -938
rect 2823 -878 2883 114
rect 3006 30 3066 399
rect 3099 -790 3159 114
rect 3282 30 3342 487
rect 3375 -702 3435 114
rect 3558 30 3618 575
rect 3651 -614 3711 114
rect 3834 30 3894 663
rect 3927 -526 3987 114
rect 4110 30 4170 751
rect 5518 811 5578 817
rect 5242 723 5302 729
rect 4966 635 5026 641
rect 4690 547 4750 553
rect 4414 459 4474 465
rect 3927 -592 3987 -586
rect 4231 -526 4291 114
rect 4414 30 4474 399
rect 4507 -438 4567 114
rect 4690 30 4750 487
rect 4783 -350 4843 114
rect 4966 30 5026 575
rect 5059 -262 5119 114
rect 5242 30 5302 663
rect 5335 -174 5395 114
rect 5518 30 5578 751
rect 5335 -240 5395 -234
rect 5059 -328 5119 -322
rect 4783 -416 4843 -410
rect 4507 -504 4567 -498
rect 4231 -592 4291 -586
rect 3651 -680 3711 -674
rect 3375 -768 3435 -762
rect 3099 -856 3159 -850
rect 2823 -944 2883 -938
rect 2243 -1032 2303 -1026
rect 1967 -1120 2027 -1114
rect 1691 -1208 1751 -1202
rect 1415 -1296 1475 -1290
rect 835 -1384 895 -1378
rect 559 -1472 619 -1466
rect 283 -1560 343 -1554
rect 7 -1648 67 -1642
<< via1 >>
rect 1294 751 1354 811
rect 1018 663 1078 723
rect 742 575 802 635
rect 466 487 526 547
rect 190 399 250 459
rect 2702 751 2762 811
rect 2426 663 2486 723
rect 2150 575 2210 635
rect 1874 487 1934 547
rect 1598 399 1658 459
rect 1111 -1290 1171 -1230
rect 4110 751 4170 811
rect 3834 663 3894 723
rect 3558 575 3618 635
rect 3282 487 3342 547
rect 3006 399 3066 459
rect 2519 -938 2579 -878
rect 5518 751 5578 811
rect 5242 663 5302 723
rect 4966 575 5026 635
rect 4690 487 4750 547
rect 4414 399 4474 459
rect 3927 -586 3987 -526
rect 5335 -234 5395 -174
rect 5059 -322 5119 -262
rect 4783 -410 4843 -350
rect 4507 -498 4567 -438
rect 4231 -586 4291 -526
rect 3651 -674 3711 -614
rect 3375 -762 3435 -702
rect 3099 -850 3159 -790
rect 2823 -938 2883 -878
rect 2243 -1026 2303 -966
rect 1967 -1114 2027 -1054
rect 1691 -1202 1751 -1142
rect 1415 -1290 1475 -1230
rect 835 -1378 895 -1318
rect 559 -1466 619 -1406
rect 283 -1554 343 -1494
rect 7 -1642 67 -1582
<< metal2 >>
rect 1288 751 1294 811
rect 1354 751 2702 811
rect 2762 751 4110 811
rect 4170 751 5518 811
rect 5578 751 5584 811
rect 1012 663 1018 723
rect 1078 663 2426 723
rect 2486 663 3834 723
rect 3894 663 5242 723
rect 5302 663 5308 723
rect 736 575 742 635
rect 802 575 2150 635
rect 2210 575 3558 635
rect 3618 575 4966 635
rect 5026 575 5032 635
rect 460 487 466 547
rect 526 487 1874 547
rect 1934 487 3282 547
rect 3342 487 4690 547
rect 4750 487 4756 547
rect 184 399 190 459
rect 250 399 1598 459
rect 1658 399 3006 459
rect 3066 399 4414 459
rect 4474 399 4480 459
use hnmos_1  hnmos_1_0
timestamp 1750900893
transform 1 0 2531 0 1 1
box -41 3 235 201
use hnmos_1  hnmos_1_1
timestamp 1750900893
transform 1 0 1123 0 1 1
box -41 3 235 201
use hnmos_1  hnmos_1_2
timestamp 1750900893
transform 1 0 3939 0 1 1
box -41 3 235 201
use hnmos_1  hnmos_1_3
timestamp 1750900893
transform 1 0 5347 0 1 1
box -41 3 235 201
use hnmos_4  hnmos_4_0
timestamp 1750900893
transform 1 0 -14 0 1 4
box -8 0 1096 198
use hnmos_4  hnmos_4_1
timestamp 1750900893
transform 1 0 1394 0 1 4
box -8 0 1096 198
use hnmos_4  hnmos_4_2
timestamp 1750900893
transform 1 0 2802 0 1 4
box -8 0 1096 198
use hnmos_4  hnmos_4_3
timestamp 1750900893
transform 1 0 4210 0 1 4
box -8 0 1096 198
<< end >>
