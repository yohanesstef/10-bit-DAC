* NGSPICE file created from top_segment_3.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_SEMVNL a_n141_n733# a_n141_301# VSUBS
X0 a_n141_301# a_n141_n733# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.17
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_SEMXNL a_n141_n733# a_n141_301# VSUBS
X0 a_n141_301# a_n141_n733# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.17
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_GLTCMD a_n141_311# a_n141_n743# VSUBS
X0 a_n141_311# a_n141_n743# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.27
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_42QADH a_n141_n748# a_n141_316# VSUBS
X0 a_n141_316# a_n141_n748# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.32
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_GVNVJY a_n141_n753# a_n141_321# VSUBS
X0 a_n141_321# a_n141_n753# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.37
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_AFTT8S a_n141_n769# a_n141_337# VSUBS
X0 a_n141_337# a_n141_n769# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.53
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_DZKNT5 a_n141_367# a_n141_n799# VSUBS
X0 a_n141_367# a_n141_n799# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.83
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_J5YLPL a_n141_n774# a_n141_342# VSUBS
X0 a_n141_342# a_n141_n774# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.58
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_47PAZ6 a_n141_n784# a_n141_352# VSUBS
X0 a_n141_352# a_n141_n784# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.68
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_DZKLT5 a_n141_367# a_n141_n799# VSUBS
X0 a_n141_367# a_n141_n799# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.83
.ends

.subckt rseg_3_1 sky130_fd_pr__res_xhigh_po_1p41_DZKNT5_0/a_n141_367# XR1/a_n141_n733#
+ sky130_fd_pr__res_xhigh_po_1p41_SEMVNL_0/a_n141_301# sky130_fd_pr__res_xhigh_po_1p41_DZKNT5_0/a_n141_n799#
+ m1_4812_n3449# m1_6357_n4745# sky130_fd_pr__res_xhigh_po_1p41_SEMVNL_0/a_n141_n733#
+ m1_6332_n4421# m1_4786_n4097# m1_6301_n2801# m1_6311_n3773# m1_4827_n2539# VSUBS
+ m1_4745_n4745#
Xsky130_fd_pr__res_xhigh_po_1p41_SEMVNL_0 sky130_fd_pr__res_xhigh_po_1p41_SEMVNL_0/a_n141_n733#
+ sky130_fd_pr__res_xhigh_po_1p41_SEMVNL_0/a_n141_301# VSUBS sky130_fd_pr__res_xhigh_po_1p41_SEMVNL
XXR1 XR1/a_n141_n733# m1_4827_n2539# VSUBS sky130_fd_pr__res_xhigh_po_1p41_SEMXNL
XXR2 m1_4827_n2539# m1_6301_n2801# VSUBS sky130_fd_pr__res_xhigh_po_1p41_GLTCMD
XXR3 m1_6301_n2801# m1_4812_n3449# VSUBS sky130_fd_pr__res_xhigh_po_1p41_42QADH
XXR4 m1_6311_n3773# m1_4812_n3449# VSUBS sky130_fd_pr__res_xhigh_po_1p41_GVNVJY
XXR5 m1_6311_n3773# m1_4786_n4097# VSUBS sky130_fd_pr__res_xhigh_po_1p41_AFTT8S
Xsky130_fd_pr__res_xhigh_po_1p41_DZKNT5_0 sky130_fd_pr__res_xhigh_po_1p41_DZKNT5_0/a_n141_367#
+ sky130_fd_pr__res_xhigh_po_1p41_DZKNT5_0/a_n141_n799# VSUBS sky130_fd_pr__res_xhigh_po_1p41_DZKNT5
XXR6 m1_6332_n4421# m1_4786_n4097# VSUBS sky130_fd_pr__res_xhigh_po_1p41_J5YLPL
XXR7 m1_6332_n4421# m1_4745_n4745# VSUBS sky130_fd_pr__res_xhigh_po_1p41_47PAZ6
XXR8 m1_4745_n4745# m1_6357_n4745# VSUBS sky130_fd_pr__res_xhigh_po_1p41_DZKLT5
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_QX57C3 a_n141_n825# a_n141_393# VSUBS
X0 a_n141_393# a_n141_n825# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=4.09
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_H2U5BC a_n141_n835# a_n141_403# VSUBS
X0 a_n141_403# a_n141_n835# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=4.19
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_E2U9YT a_n141_n861# a_n141_429# VSUBS
X0 a_n141_429# a_n141_n861# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=4.45
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_YY58WS a_n141_378# a_n141_n810# VSUBS
X0 a_n141_378# a_n141_n810# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.94
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_KLD4QF a_n141_n902# a_n141_470# VSUBS
X0 a_n141_470# a_n141_n902# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=4.86
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_4F76E7 a_n141_n876# a_n141_444# VSUBS
X0 a_n141_444# a_n141_n876# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=4.6
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_HDPFLR a_n141_n928# a_n141_496# VSUBS
X0 a_n141_496# a_n141_n928# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=5.12
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_5X53DF a_n141_526# a_n141_n958# VSUBS
X0 a_n141_526# a_n141_n958# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=5.42
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_YY56WS a_n141_378# a_n141_n810# VSUBS
X0 a_n141_378# a_n141_n810# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=3.94
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF a_n141_526# a_n141_n958# VSUBS
X0 a_n141_526# a_n141_n958# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=5.42
.ends

.subckt rseg_3_2 XR9/a_n141_n810# m1_8330_n3320# sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF_0/a_n141_526#
+ XR16/a_n141_n958# sky130_fd_pr__res_xhigh_po_1p41_YY58WS_0/a_n141_n810# m1_8304_n3968#
+ sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF_0/a_n141_n958# m1_10152_n3644# m1_8375_n2410#
+ m1_10116_n4292# m1_10193_n2996# m1_8263_n4616# sky130_fd_pr__res_xhigh_po_1p41_YY58WS_0/a_n141_378#
+ VSUBS
XXR10 m1_10116_n4292# m1_8263_n4616# VSUBS sky130_fd_pr__res_xhigh_po_1p41_QX57C3
XXR11 m1_10116_n4292# m1_8304_n3968# VSUBS sky130_fd_pr__res_xhigh_po_1p41_H2U5BC
XXR12 m1_10152_n3644# m1_8304_n3968# VSUBS sky130_fd_pr__res_xhigh_po_1p41_E2U9YT
Xsky130_fd_pr__res_xhigh_po_1p41_YY58WS_0 sky130_fd_pr__res_xhigh_po_1p41_YY58WS_0/a_n141_378#
+ sky130_fd_pr__res_xhigh_po_1p41_YY58WS_0/a_n141_n810# VSUBS sky130_fd_pr__res_xhigh_po_1p41_YY58WS
XXR14 m1_10193_n2996# m1_8330_n3320# VSUBS sky130_fd_pr__res_xhigh_po_1p41_KLD4QF
XXR13 m1_10152_n3644# m1_8330_n3320# VSUBS sky130_fd_pr__res_xhigh_po_1p41_4F76E7
XXR15 m1_10193_n2996# m1_8375_n2410# VSUBS sky130_fd_pr__res_xhigh_po_1p41_HDPFLR
XXR16 m1_8375_n2410# XR16/a_n141_n958# VSUBS sky130_fd_pr__res_xhigh_po_1p41_5X53DF
XXR9 m1_8263_n4616# XR9/a_n141_n810# VSUBS sky130_fd_pr__res_xhigh_po_1p41_YY56WS
Xsky130_fd_pr__res_xhigh_po_1p41_5X5ZCF_0 sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF_0/a_n141_526#
+ sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF_0/a_n141_n958# VSUBS sky130_fd_pr__res_xhigh_po_1p41_5X5ZCF
.ends

.subckt rseg_3_v3 v0 v1 v2 v4 v5 v6 v7 v8 v9 v11 v13 v15 gnd v16 v14 v10 v3 v12
Xrseg_3_1_0 gnd v0 gnd gnd v3 v8 gnd v6 v5 v2 v4 v1 gnd v7 rseg_3_1
Xrseg_3_2_0 v8 v13 gnd v16 gnd v11 gnd v12 v15 v10 v14 v9 gnd gnd rseg_3_2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WJ97JY w_n144_n140# a_n50_n104# a_n108_n78# a_50_n78#
X0 a_50_n78# a_n50_n104# a_n108_n78# w_n144_n140# sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
.ends

.subckt hpmos_1 XM1/a_50_n78# XM1/w_n144_n140# XM1/a_n108_n78# m1_1998_n3033#
XXM1 XM1/w_n144_n140# m1_1998_n3033# XM1/a_n108_n78# XM1/a_50_n78# sky130_fd_pr__pfet_g5v0d10v5_WJ97JY
.ends

.subckt hpmos_2 hpmos_1_1/XM1/a_n108_n78# hpmos_1_1/XM1/a_50_n78# hpmos_1_0/XM1/a_n108_n78#
+ hpmos_1_1/m1_1998_n3033# hpmos_1_0/XM1/a_50_n78# hpmos_1_1/XM1/w_n144_n140#
Xhpmos_1_0 hpmos_1_0/XM1/a_50_n78# hpmos_1_1/XM1/w_n144_n140# hpmos_1_0/XM1/a_n108_n78#
+ hpmos_1_1/m1_1998_n3033# hpmos_1
Xhpmos_1_1 hpmos_1_1/XM1/a_50_n78# hpmos_1_1/XM1/w_n144_n140# hpmos_1_1/XM1/a_n108_n78#
+ hpmos_1_1/m1_1998_n3033# hpmos_1
.ends

.subckt hpmos_4 hpmos_2_0/hpmos_1_0/XM1/a_50_n78# hpmos_2_0/hpmos_1_0/XM1/a_n108_n78#
+ hpmos_2_1/hpmos_1_1/XM1/a_n108_n78# hpmos_2_1/hpmos_1_0/XM1/a_50_n78# hpmos_2_1/hpmos_1_1/XM1/w_n144_n140#
+ hpmos_2_1/hpmos_1_0/XM1/a_n108_n78# hpmos_2_0/hpmos_1_1/XM1/a_50_n78# hpmos_2_1/hpmos_1_1/XM1/a_50_n78#
+ hpmos_2_0/hpmos_1_1/XM1/a_n108_n78# hpmos_2_1/hpmos_1_1/m1_1998_n3033#
Xhpmos_2_0 hpmos_2_0/hpmos_1_1/XM1/a_n108_n78# hpmos_2_0/hpmos_1_1/XM1/a_50_n78# hpmos_2_0/hpmos_1_0/XM1/a_n108_n78#
+ hpmos_2_1/hpmos_1_1/m1_1998_n3033# hpmos_2_0/hpmos_1_0/XM1/a_50_n78# hpmos_2_1/hpmos_1_1/XM1/w_n144_n140#
+ hpmos_2
Xhpmos_2_1 hpmos_2_1/hpmos_1_1/XM1/a_n108_n78# hpmos_2_1/hpmos_1_1/XM1/a_50_n78# hpmos_2_1/hpmos_1_0/XM1/a_n108_n78#
+ hpmos_2_1/hpmos_1_1/m1_1998_n3033# hpmos_2_1/hpmos_1_0/XM1/a_50_n78# hpmos_2_1/hpmos_1_1/XM1/w_n144_n140#
+ hpmos_2
.ends

.subckt hpmos_5 m1_292_56# m1_568_56# hpmos_4_0/hpmos_2_0/hpmos_1_0/XM1/a_50_n78#
+ hpmos_1_1/XM1/a_50_n78# m1_844_56# m1_16_56# hpmos_4_0/hpmos_2_1/hpmos_1_0/XM1/a_50_n78#
+ hpmos_4_0/hpmos_2_0/hpmos_1_1/XM1/a_50_n78# w_n156_n170# m1_1120_56# hpmos_4_0/hpmos_2_1/hpmos_1_1/XM1/a_50_n78#
+ hpmos_1_1/m1_1998_n3033#
Xhpmos_1_1 hpmos_1_1/XM1/a_50_n78# w_n156_n170# m1_1120_56# hpmos_1_1/m1_1998_n3033#
+ hpmos_1
Xhpmos_4_0 hpmos_4_0/hpmos_2_0/hpmos_1_0/XM1/a_50_n78# m1_16_56# m1_844_56# hpmos_4_0/hpmos_2_1/hpmos_1_0/XM1/a_50_n78#
+ w_n156_n170# m1_568_56# hpmos_4_0/hpmos_2_0/hpmos_1_1/XM1/a_50_n78# hpmos_4_0/hpmos_2_1/hpmos_1_1/XM1/a_50_n78#
+ m1_292_56# hpmos_1_1/m1_1998_n3033# hpmos_4
.ends

.subckt tps3_switch_10 hpmos_5_1/hpmos_1_1/m1_1998_n3033# hpmos_5_0/m1_844_56# hpmos_5_1/m1_844_56#
+ hpmos_5_1/m1_16_56# hpmos_5_1/hpmos_4_0/hpmos_2_0/hpmos_1_0/XM1/a_50_n78# hpmos_5_0/hpmos_1_1/XM1/a_50_n78#
+ hpmos_5_0/hpmos_4_0/hpmos_2_0/hpmos_1_0/XM1/a_50_n78# hpmos_5_1/w_n156_n170# hpmos_5_1/hpmos_4_0/hpmos_2_1/hpmos_1_0/XM1/a_50_n78#
+ hpmos_5_0/hpmos_4_0/hpmos_2_1/hpmos_1_0/XM1/a_50_n78# hpmos_5_1/hpmos_1_1/XM1/a_50_n78#
+ hpmos_5_0/hpmos_1_1/m1_1998_n3033# hpmos_5_0/m1_1120_56# hpmos_5_1/m1_1120_56# hpmos_5_1/hpmos_4_0/hpmos_2_0/hpmos_1_1/XM1/a_50_n78#
+ hpmos_5_0/hpmos_4_0/hpmos_2_0/hpmos_1_1/XM1/a_50_n78# hpmos_5_0/m1_292_56# hpmos_5_0/m1_568_56#
+ hpmos_5_1/m1_292_56# hpmos_5_1/m1_568_56# hpmos_5_1/hpmos_4_0/hpmos_2_1/hpmos_1_1/XM1/a_50_n78#
+ hpmos_5_0/hpmos_4_0/hpmos_2_1/hpmos_1_1/XM1/a_50_n78# hpmos_5_0/m1_16_56#
Xhpmos_5_0 hpmos_5_0/m1_292_56# hpmos_5_0/m1_568_56# hpmos_5_0/hpmos_4_0/hpmos_2_0/hpmos_1_0/XM1/a_50_n78#
+ hpmos_5_0/hpmos_1_1/XM1/a_50_n78# hpmos_5_0/m1_844_56# hpmos_5_0/m1_16_56# hpmos_5_0/hpmos_4_0/hpmos_2_1/hpmos_1_0/XM1/a_50_n78#
+ hpmos_5_0/hpmos_4_0/hpmos_2_0/hpmos_1_1/XM1/a_50_n78# hpmos_5_1/w_n156_n170# hpmos_5_0/m1_1120_56#
+ hpmos_5_0/hpmos_4_0/hpmos_2_1/hpmos_1_1/XM1/a_50_n78# hpmos_5_0/hpmos_1_1/m1_1998_n3033#
+ hpmos_5
Xhpmos_5_1 hpmos_5_1/m1_292_56# hpmos_5_1/m1_568_56# hpmos_5_1/hpmos_4_0/hpmos_2_0/hpmos_1_0/XM1/a_50_n78#
+ hpmos_5_1/hpmos_1_1/XM1/a_50_n78# hpmos_5_1/m1_844_56# hpmos_5_1/m1_16_56# hpmos_5_1/hpmos_4_0/hpmos_2_1/hpmos_1_0/XM1/a_50_n78#
+ hpmos_5_1/hpmos_4_0/hpmos_2_0/hpmos_1_1/XM1/a_50_n78# hpmos_5_1/w_n156_n170# hpmos_5_1/m1_1120_56#
+ hpmos_5_1/hpmos_4_0/hpmos_2_1/hpmos_1_1/XM1/a_50_n78# hpmos_5_1/hpmos_1_1/m1_1998_n3033#
+ hpmos_5
.ends

.subckt tps3_switch_final_stage hpmos_2_0/hpmos_1_0/XM1/a_50_n78# hpmos_1_1/XM1/a_n108_n78#
+ hpmos_2_0/hpmos_1_0/XM1/a_n108_n78# hpmos_1_1/XM1/a_50_n78# hpmos_2_3/hpmos_1_1/XM1/a_50_n78#
+ hpmos_1_0/m1_1998_n3033# hpmos_2_1/hpmos_1_1/XM1/a_n108_n78# hpmos_1_0/XM1/a_n108_n78#
+ hpmos_2_1/hpmos_1_0/XM1/a_50_n78# hpmos_2_0/hpmos_1_1/XM1/a_50_n78# hpmos_2_1/hpmos_1_0/XM1/a_n108_n78#
+ w_n1308_n166# hpmos_2_2/hpmos_1_1/m1_1998_n3033# hpmos_2_2/hpmos_1_1/XM1/a_n108_n78#
+ hpmos_2_2/hpmos_1_0/XM1/a_50_n78# hpmos_2_1/hpmos_1_1/XM1/a_50_n78# hpmos_2_2/hpmos_1_0/XM1/a_n108_n78#
+ hpmos_2_3/hpmos_1_1/m1_1998_n3033# hpmos_1_0/XM1/a_50_n78# hpmos_2_3/hpmos_1_1/XM1/a_n108_n78#
+ hpmos_2_3/hpmos_1_0/XM1/a_50_n78# hpmos_1_1/m1_1998_n3033# hpmos_2_2/hpmos_1_1/XM1/a_50_n78#
+ hpmos_2_0/hpmos_1_1/XM1/a_n108_n78# hpmos_2_3/hpmos_1_0/XM1/a_n108_n78#
Xhpmos_1_0 hpmos_1_0/XM1/a_50_n78# w_n1308_n166# hpmos_1_0/XM1/a_n108_n78# hpmos_1_0/m1_1998_n3033#
+ hpmos_1
Xhpmos_1_1 hpmos_1_1/XM1/a_50_n78# w_n1308_n166# hpmos_1_1/XM1/a_n108_n78# hpmos_1_1/m1_1998_n3033#
+ hpmos_1
Xhpmos_2_0 hpmos_2_0/hpmos_1_1/XM1/a_n108_n78# hpmos_2_0/hpmos_1_1/XM1/a_50_n78# hpmos_2_0/hpmos_1_0/XM1/a_n108_n78#
+ hpmos_1_1/m1_1998_n3033# hpmos_2_0/hpmos_1_0/XM1/a_50_n78# w_n1308_n166# hpmos_2
Xhpmos_2_1 hpmos_2_1/hpmos_1_1/XM1/a_n108_n78# hpmos_2_1/hpmos_1_1/XM1/a_50_n78# hpmos_2_1/hpmos_1_0/XM1/a_n108_n78#
+ hpmos_1_0/m1_1998_n3033# hpmos_2_1/hpmos_1_0/XM1/a_50_n78# w_n1308_n166# hpmos_2
Xhpmos_2_2 hpmos_2_2/hpmos_1_1/XM1/a_n108_n78# hpmos_2_2/hpmos_1_1/XM1/a_50_n78# hpmos_2_2/hpmos_1_0/XM1/a_n108_n78#
+ hpmos_2_2/hpmos_1_1/m1_1998_n3033# hpmos_2_2/hpmos_1_0/XM1/a_50_n78# w_n1308_n166#
+ hpmos_2
Xhpmos_2_3 hpmos_2_3/hpmos_1_1/XM1/a_n108_n78# hpmos_2_3/hpmos_1_1/XM1/a_50_n78# hpmos_2_3/hpmos_1_0/XM1/a_n108_n78#
+ hpmos_2_3/hpmos_1_1/m1_1998_n3033# hpmos_2_3/hpmos_1_0/XM1/a_50_n78# w_n1308_n166#
+ hpmos_2
.ends

.subckt hpmos_9 hpmos_4_1/hpmos_2_0/hpmos_1_0/XM1/a_50_n78# hpmos_4_0/hpmos_2_0/hpmos_1_0/XM1/a_50_n78#
+ m1_4315_962# hpmos_1_1/XM1/a_50_n78# m1_2452_962# hpmos_4_1/hpmos_2_1/hpmos_1_0/XM1/a_50_n78#
+ hpmos_4_0/hpmos_2_1/hpmos_1_0/XM1/a_50_n78# hpmos_4_1/hpmos_2_0/hpmos_1_1/XM1/a_50_n78#
+ m1_2659_962# hpmos_4_0/hpmos_2_0/hpmos_1_1/XM1/a_50_n78# m1_3487_962# m1_2935_962#
+ hpmos_4_1/hpmos_2_1/hpmos_1_1/XM1/a_50_n78# m1_3763_962# hpmos_4_0/hpmos_2_1/hpmos_1_1/XM1/a_50_n78#
+ m1_3211_962# m1_4591_962# hpmos_1_1/m1_1998_n3033# w_2208_736# m1_4039_962#
Xhpmos_1_1 hpmos_1_1/XM1/a_50_n78# w_2208_736# m1_4591_962# hpmos_1_1/m1_1998_n3033#
+ hpmos_1
Xhpmos_4_0 hpmos_4_0/hpmos_2_0/hpmos_1_0/XM1/a_50_n78# m1_2452_962# m1_3211_962# hpmos_4_0/hpmos_2_1/hpmos_1_0/XM1/a_50_n78#
+ w_2208_736# m1_2935_962# hpmos_4_0/hpmos_2_0/hpmos_1_1/XM1/a_50_n78# hpmos_4_0/hpmos_2_1/hpmos_1_1/XM1/a_50_n78#
+ m1_2659_962# hpmos_1_1/m1_1998_n3033# hpmos_4
Xhpmos_4_1 hpmos_4_1/hpmos_2_0/hpmos_1_0/XM1/a_50_n78# m1_3487_962# m1_4315_962# hpmos_4_1/hpmos_2_1/hpmos_1_0/XM1/a_50_n78#
+ w_2208_736# m1_4039_962# hpmos_4_1/hpmos_2_0/hpmos_1_1/XM1/a_50_n78# hpmos_4_1/hpmos_2_1/hpmos_1_1/XM1/a_50_n78#
+ m1_3763_962# hpmos_1_1/m1_1998_n3033# hpmos_4
.ends

.subckt top_segment_3 V0 V16 b[3] b[4] b[5] b[6] bb[3] bb[4] bb[5] bb[6] VH VL GND
+ VPB
Xrseg_3_v3_0 V0 rseg_3_v3_0/v1 rseg_3_v3_0/v2 rseg_3_v3_0/v4 rseg_3_v3_0/v5 rseg_3_v3_0/v6
+ rseg_3_v3_0/v7 rseg_3_v3_0/v8 rseg_3_v3_0/v9 rseg_3_v3_0/v11 rseg_3_v3_0/v13 rseg_3_v3_0/v15
+ GND V16 rseg_3_v3_0/v14 rseg_3_v3_0/v10 rseg_3_v3_0/v3 rseg_3_v3_0/v12 rseg_3_v3
Xtps3_switch_10_0 bb[5] m1_6825_5928# m1_6825_5928# m1_7957_5928# m1_9455_5394# m1_9455_5394#
+ m1_8351_5042# VPB m1_10275_5570# m1_8903_5218# m1_9723_5746# b[5] m1_6549_5928#
+ m1_6549_5928# m1_10551_5482# m1_8627_5130# m1_7681_5928# m1_7101_5928# m1_7681_5928#
+ m1_7101_5928# m1_9999_5658# m1_9179_5306# m1_7957_5928# tps3_switch_10
Xtps3_switch_final_stage_0 m1_6549_5928# m1_6245_5928# m1_5389_5928# m1_7101_5928#
+ m1_5665_5928# b[4] m1_5665_5928# m1_6245_5928# m1_7101_5928# m1_6825_5928# m1_5389_5928#
+ VPB b[3] VL m1_5665_5928# m1_7681_5928# VH bb[3] m1_7957_5928# VL m1_5389_5928#
+ bb[4] m1_6245_5928# m1_5665_5928# VH tps3_switch_final_stage
Xhpmos_9_0 rseg_3_v3_0/v4 V0 m1_9999_5658# rseg_3_v3_0/v8 m1_8351_5042# rseg_3_v3_0/v6
+ rseg_3_v3_0/v2 rseg_3_v3_0/v5 m1_8627_5130# rseg_3_v3_0/v1 m1_9455_5394# m1_8903_5218#
+ rseg_3_v3_0/v7 m1_10551_5482# rseg_3_v3_0/v3 m1_9179_5306# m1_9723_5746# bb[6] VPB
+ m1_10275_5570# hpmos_9
Xhpmos_9_1 rseg_3_v3_0/v12 rseg_3_v3_0/v8 m1_9999_5658# V16 m1_8351_5042# rseg_3_v3_0/v14
+ rseg_3_v3_0/v10 rseg_3_v3_0/v13 m1_8627_5130# rseg_3_v3_0/v9 m1_9455_5394# m1_8903_5218#
+ rseg_3_v3_0/v15 m1_10551_5482# rseg_3_v3_0/v11 m1_9179_5306# m1_9723_5746# b[6]
+ VPB m1_10275_5570# hpmos_9
.ends

