magic
tech sky130A
magscale 1 2
timestamp 1749630286
<< pwell >>
rect 10163 -19548 24372 -15966
<< psubdiff >>
rect 10199 -16062 10459 -16002
rect 24076 -16062 24336 -16002
rect 10199 -16262 10259 -16062
rect 10199 -19452 10259 -19252
rect 24276 -16262 24336 -16062
rect 24276 -19452 24336 -19252
rect 10199 -19512 10459 -19452
rect 24076 -19512 24336 -19452
<< psubdiffcont >>
rect 10459 -16062 24076 -16002
rect 10199 -19252 10259 -16262
rect 24276 -19252 24336 -16262
rect 10459 -19512 24076 -19452
<< locali >>
rect 10199 -16062 10459 -16002
rect 24076 -16062 24336 -16002
rect 10199 -16262 10259 -16062
rect 10613 -16158 11045 -16062
rect 11985 -16158 12417 -16062
rect 13054 -16158 13486 -16062
rect 13790 -16158 14222 -16062
rect 14766 -16158 15198 -16062
rect 15482 -16158 15914 -16062
rect 16546 -16158 16978 -16062
rect 17160 -16158 17592 -16062
rect 18136 -16158 18568 -16062
rect 18740 -16158 19172 -16062
rect 19809 -16158 20241 -16062
rect 20361 -16158 20793 -16062
rect 21337 -16158 21769 -16062
rect 21899 -16158 22331 -16062
rect 22968 -16158 23400 -16062
rect 23490 -16158 23922 -16062
rect 10199 -19452 10259 -19252
rect 24276 -16262 24336 -16062
rect 10849 -19452 11281 -19356
rect 11749 -19452 12181 -19356
rect 12987 -19452 13419 -19356
rect 13857 -19452 14289 -19356
rect 14792 -19452 15224 -19356
rect 15456 -19452 15888 -19356
rect 16531 -19452 16963 -19356
rect 17175 -19452 17607 -19356
rect 18152 -19452 18584 -19356
rect 18724 -19452 19156 -19356
rect 19794 -19452 20226 -19356
rect 20376 -19452 20808 -19356
rect 21347 -19452 21779 -19356
rect 21889 -19452 22321 -19356
rect 22958 -19452 23390 -19356
rect 23500 -19452 23932 -19356
rect 24276 -19452 24336 -19252
rect 10199 -19512 10459 -19452
rect 24076 -19512 24336 -19452
<< metal1 >>
rect 12763 -19022 12769 -18760
<< via1 >>
rect 12345 -16754 12405 -16492
rect 14150 -16754 14210 -16492
rect 15842 -16754 15902 -16492
rect 17520 -16754 17580 -16492
rect 19100 -16754 19160 -16492
rect 20721 -16754 20781 -16492
rect 22259 -16754 22319 -16492
rect 23849 -16754 23909 -16492
rect 12703 -19022 12763 -18760
rect 14217 -19022 14277 -18760
rect 16194 -19022 16254 -18760
rect 17535 -19022 17595 -18760
rect 19452 -19022 19512 -18760
rect 20736 -19022 20796 -18760
rect 22611 -19022 22671 -18760
rect 23860 -19022 23920 -18760
<< metal2 >>
rect 11487 -16024 12186 -15964
rect 15638 -16024 15689 -15964
rect 13924 -16112 14059 -16052
rect 17413 -16112 17440 -16052
rect 11487 -16200 12186 -16140
rect 13924 -16200 14059 -16140
rect 15637 -16200 15688 -16140
rect 17417 -16200 17444 -16140
rect 13923 -16288 14058 -16228
rect 17416 -16288 17443 -16228
rect 11487 -16376 12186 -16316
rect 15638 -16376 15689 -16316
rect 10163 -16754 12345 -16492
rect 12405 -16754 12411 -16492
rect 14144 -16754 14150 -16492
rect 14210 -16754 15842 -16492
rect 15902 -16754 15908 -16492
rect 17514 -16754 17520 -16492
rect 17580 -16754 19100 -16492
rect 19160 -16754 19166 -16492
rect 20715 -16754 20721 -16492
rect 20781 -16754 22259 -16492
rect 22319 -16754 22325 -16492
rect 23843 -16754 23849 -16492
rect 23909 -16754 24372 -16492
rect 12697 -19022 12703 -18760
rect 12763 -19022 14217 -18760
rect 14277 -19022 14283 -18760
rect 16188 -19022 16194 -18760
rect 16254 -19022 17535 -18760
rect 17595 -19022 17601 -18760
rect 19446 -19022 19452 -18760
rect 19512 -19022 20736 -18760
rect 20796 -19022 20802 -18760
rect 22604 -19022 22611 -18760
rect 22671 -19022 23860 -18760
rect 23920 -19022 23926 -18760
use pin_8_even  pin_8_even_0
timestamp 1749382758
transform 1 0 11128 0 1 -19447
box 1569 2955 2796 3659
use pin_8_even  pin_8_even_1
timestamp 1749382758
transform 1 0 17883 0 1 -19447
box 1569 2955 2796 3659
use pin_8_even  pin_8_even_2
timestamp 1749382758
transform 1 0 14625 0 1 -19447
box 1569 2955 2796 3659
use pin_8_even  pin_8_even_3
timestamp 1749382758
transform 1 0 21042 0 1 -19447
box 1569 2955 2796 3659
use pin_8_even_rigth  pin_8_even_rigth_0
timestamp 1749382774
transform 1 0 14707 0 1 -19447
box 2721 2955 3149 3401
use pin_8_even_rigth  pin_8_even_rigth_1
timestamp 1749382774
transform 1 0 17908 0 1 -19447
box 2721 2955 3149 3401
use pin_8_even_rigth  pin_8_even_rigth_2
timestamp 1749382774
transform 1 0 21037 0 1 -19447
box 2721 2955 3149 3401
use pin_8_even_rigth  pin_8_even_rigth_3
timestamp 1749382774
transform 1 0 11337 0 1 -19447
box 2721 2955 3149 3401
use pin_8_odd  pin_8_odd_0
timestamp 1749375316
transform 1 0 10266 0 1 -19447
box 83 2955 1221 3659
use pin_8_odd  pin_8_odd_1
timestamp 1749375316
transform 1 0 14419 0 1 -19447
box 83 2955 1221 3659
use pin_8_odd  pin_8_odd_2
timestamp 1749375316
transform 1 0 17789 0 1 -19447
box 83 2955 1221 3659
use pin_8_odd  pin_8_odd_3
timestamp 1749375316
transform 1 0 20990 0 1 -19447
box 83 2955 1221 3659
use pin_8_odd_right  pin_8_odd_right_0
timestamp 1749376058
transform 1 0 11128 0 1 -19447
box 1057 2955 1553 3489
use pin_8_odd_right  pin_8_odd_right_1
timestamp 1749376058
transform 1 0 14625 0 1 -19447
box 1057 2955 1553 3489
use pin_8_odd_right  pin_8_odd_right_2
timestamp 1749376058
transform 1 0 17883 0 1 -19447
box 1057 2955 1553 3489
use pin_8_odd_right  pin_8_odd_right_3
timestamp 1749376058
transform 1 0 21042 0 1 -19447
box 1057 2955 1553 3489
use rseg_1_1  rseg_1_1_1
timestamp 1749538868
transform 1 0 8815 0 1 6272
box 1540 -25628 3948 -22430
use rseg_1_2  rseg_1_2_1
timestamp 1749538868
transform 1 0 1523 0 1 4689
box 11268 -24045 12957 -20847
use rseg_1_3  rseg_1_3_0
timestamp 1749538868
transform 1 0 -191 0 1 4228
box 14699 -23584 16451 -20386
use rseg_1_4  rseg_1_4_0
timestamp 1749538868
transform 1 0 2239 0 1 4689
box 14049 -24045 15611 -20847
use rseg_1_5  rseg_1_5_0
timestamp 1749538868
transform 1 0 2701 0 1 4689
box 15177 -24045 16817 -20847
use rseg_1_6  rseg_1_6_0
timestamp 1749538868
transform 1 0 3240 0 1 4689
box 16306 -24045 17811 -20847
use rseg_1_7  rseg_1_7_0
timestamp 1749538868
transform 1 0 3721 0 1 4689
box 17358 -24045 18956 -20847
use rseg_1_8  rseg_1_8_0
timestamp 1749538868
transform 1 0 4243 0 1 4689
box 18462 -24045 19937 -20847
<< labels >>
flabel metal1 s 13060 -16492 13060 -16492 2 FreeSans 240 0 0 0 v15
port 15 ne
flabel metal1 s 23856 -16492 23856 -16492 2 FreeSans 240 0 0 0 v64
port 64 ne
flabel metal1 s 22969 -16492 22969 -16492 2 FreeSans 240 0 0 0 v63
port 63 ne
flabel metal1 s 23944 -16492 23944 -16492 2 FreeSans 240 0 0 0 v62
port 62 ne
flabel metal1 s 22881 -16492 22881 -16492 2 FreeSans 240 0 0 0 v61
port 61 ne
flabel metal1 s 24032 -16492 24032 -16492 2 FreeSans 240 0 0 0 v60
port 60 ne
flabel metal1 s 22793 -16492 22793 -16492 2 FreeSans 240 0 0 0 v59
port 59 ne
flabel metal1 s 24120 -16492 24120 -16492 2 FreeSans 240 0 0 0 v58
port 58 ne
flabel metal1 s 22705 -16492 22705 -16492 2 FreeSans 240 0 0 0 v57
port 57 ne
flabel metal1 s 22617 -16492 22617 -16492 2 FreeSans 240 0 0 0 v56
port 56 ne
flabel metal1 s 21079 -16492 21079 -16492 2 FreeSans 240 0 0 0 v55
port 55 ne
flabel metal1 s 22529 -16492 22529 -16492 2 FreeSans 240 0 0 0 v54
port 54 ne
flabel metal1 s 21167 -16492 21167 -16492 2 FreeSans 240 0 0 0 v53
port 53 ne
flabel metal1 s 22441 -16492 22441 -16492 2 FreeSans 240 0 0 0 v52
port 52 ne
flabel metal1 s 21255 -16492 21255 -16492 2 FreeSans 240 0 0 0 v51
port 51 ne
flabel metal1 s 22353 -16492 22353 -16492 2 FreeSans 240 0 0 0 v50
port 50 ne
flabel metal1 s 21343 -16492 21343 -16492 2 FreeSans 240 0 0 0 v49
port 49 ne
flabel metal1 s 20727 -16492 20727 -16492 2 FreeSans 240 0 0 0 v48
port 48 ne
flabel metal1 s 19810 -16492 19810 -16492 2 FreeSans 240 0 0 0 v47
port 47 ne
flabel metal1 s 20815 -16492 20815 -16492 2 FreeSans 240 0 0 0 v46
port 46 ne
flabel metal1 s 19722 -16492 19722 -16492 2 FreeSans 240 0 0 0 v45
port 45 ne
flabel metal1 s 20903 -16492 20903 -16492 2 FreeSans 240 0 0 0 v44
port 44 ne
flabel metal1 s 19634 -16492 19634 -16492 2 FreeSans 240 0 0 0 v43
port 43 ne
flabel metal1 s 20991 -16492 20991 -16492 2 FreeSans 240 0 0 0 v42
port 42 ne
flabel metal1 s 19546 -16492 19546 -16492 2 FreeSans 240 0 0 0 v41
port 41 ne
flabel metal1 s 19458 -16492 19458 -16492 2 FreeSans 240 0 0 0 v40
port 40 ne
flabel metal1 s 17878 -16492 17878 -16492 2 FreeSans 240 0 0 0 v39
port 39 ne
flabel metal1 s 19370 -16492 19370 -16492 2 FreeSans 240 0 0 0 v38
port 38 ne
flabel metal1 s 17966 -16492 17966 -16492 2 FreeSans 240 0 0 0 v37
port 37 ne
flabel metal1 s 19282 -16492 19282 -16492 2 FreeSans 240 0 0 0 v36
port 36 ne
flabel metal1 s 18054 -16493 18054 -16493 2 FreeSans 240 0 0 0 v35
port 35 ne
flabel metal1 s 19194 -16492 19194 -16492 2 FreeSans 240 0 0 0 v34
port 34 ne
flabel metal1 s 18142 -16492 18142 -16492 2 FreeSans 240 0 0 0 v33
port 33 ne
flabel metal1 s 17526 -16492 17526 -16492 2 FreeSans 240 0 0 0 v32
port 32 ne
flabel metal1 s 16552 -16492 16552 -16492 2 FreeSans 240 0 0 0 v31
port 31 ne
flabel metal1 s 17614 -16492 17614 -16492 2 FreeSans 240 0 0 0 v30
port 30 ne
flabel metal1 s 16464 -16492 16464 -16492 2 FreeSans 240 0 0 0 v29
port 29 ne
flabel metal1 s 17702 -16492 17702 -16492 2 FreeSans 240 0 0 0 v28
port 28 ne
flabel metal1 s 16376 -16492 16376 -16492 2 FreeSans 240 0 0 0 v27
port 27 ne
flabel metal1 s 17790 -16492 17790 -16492 2 FreeSans 240 0 0 0 v26
port 26 ne
flabel metal1 s 16288 -16492 16288 -16492 2 FreeSans 240 0 0 0 v25
port 25 ne
flabel metal1 s 16200 -16492 16200 -16492 2 FreeSans 240 0 0 0 v24
port 24 ne
flabel metal1 s 14508 -16492 14508 -16492 2 FreeSans 240 0 0 0 v23
port 23 ne
flabel metal1 s 16112 -16492 16112 -16492 2 FreeSans 240 0 0 0 v22
port 22 ne
flabel metal1 s 14596 -16492 14596 -16492 2 FreeSans 240 0 0 0 v21
port 21 ne
flabel metal1 s 16024 -16492 16024 -16492 2 FreeSans 240 0 0 0 v20
port 20 ne
flabel metal1 s 14684 -16492 14684 -16492 2 FreeSans 240 0 0 0 v19
port 19 ne
flabel metal1 s 15936 -16492 15936 -16492 2 FreeSans 240 0 0 0 v18
port 18 ne
flabel metal1 s 14772 -16492 14772 -16492 2 FreeSans 240 0 0 0 v17
port 17 ne
flabel metal1 s 14156 -16492 14156 -16492 2 FreeSans 240 0 0 0 v16
port 16 ne
flabel metal1 s 14244 -16492 14244 -16492 2 FreeSans 240 0 0 0 v14
port 14 ne
flabel metal1 s 12967 -16492 12967 -16492 2 FreeSans 240 0 0 0 v13
port 13 ne
flabel metal1 s 14332 -16492 14332 -16492 2 FreeSans 240 0 0 0 v12
port 12 ne
flabel metal1 s 12879 -16492 12879 -16492 2 FreeSans 240 0 0 0 v11
port 11 ne
flabel metal1 s 14420 -16492 14420 -16492 2 FreeSans 240 0 0 0 v10
port 10 ne
flabel metal1 s 12791 -16492 12791 -16492 2 FreeSans 240 0 0 0 v9
port 9 ne
flabel metal1 s 12703 -16492 12703 -16492 2 FreeSans 240 0 0 0 v8
port 8 ne
flabel metal1 s 10355 -16492 10355 -16492 2 FreeSans 240 0 0 0 v7
port 7 ne
flabel metal1 s 12615 -16492 12615 -16492 2 FreeSans 240 0 0 0 v6
port 6 ne
flabel metal1 s 10443 -16492 10443 -16492 2 FreeSans 240 0 0 0 v5
port 5 ne
flabel metal1 s 12527 -16492 12527 -16492 2 FreeSans 240 0 0 0 v4
port 4 ne
flabel metal1 s 12439 -16492 12439 -16492 2 FreeSans 240 0 0 0 v2
port 2 ne
flabel metal1 s 10531 -16492 10531 -16492 2 FreeSans 240 0 0 0 v3
port 3 ne
flabel metal1 s 10619 -16492 10619 -16492 2 FreeSans 240 0 0 0 v1
port 1 ne
flabel locali s 10199 -19512 10199 -19512 2 FreeSans 1600 0 0 0 gnd
port 65 ne
flabel metal2 s 10163 -16754 10163 -16754 2 FreeSans 1600 0 0 0 v0
port 0 ne
<< end >>
