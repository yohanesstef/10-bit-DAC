magic
tech sky130A
magscale 1 2
timestamp 1749147130
<< pwell >>
rect -307 -740 307 740
<< psubdiff >>
rect -271 670 -175 704
rect 175 670 271 704
rect -271 608 -237 670
rect 237 608 271 670
rect -271 -670 -237 -608
rect 237 -670 271 -608
rect -271 -704 -175 -670
rect 175 -704 271 -670
<< psubdiffcont >>
rect -175 670 175 704
rect -271 -608 -237 608
rect 237 -608 271 608
rect -175 -704 175 -670
<< xpolycontact >>
rect -141 142 141 574
rect -141 -574 141 -142
<< xpolyres >>
rect -141 -142 141 142
<< locali >>
rect -271 670 -175 704
rect 175 670 271 704
rect -271 608 -237 670
rect 237 608 271 670
rect -271 -670 -237 -608
rect 237 -670 271 -608
rect -271 -704 -175 -670
rect 175 -704 271 -670
<< viali >>
rect -125 159 125 556
rect -125 -556 125 -159
<< metal1 >>
rect -131 556 131 568
rect -131 159 -125 556
rect 125 159 131 556
rect -131 147 131 159
rect -131 -159 131 -147
rect -131 -556 -125 -159
rect 125 -556 131 -159
rect -131 -568 131 -556
<< properties >>
string FIXED_BBOX -254 -687 254 687
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.579 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 2.506k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
