magic
tech sky130A
magscale 1 2
timestamp 1750828667
<< viali >>
rect 503 2548 537 2582
rect 647 2548 681 2582
<< metal1 >>
rect 77 2788 1067 2936
rect 490 2594 550 2600
rect 490 2528 550 2534
rect 634 2594 694 2600
rect 634 2528 694 2534
rect 77 1968 1067 2224
<< via1 >>
rect 490 2582 550 2594
rect 490 2548 503 2582
rect 503 2548 537 2582
rect 537 2548 550 2582
rect 490 2534 550 2548
rect 634 2582 694 2594
rect 634 2548 647 2582
rect 647 2548 681 2582
rect 681 2548 694 2582
rect 634 2534 694 2548
<< metal2 >>
rect 490 2594 550 2600
rect 490 2142 550 2534
rect 634 2594 694 2936
rect 634 2528 694 2534
rect 490 2086 492 2142
rect 548 2086 550 2142
rect 490 2077 550 2086
<< via2 >>
rect 492 2086 548 2142
rect 492 1474 548 1530
<< metal3 >>
rect 487 2142 553 2147
rect 487 2086 492 2142
rect 548 2086 553 2142
rect 487 1530 553 2086
rect 487 1474 492 1530
rect 548 1474 553 1530
rect 487 1469 553 1474
use lvsf  lvsf_0
timestamp 1750828667
transform 1 0 -2560 0 1 1768
box 2571 -1765 3693 326
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1704896540
transform 1 0 428 0 -1 2913
box -66 -43 354 897
<< end >>
