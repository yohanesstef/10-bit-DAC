magic
tech sky130A
magscale 1 2
timestamp 1749844197
<< error_p >>
rect 12636 54467 12663 54477
rect 12610 54407 12663 54467
rect 12636 54397 12663 54407
rect 12664 54467 12691 54477
rect 14141 54467 14168 54477
rect 12664 54407 12717 54467
rect 14115 54407 14168 54467
rect 12664 54397 12691 54407
rect 14141 54397 14168 54407
rect 14169 54467 14196 54477
rect 15646 54467 15673 54477
rect 14169 54407 14222 54467
rect 15620 54407 15673 54467
rect 14169 54397 14196 54407
rect 15646 54397 15673 54407
rect 15674 54467 15701 54477
rect 17151 54467 17178 54477
rect 15674 54407 15727 54467
rect 17125 54407 17178 54467
rect 15674 54397 15701 54407
rect 17151 54397 17178 54407
rect 17179 54467 17206 54477
rect 18656 54467 18683 54477
rect 17179 54407 17232 54467
rect 18630 54407 18683 54467
rect 17179 54397 17206 54407
rect 18656 54397 18683 54407
rect 18684 54467 18711 54477
rect 18684 54407 18737 54467
rect 18684 54397 18711 54407
rect 12636 54309 12663 54369
rect 12664 54309 12691 54369
rect 14141 54309 14168 54369
rect 14169 54309 14196 54369
rect 15646 54309 15673 54369
rect 15674 54309 15701 54369
rect 17151 54309 17178 54369
rect 17179 54309 17206 54369
rect 18656 54309 18683 54369
rect 18684 54309 18711 54369
rect 12636 53381 12663 53441
rect 12664 53381 12691 53441
rect 14141 53381 14168 53441
rect 14169 53381 14196 53441
rect 15646 53381 15673 53441
rect 15674 53381 15701 53441
rect 17151 53381 17178 53441
rect 17179 53381 17206 53441
rect 18656 53381 18683 53441
rect 18684 53381 18711 53441
rect 12636 53343 12663 53353
rect 12610 53283 12663 53343
rect 12636 53273 12663 53283
rect 12664 53343 12691 53353
rect 14141 53343 14168 53353
rect 12664 53283 12717 53343
rect 14115 53283 14168 53343
rect 12664 53273 12691 53283
rect 14141 53273 14168 53283
rect 14169 53343 14196 53353
rect 15646 53343 15673 53353
rect 14169 53283 14222 53343
rect 15620 53283 15673 53343
rect 14169 53273 14196 53283
rect 15646 53273 15673 53283
rect 15674 53343 15701 53353
rect 17151 53343 17178 53353
rect 15674 53283 15727 53343
rect 17125 53283 17178 53343
rect 15674 53273 15701 53283
rect 17151 53273 17178 53283
rect 17179 53343 17206 53353
rect 18656 53343 18683 53353
rect 17179 53283 17232 53343
rect 18630 53283 18683 53343
rect 17179 53273 17206 53283
rect 18656 53273 18683 53283
rect 18684 53343 18711 53353
rect 18684 53283 18737 53343
rect 18684 53273 18711 53283
rect 12636 53185 12663 53245
rect 12664 53185 12691 53245
rect 14141 53185 14168 53245
rect 14169 53185 14196 53245
rect 15646 53185 15673 53245
rect 15674 53185 15701 53245
rect 17151 53185 17178 53245
rect 17179 53185 17206 53245
rect 18656 53185 18683 53245
rect 18684 53185 18711 53245
rect 12636 52257 12663 52317
rect 12664 52257 12691 52317
rect 14141 52257 14168 52317
rect 14169 52257 14196 52317
rect 15646 52257 15673 52317
rect 15674 52257 15701 52317
rect 17151 52257 17178 52317
rect 17179 52257 17206 52317
rect 18656 52257 18683 52317
rect 18684 52257 18711 52317
rect 12636 52219 12663 52229
rect 12610 52159 12663 52219
rect 12636 52149 12663 52159
rect 12664 52219 12691 52229
rect 14141 52219 14168 52229
rect 12664 52159 12717 52219
rect 14115 52159 14168 52219
rect 12664 52149 12691 52159
rect 14141 52149 14168 52159
rect 14169 52219 14196 52229
rect 15646 52219 15673 52229
rect 14169 52159 14222 52219
rect 15620 52159 15673 52219
rect 14169 52149 14196 52159
rect 15646 52149 15673 52159
rect 15674 52219 15701 52229
rect 17151 52219 17178 52229
rect 15674 52159 15727 52219
rect 17125 52159 17178 52219
rect 15674 52149 15701 52159
rect 17151 52149 17178 52159
rect 17179 52219 17206 52229
rect 18656 52219 18683 52229
rect 17179 52159 17232 52219
rect 18630 52159 18683 52219
rect 17179 52149 17206 52159
rect 18656 52149 18683 52159
rect 18684 52219 18711 52229
rect 18684 52159 18737 52219
rect 18684 52149 18711 52159
rect 1002 50345 1029 50355
rect 976 50285 1029 50345
rect 1002 50275 1029 50285
rect 1030 50345 1057 50355
rect 2507 50345 2534 50355
rect 1030 50285 1083 50345
rect 2481 50285 2534 50345
rect 1030 50275 1057 50285
rect 2507 50275 2534 50285
rect 2535 50345 2562 50355
rect 4012 50345 4039 50355
rect 2535 50285 2588 50345
rect 3986 50285 4039 50345
rect 2535 50275 2562 50285
rect 4012 50275 4039 50285
rect 4040 50345 4067 50355
rect 5517 50345 5544 50355
rect 4040 50285 4093 50345
rect 5491 50285 5544 50345
rect 4040 50275 4067 50285
rect 5517 50275 5544 50285
rect 5545 50345 5572 50355
rect 7022 50345 7049 50355
rect 5545 50285 5598 50345
rect 6996 50285 7049 50345
rect 5545 50275 5572 50285
rect 7022 50275 7049 50285
rect 7050 50345 7077 50355
rect 7050 50285 7103 50345
rect 7050 50275 7077 50285
rect 1002 50187 1029 50247
rect 1030 50187 1057 50247
rect 2507 50187 2534 50247
rect 2535 50187 2562 50247
rect 4012 50187 4039 50247
rect 4040 50187 4067 50247
rect 5517 50187 5544 50247
rect 5545 50187 5572 50247
rect 7022 50187 7049 50247
rect 7050 50187 7077 50247
rect 1002 49259 1029 49319
rect 1030 49259 1057 49319
rect 2507 49259 2534 49319
rect 2535 49259 2562 49319
rect 4012 49259 4039 49319
rect 4040 49259 4067 49319
rect 5517 49259 5544 49319
rect 5545 49259 5572 49319
rect 7022 49259 7049 49319
rect 7050 49259 7077 49319
rect 1002 49221 1029 49231
rect 976 49161 1029 49221
rect 1002 49151 1029 49161
rect 1030 49221 1057 49231
rect 2507 49221 2534 49231
rect 1030 49161 1083 49221
rect 2481 49161 2534 49221
rect 1030 49151 1057 49161
rect 2507 49151 2534 49161
rect 2535 49221 2562 49231
rect 4012 49221 4039 49231
rect 2535 49161 2588 49221
rect 3986 49161 4039 49221
rect 2535 49151 2562 49161
rect 4012 49151 4039 49161
rect 4040 49221 4067 49231
rect 5517 49221 5544 49231
rect 4040 49161 4093 49221
rect 5491 49161 5544 49221
rect 4040 49151 4067 49161
rect 5517 49151 5544 49161
rect 5545 49221 5572 49231
rect 7022 49221 7049 49231
rect 5545 49161 5598 49221
rect 6996 49161 7049 49221
rect 5545 49151 5572 49161
rect 7022 49151 7049 49161
rect 7050 49221 7077 49231
rect 7050 49161 7103 49221
rect 7050 49151 7077 49161
rect 1002 49063 1029 49123
rect 1030 49063 1057 49123
rect 2507 49063 2534 49123
rect 2535 49063 2562 49123
rect 4012 49063 4039 49123
rect 4040 49063 4067 49123
rect 5517 49063 5544 49123
rect 5545 49063 5572 49123
rect 7022 49063 7049 49123
rect 7050 49063 7077 49123
rect 1002 48135 1029 48195
rect 1030 48135 1057 48195
rect 2507 48135 2534 48195
rect 2535 48135 2562 48195
rect 4012 48135 4039 48195
rect 4040 48135 4067 48195
rect 5517 48135 5544 48195
rect 5545 48135 5572 48195
rect 7022 48135 7049 48195
rect 7050 48135 7077 48195
rect 1002 48097 1029 48107
rect 976 48064 1029 48097
rect -464 48037 1029 48064
rect -438 48027 1029 48037
rect 1030 48097 1057 48107
rect 2507 48097 2534 48107
rect 1030 48064 1083 48097
rect 2481 48064 2534 48097
rect 1030 48027 2534 48064
rect 2535 48097 2562 48107
rect 4012 48097 4039 48107
rect 2535 48064 2588 48097
rect 3986 48064 4039 48097
rect 2535 48027 4039 48064
rect 4040 48097 4067 48107
rect 5517 48097 5544 48107
rect 4040 48064 4093 48097
rect 5491 48064 5544 48097
rect 4040 48027 5544 48064
rect 5545 48097 5572 48107
rect 7022 48097 7049 48107
rect 5545 48064 5598 48097
rect 6996 48064 7049 48097
rect 5545 48027 7049 48064
rect 7050 48097 7077 48107
rect 7050 48064 7103 48097
rect 7050 48027 8554 48064
rect -410 47983 1094 48020
rect 1041 47950 1094 47983
rect 1067 47940 1094 47950
rect 1095 47983 2599 48020
rect 1095 47950 1148 47983
rect 2546 47950 2599 47983
rect 1095 47940 1122 47950
rect 2572 47940 2599 47950
rect 2600 47983 4104 48020
rect 2600 47950 2653 47983
rect 4051 47950 4104 47983
rect 2600 47940 2627 47950
rect 4077 47940 4104 47950
rect 4105 47983 5609 48020
rect 4105 47950 4158 47983
rect 5556 47950 5609 47983
rect 4105 47940 4132 47950
rect 5582 47940 5609 47950
rect 5610 47983 7114 48020
rect 5610 47950 5663 47983
rect 7061 47950 7114 47983
rect 5610 47940 5637 47950
rect 7087 47940 7114 47950
rect 7115 48010 8582 48020
rect 7115 47983 8608 48010
rect 7115 47950 7168 47983
rect 7115 47940 7142 47950
rect 1067 47852 1094 47912
rect 1095 47852 1122 47912
rect 2572 47852 2599 47912
rect 2600 47852 2627 47912
rect 4077 47852 4104 47912
rect 4105 47852 4132 47912
rect 5582 47852 5609 47912
rect 5610 47852 5637 47912
rect 7087 47852 7114 47912
rect 7115 47852 7142 47912
rect 1067 46924 1094 46984
rect 1095 46924 1122 46984
rect 2572 46924 2599 46984
rect 2600 46924 2627 46984
rect 4077 46924 4104 46984
rect 4105 46924 4132 46984
rect 5582 46924 5609 46984
rect 5610 46924 5637 46984
rect 7087 46924 7114 46984
rect 7115 46924 7142 46984
rect 1067 46886 1094 46896
rect 1041 46826 1094 46886
rect 1067 46816 1094 46826
rect 1095 46886 1122 46896
rect 2572 46886 2599 46896
rect 1095 46826 1148 46886
rect 2546 46826 2599 46886
rect 1095 46816 1122 46826
rect 2572 46816 2599 46826
rect 2600 46886 2627 46896
rect 4077 46886 4104 46896
rect 2600 46826 2653 46886
rect 4051 46826 4104 46886
rect 2600 46816 2627 46826
rect 4077 46816 4104 46826
rect 4105 46886 4132 46896
rect 5582 46886 5609 46896
rect 4105 46826 4158 46886
rect 5556 46826 5609 46886
rect 4105 46816 4132 46826
rect 5582 46816 5609 46826
rect 5610 46886 5637 46896
rect 7087 46886 7114 46896
rect 5610 46826 5663 46886
rect 7061 46826 7114 46886
rect 5610 46816 5637 46826
rect 7087 46816 7114 46826
rect 7115 46886 7142 46896
rect 7115 46826 7168 46886
rect 7115 46816 7142 46826
rect 1067 46728 1094 46788
rect 1095 46728 1122 46788
rect 2572 46728 2599 46788
rect 2600 46728 2627 46788
rect 4077 46728 4104 46788
rect 4105 46728 4132 46788
rect 5582 46728 5609 46788
rect 5610 46728 5637 46788
rect 7087 46728 7114 46788
rect 7115 46728 7142 46788
rect 1067 45834 1094 45860
rect 1095 45834 1122 45860
rect 2572 45834 2599 45860
rect 2600 45834 2627 45860
rect 4077 45834 4104 45860
rect 4105 45834 4132 45860
rect 5582 45834 5609 45860
rect 5610 45834 5637 45860
rect 7087 45834 7114 45860
rect 7115 45834 7142 45860
rect 1067 45824 1124 45834
rect 2572 45824 2629 45834
rect 4077 45824 4134 45834
rect 5582 45824 5639 45834
rect 7087 45824 7144 45834
rect -333 45816 -100 45824
rect 43 45816 276 45824
rect 419 45816 652 45824
rect 795 45816 1028 45824
rect 1043 45816 1150 45824
rect 1172 45816 1405 45824
rect 1548 45816 1781 45824
rect 1924 45816 2157 45824
rect 2300 45816 2533 45824
rect 2548 45816 2655 45824
rect 2677 45816 2910 45824
rect 3053 45816 3286 45824
rect 3429 45816 3662 45824
rect 3805 45816 4038 45824
rect 4053 45816 4160 45824
rect 4182 45816 4415 45824
rect 4558 45816 4791 45824
rect 4934 45816 5167 45824
rect 5310 45816 5543 45824
rect 5558 45816 5665 45824
rect 5687 45816 5920 45824
rect 6063 45816 6296 45824
rect 6439 45816 6672 45824
rect 6815 45816 7048 45824
rect 7063 45816 7170 45824
rect 7192 45816 7425 45824
rect 7568 45816 7801 45824
rect 7944 45816 8177 45824
rect 8320 45816 8553 45824
rect -408 45800 8621 45816
rect -408 45782 1096 45800
rect 1097 45782 2601 45800
rect 2602 45782 4106 45800
rect 4107 45782 5611 45800
rect 5612 45782 7116 45800
rect 7117 45782 8621 45800
rect -408 45772 8621 45782
rect -408 45764 1096 45772
rect 1097 45764 2601 45772
rect 2602 45764 4106 45772
rect 4107 45764 5611 45772
rect 5612 45764 7116 45772
rect 7117 45764 8621 45772
rect -410 45726 1094 45762
rect 1095 45726 2599 45762
rect 2600 45726 4104 45762
rect 4105 45726 5609 45762
rect 5610 45726 7114 45762
rect 7115 45726 8619 45762
rect -410 45710 8619 45726
rect -331 45702 -98 45710
rect 45 45702 278 45710
rect 421 45702 654 45710
rect 797 45702 1030 45710
rect 1041 45702 1148 45710
rect 1174 45702 1407 45710
rect 1550 45702 1783 45710
rect 1926 45702 2159 45710
rect 2302 45702 2535 45710
rect 2546 45702 2653 45710
rect 2679 45702 2912 45710
rect 3055 45702 3288 45710
rect 3431 45702 3664 45710
rect 3807 45702 4040 45710
rect 4051 45702 4158 45710
rect 4184 45702 4417 45710
rect 4560 45702 4793 45710
rect 4936 45702 5169 45710
rect 5312 45702 5545 45710
rect 5556 45702 5663 45710
rect 5689 45702 5922 45710
rect 6065 45702 6298 45710
rect 6441 45702 6674 45710
rect 6817 45702 7050 45710
rect 7061 45702 7168 45710
rect 7194 45702 7427 45710
rect 7570 45702 7803 45710
rect 7946 45702 8179 45710
rect 8322 45702 8555 45710
rect 1067 45692 1124 45702
rect 2572 45692 2629 45702
rect 4077 45692 4134 45702
rect 5582 45692 5639 45702
rect 7087 45692 7144 45702
rect 1069 45666 1096 45692
rect 1097 45666 1124 45692
rect 2574 45666 2601 45692
rect 2602 45666 2629 45692
rect 4079 45666 4106 45692
rect 4107 45666 4134 45692
rect 5584 45666 5611 45692
rect 5612 45666 5639 45692
rect 7089 45666 7116 45692
rect 7117 45666 7144 45692
rect 1069 44738 1096 44798
rect 1097 44738 1124 44798
rect 2574 44738 2601 44798
rect 2602 44738 2629 44798
rect 4079 44738 4106 44798
rect 4107 44738 4134 44798
rect 5584 44738 5611 44798
rect 5612 44738 5639 44798
rect 7089 44738 7116 44798
rect 7117 44738 7144 44798
rect 1069 44700 1096 44710
rect 1043 44640 1096 44700
rect 1069 44630 1096 44640
rect 1097 44700 1124 44710
rect 2574 44700 2601 44710
rect 1097 44640 1150 44700
rect 2548 44640 2601 44700
rect 1097 44630 1124 44640
rect 2574 44630 2601 44640
rect 2602 44700 2629 44710
rect 4079 44700 4106 44710
rect 2602 44640 2655 44700
rect 4053 44640 4106 44700
rect 2602 44630 2629 44640
rect 4079 44630 4106 44640
rect 4107 44700 4134 44710
rect 5584 44700 5611 44710
rect 4107 44640 4160 44700
rect 5558 44640 5611 44700
rect 4107 44630 4134 44640
rect 5584 44630 5611 44640
rect 5612 44700 5639 44710
rect 7089 44700 7116 44710
rect 5612 44640 5665 44700
rect 7063 44640 7116 44700
rect 5612 44630 5639 44640
rect 7089 44630 7116 44640
rect 7117 44700 7144 44710
rect 7117 44640 7170 44700
rect 7117 44630 7144 44640
rect 1069 44542 1096 44602
rect 1097 44542 1124 44602
rect 2574 44542 2601 44602
rect 2602 44542 2629 44602
rect 4079 44542 4106 44602
rect 4107 44542 4134 44602
rect 5584 44542 5611 44602
rect 5612 44542 5639 44602
rect 7089 44542 7116 44602
rect 7117 44542 7144 44602
rect 1069 43614 1096 43674
rect 1097 43614 1124 43674
rect 2574 43614 2601 43674
rect 2602 43614 2629 43674
rect 4079 43614 4106 43674
rect 4107 43614 4134 43674
rect 5584 43614 5611 43674
rect 5612 43614 5639 43674
rect 7089 43614 7116 43674
rect 7117 43614 7144 43674
rect 1069 43576 1096 43586
rect 1043 43516 1096 43576
rect 1069 43506 1096 43516
rect 1097 43576 1124 43586
rect 2574 43576 2601 43586
rect 1097 43516 1150 43576
rect 2548 43516 2601 43576
rect 1097 43506 1124 43516
rect 2574 43506 2601 43516
rect 2602 43576 2629 43586
rect 4079 43576 4106 43586
rect 2602 43516 2655 43576
rect 4053 43516 4106 43576
rect 2602 43506 2629 43516
rect 4079 43506 4106 43516
rect 4107 43576 4134 43586
rect 5584 43576 5611 43586
rect 4107 43516 4160 43576
rect 5558 43516 5611 43576
rect 4107 43506 4134 43516
rect 5584 43506 5611 43516
rect 5612 43576 5639 43586
rect 7089 43576 7116 43586
rect 5612 43516 5665 43576
rect 7063 43516 7116 43576
rect 5612 43506 5639 43516
rect 7089 43506 7116 43516
rect 7117 43576 7144 43586
rect 7117 43516 7170 43576
rect 7117 43506 7144 43516
rect 34378 18299 34405 18309
rect 34352 18239 34405 18299
rect 34378 18229 34405 18239
rect 34406 18299 34433 18309
rect 35883 18299 35910 18309
rect 34406 18239 34459 18299
rect 35857 18239 35910 18299
rect 34406 18229 34433 18239
rect 35883 18229 35910 18239
rect 35911 18299 35938 18309
rect 37388 18299 37415 18309
rect 35911 18239 35964 18299
rect 37362 18239 37415 18299
rect 35911 18229 35938 18239
rect 37388 18229 37415 18239
rect 37416 18299 37443 18309
rect 38893 18299 38920 18309
rect 37416 18239 37469 18299
rect 38867 18239 38920 18299
rect 37416 18229 37443 18239
rect 38893 18229 38920 18239
rect 38921 18299 38948 18309
rect 40398 18299 40425 18309
rect 38921 18239 38974 18299
rect 40372 18239 40425 18299
rect 38921 18229 38948 18239
rect 40398 18229 40425 18239
rect 40426 18299 40453 18309
rect 40426 18239 40479 18299
rect 40426 18229 40453 18239
rect 34378 18141 34405 18201
rect 34406 18141 34433 18201
rect 35883 18141 35910 18201
rect 35911 18141 35938 18201
rect 37388 18141 37415 18201
rect 37416 18141 37443 18201
rect 38893 18141 38920 18201
rect 38921 18141 38948 18201
rect 40398 18141 40425 18201
rect 40426 18141 40453 18201
rect 34378 17213 34405 17273
rect 34406 17213 34433 17273
rect 35883 17213 35910 17273
rect 35911 17213 35938 17273
rect 37388 17213 37415 17273
rect 37416 17213 37443 17273
rect 38893 17213 38920 17273
rect 38921 17213 38948 17273
rect 40398 17213 40425 17273
rect 40426 17213 40453 17273
rect 34378 17175 34405 17185
rect 34352 17115 34405 17175
rect 34378 17105 34405 17115
rect 34406 17175 34433 17185
rect 35883 17175 35910 17185
rect 34406 17115 34459 17175
rect 35857 17115 35910 17175
rect 34406 17105 34433 17115
rect 35883 17105 35910 17115
rect 35911 17175 35938 17185
rect 37388 17175 37415 17185
rect 35911 17115 35964 17175
rect 37362 17115 37415 17175
rect 35911 17105 35938 17115
rect 37388 17105 37415 17115
rect 37416 17175 37443 17185
rect 38893 17175 38920 17185
rect 37416 17115 37469 17175
rect 38867 17115 38920 17175
rect 37416 17105 37443 17115
rect 38893 17105 38920 17115
rect 38921 17175 38948 17185
rect 40398 17175 40425 17185
rect 38921 17115 38974 17175
rect 40372 17115 40425 17175
rect 38921 17105 38948 17115
rect 40398 17105 40425 17115
rect 40426 17175 40453 17185
rect 40426 17115 40479 17175
rect 40426 17105 40453 17115
rect 34378 17017 34405 17077
rect 34406 17017 34433 17077
rect 35883 17017 35910 17077
rect 35911 17017 35938 17077
rect 37388 17017 37415 17077
rect 37416 17017 37443 17077
rect 38893 17017 38920 17077
rect 38921 17017 38948 17077
rect 40398 17017 40425 17077
rect 40426 17017 40453 17077
rect 34378 16089 34405 16149
rect 34406 16089 34433 16149
rect 35883 16089 35910 16149
rect 35911 16089 35938 16149
rect 37388 16089 37415 16149
rect 37416 16089 37443 16149
rect 38893 16089 38920 16149
rect 38921 16089 38948 16149
rect 40398 16089 40425 16149
rect 40426 16089 40453 16149
rect 34378 16051 34405 16061
rect 34352 15991 34405 16051
rect 34378 15981 34405 15991
rect 34406 16051 34433 16061
rect 35883 16051 35910 16061
rect 34406 15991 34459 16051
rect 35857 15991 35910 16051
rect 34406 15981 34433 15991
rect 35883 15981 35910 15991
rect 35911 16051 35938 16061
rect 37388 16051 37415 16061
rect 35911 15991 35964 16051
rect 37362 15991 37415 16051
rect 35911 15981 35938 15991
rect 37388 15981 37415 15991
rect 37416 16051 37443 16061
rect 38893 16051 38920 16061
rect 37416 15991 37469 16051
rect 38867 15991 38920 16051
rect 37416 15981 37443 15991
rect 38893 15981 38920 15991
rect 38921 16051 38948 16061
rect 40398 16051 40425 16061
rect 38921 15991 38974 16051
rect 40372 15991 40425 16051
rect 38921 15981 38948 15991
rect 40398 15981 40425 15991
rect 40426 16051 40453 16061
rect 40426 15991 40479 16051
rect 40426 15981 40453 15991
rect 22744 14177 22771 14187
rect 22718 14117 22771 14177
rect 22744 14107 22771 14117
rect 22772 14177 22799 14187
rect 24249 14177 24276 14187
rect 22772 14117 22825 14177
rect 24223 14117 24276 14177
rect 22772 14107 22799 14117
rect 24249 14107 24276 14117
rect 24277 14177 24304 14187
rect 25754 14177 25781 14187
rect 24277 14117 24330 14177
rect 25728 14117 25781 14177
rect 24277 14107 24304 14117
rect 25754 14107 25781 14117
rect 25782 14177 25809 14187
rect 27259 14177 27286 14187
rect 25782 14117 25835 14177
rect 27233 14117 27286 14177
rect 25782 14107 25809 14117
rect 27259 14107 27286 14117
rect 27287 14177 27314 14187
rect 28764 14177 28791 14187
rect 27287 14117 27340 14177
rect 28738 14117 28791 14177
rect 27287 14107 27314 14117
rect 28764 14107 28791 14117
rect 28792 14177 28819 14187
rect 28792 14117 28845 14177
rect 28792 14107 28819 14117
rect 22744 14019 22771 14079
rect 22772 14019 22799 14079
rect 24249 14019 24276 14079
rect 24277 14019 24304 14079
rect 25754 14019 25781 14079
rect 25782 14019 25809 14079
rect 27259 14019 27286 14079
rect 27287 14019 27314 14079
rect 28764 14019 28791 14079
rect 28792 14019 28819 14079
rect 22744 13091 22771 13151
rect 22772 13091 22799 13151
rect 24249 13091 24276 13151
rect 24277 13091 24304 13151
rect 25754 13091 25781 13151
rect 25782 13091 25809 13151
rect 27259 13091 27286 13151
rect 27287 13091 27314 13151
rect 28764 13091 28791 13151
rect 28792 13091 28819 13151
rect 22744 13053 22771 13063
rect 22718 12993 22771 13053
rect 22744 12983 22771 12993
rect 22772 13053 22799 13063
rect 24249 13053 24276 13063
rect 22772 12993 22825 13053
rect 24223 12993 24276 13053
rect 22772 12983 22799 12993
rect 24249 12983 24276 12993
rect 24277 13053 24304 13063
rect 25754 13053 25781 13063
rect 24277 12993 24330 13053
rect 25728 12993 25781 13053
rect 24277 12983 24304 12993
rect 25754 12983 25781 12993
rect 25782 13053 25809 13063
rect 27259 13053 27286 13063
rect 25782 12993 25835 13053
rect 27233 12993 27286 13053
rect 25782 12983 25809 12993
rect 27259 12983 27286 12993
rect 27287 13053 27314 13063
rect 28764 13053 28791 13063
rect 27287 12993 27340 13053
rect 28738 12993 28791 13053
rect 27287 12983 27314 12993
rect 28764 12983 28791 12993
rect 28792 13053 28819 13063
rect 28792 12993 28845 13053
rect 28792 12983 28819 12993
rect 22744 12895 22771 12955
rect 22772 12895 22799 12955
rect 24249 12895 24276 12955
rect 24277 12895 24304 12955
rect 25754 12895 25781 12955
rect 25782 12895 25809 12955
rect 27259 12895 27286 12955
rect 27287 12895 27314 12955
rect 28764 12895 28791 12955
rect 28792 12895 28819 12955
rect 22744 11967 22771 12027
rect 22772 11967 22799 12027
rect 24249 11967 24276 12027
rect 24277 11967 24304 12027
rect 25754 11967 25781 12027
rect 25782 11967 25809 12027
rect 27259 11967 27286 12027
rect 27287 11967 27314 12027
rect 28764 11967 28791 12027
rect 28792 11967 28819 12027
rect 22744 11929 22771 11939
rect 22718 11896 22771 11929
rect 21527 11859 22771 11896
rect 22772 11929 22799 11939
rect 24249 11929 24276 11939
rect 22772 11896 22825 11929
rect 24223 11896 24276 11929
rect 22772 11859 24276 11896
rect 24277 11929 24304 11939
rect 25754 11929 25781 11939
rect 24277 11896 24330 11929
rect 25728 11896 25781 11929
rect 24277 11859 25781 11896
rect 25782 11929 25809 11939
rect 27259 11929 27286 11939
rect 25782 11896 25835 11929
rect 27233 11896 27286 11929
rect 25782 11859 27286 11896
rect 27287 11929 27314 11939
rect 28764 11929 28791 11939
rect 27287 11896 27340 11929
rect 28738 11896 28791 11929
rect 27287 11859 28791 11896
rect 28792 11929 28819 11939
rect 28792 11896 28845 11929
rect 28792 11859 30296 11896
rect 21527 11815 22836 11852
rect 22783 11782 22836 11815
rect 22809 11772 22836 11782
rect 22837 11815 24341 11852
rect 22837 11782 22890 11815
rect 24288 11782 24341 11815
rect 22837 11772 22864 11782
rect 24314 11772 24341 11782
rect 24342 11815 25846 11852
rect 24342 11782 24395 11815
rect 25793 11782 25846 11815
rect 24342 11772 24369 11782
rect 25819 11772 25846 11782
rect 25847 11815 27351 11852
rect 25847 11782 25900 11815
rect 27298 11782 27351 11815
rect 25847 11772 25874 11782
rect 27324 11772 27351 11782
rect 27352 11815 28856 11852
rect 27352 11782 27405 11815
rect 28803 11782 28856 11815
rect 27352 11772 27379 11782
rect 28829 11772 28856 11782
rect 28857 11842 30324 11852
rect 28857 11815 30350 11842
rect 28857 11782 28910 11815
rect 28857 11772 28884 11782
rect 22809 11684 22836 11744
rect 22837 11684 22864 11744
rect 24314 11684 24341 11744
rect 24342 11684 24369 11744
rect 25819 11684 25846 11744
rect 25847 11684 25874 11744
rect 27324 11684 27351 11744
rect 27352 11684 27379 11744
rect 28829 11684 28856 11744
rect 28857 11684 28884 11744
rect 22809 10756 22836 10816
rect 22837 10756 22864 10816
rect 24314 10756 24341 10816
rect 24342 10756 24369 10816
rect 25819 10756 25846 10816
rect 25847 10756 25874 10816
rect 27324 10756 27351 10816
rect 27352 10756 27379 10816
rect 28829 10756 28856 10816
rect 28857 10756 28884 10816
rect 22809 10718 22836 10728
rect 22783 10658 22836 10718
rect 22809 10648 22836 10658
rect 22837 10718 22864 10728
rect 24314 10718 24341 10728
rect 22837 10658 22890 10718
rect 24288 10658 24341 10718
rect 22837 10648 22864 10658
rect 24314 10648 24341 10658
rect 24342 10718 24369 10728
rect 25819 10718 25846 10728
rect 24342 10658 24395 10718
rect 25793 10658 25846 10718
rect 24342 10648 24369 10658
rect 25819 10648 25846 10658
rect 25847 10718 25874 10728
rect 27324 10718 27351 10728
rect 25847 10658 25900 10718
rect 27298 10658 27351 10718
rect 25847 10648 25874 10658
rect 27324 10648 27351 10658
rect 27352 10718 27379 10728
rect 28829 10718 28856 10728
rect 27352 10658 27405 10718
rect 28803 10658 28856 10718
rect 27352 10648 27379 10658
rect 28829 10648 28856 10658
rect 28857 10718 28884 10728
rect 28857 10658 28910 10718
rect 28857 10648 28884 10658
rect 22809 10560 22836 10620
rect 22837 10560 22864 10620
rect 24314 10560 24341 10620
rect 24342 10560 24369 10620
rect 25819 10560 25846 10620
rect 25847 10560 25874 10620
rect 27324 10560 27351 10620
rect 27352 10560 27379 10620
rect 28829 10560 28856 10620
rect 28857 10560 28884 10620
rect 22809 9666 22836 9692
rect 22837 9666 22864 9692
rect 24314 9666 24341 9692
rect 24342 9666 24369 9692
rect 25819 9666 25846 9692
rect 25847 9666 25874 9692
rect 27324 9666 27351 9692
rect 27352 9666 27379 9692
rect 28829 9666 28856 9692
rect 28857 9666 28884 9692
rect 22809 9656 22866 9666
rect 24314 9656 24371 9666
rect 25819 9656 25876 9666
rect 27324 9656 27381 9666
rect 28829 9656 28886 9666
rect 21620 9648 21642 9656
rect 21785 9648 21796 9656
rect 21620 9622 21796 9648
rect 21996 9648 22018 9656
rect 22161 9648 22172 9656
rect 21996 9622 22172 9648
rect 22372 9648 22394 9656
rect 22537 9648 22548 9656
rect 22372 9622 22548 9648
rect 22748 9648 22770 9656
rect 22785 9648 22892 9656
rect 22914 9648 23147 9656
rect 23290 9648 23523 9656
rect 23666 9648 23899 9656
rect 24042 9648 24275 9656
rect 24290 9648 24397 9656
rect 24419 9648 24652 9656
rect 24795 9648 25028 9656
rect 25171 9648 25404 9656
rect 25547 9648 25780 9656
rect 25795 9648 25902 9656
rect 25924 9648 26157 9656
rect 26300 9648 26533 9656
rect 26676 9648 26909 9656
rect 27052 9648 27285 9656
rect 27300 9648 27407 9656
rect 27429 9648 27662 9656
rect 27805 9648 28038 9656
rect 28181 9648 28414 9656
rect 28557 9648 28790 9656
rect 28805 9648 28912 9656
rect 28934 9648 29167 9656
rect 29310 9648 29543 9656
rect 29686 9648 29919 9656
rect 30062 9648 30295 9656
rect 22748 9632 30363 9648
rect 22748 9622 22838 9632
rect 21527 9614 22838 9622
rect 22839 9614 24343 9632
rect 24344 9614 25848 9632
rect 25849 9614 27353 9632
rect 27354 9614 28858 9632
rect 28859 9614 30363 9632
rect 21527 9604 30363 9614
rect 21527 9596 22838 9604
rect 22839 9596 24343 9604
rect 24344 9596 25848 9604
rect 25849 9596 27353 9604
rect 27354 9596 28858 9604
rect 28859 9596 30363 9604
rect 21527 9568 22836 9594
rect 21622 9542 21798 9568
rect 21622 9534 21644 9542
rect 21787 9534 21798 9542
rect 21998 9542 22174 9568
rect 21998 9534 22020 9542
rect 22163 9534 22174 9542
rect 22374 9542 22550 9568
rect 22374 9534 22396 9542
rect 22539 9534 22550 9542
rect 22750 9558 22836 9568
rect 22837 9558 24341 9594
rect 24342 9558 25846 9594
rect 25847 9558 27351 9594
rect 27352 9558 28856 9594
rect 28857 9558 30361 9594
rect 22750 9542 30361 9558
rect 22750 9534 22772 9542
rect 22783 9534 22890 9542
rect 22916 9534 23149 9542
rect 23292 9534 23525 9542
rect 23668 9534 23901 9542
rect 24044 9534 24277 9542
rect 24288 9534 24395 9542
rect 24421 9534 24654 9542
rect 24797 9534 25030 9542
rect 25173 9534 25406 9542
rect 25549 9534 25782 9542
rect 25793 9534 25900 9542
rect 25926 9534 26159 9542
rect 26302 9534 26535 9542
rect 26678 9534 26911 9542
rect 27054 9534 27287 9542
rect 27298 9534 27405 9542
rect 27431 9534 27664 9542
rect 27807 9534 28040 9542
rect 28183 9534 28416 9542
rect 28559 9534 28792 9542
rect 28803 9534 28910 9542
rect 28936 9534 29169 9542
rect 29312 9534 29545 9542
rect 29688 9534 29921 9542
rect 30064 9534 30297 9542
rect 22809 9524 22866 9534
rect 24314 9524 24371 9534
rect 25819 9524 25876 9534
rect 27324 9524 27381 9534
rect 28829 9524 28886 9534
rect 22811 9498 22838 9524
rect 22839 9498 22866 9524
rect 24316 9498 24343 9524
rect 24344 9498 24371 9524
rect 25821 9498 25848 9524
rect 25849 9498 25876 9524
rect 27326 9498 27353 9524
rect 27354 9498 27381 9524
rect 28831 9498 28858 9524
rect 28859 9498 28886 9524
rect 22811 8570 22838 8630
rect 22839 8570 22866 8630
rect 24316 8570 24343 8630
rect 24344 8570 24371 8630
rect 25821 8570 25848 8630
rect 25849 8570 25876 8630
rect 27326 8570 27353 8630
rect 27354 8570 27381 8630
rect 28831 8570 28858 8630
rect 28859 8570 28886 8630
rect 22811 8532 22838 8542
rect 22785 8472 22838 8532
rect 22811 8462 22838 8472
rect 22839 8532 22866 8542
rect 24316 8532 24343 8542
rect 22839 8472 22892 8532
rect 24290 8472 24343 8532
rect 22839 8462 22866 8472
rect 24316 8462 24343 8472
rect 24344 8532 24371 8542
rect 25821 8532 25848 8542
rect 24344 8472 24397 8532
rect 25795 8472 25848 8532
rect 24344 8462 24371 8472
rect 25821 8462 25848 8472
rect 25849 8532 25876 8542
rect 27326 8532 27353 8542
rect 25849 8472 25902 8532
rect 27300 8472 27353 8532
rect 25849 8462 25876 8472
rect 27326 8462 27353 8472
rect 27354 8532 27381 8542
rect 28831 8532 28858 8542
rect 27354 8472 27407 8532
rect 28805 8472 28858 8532
rect 27354 8462 27381 8472
rect 28831 8462 28858 8472
rect 28859 8532 28886 8542
rect 28859 8472 28912 8532
rect 28859 8462 28886 8472
rect 22811 8374 22838 8434
rect 22839 8374 22866 8434
rect 24316 8374 24343 8434
rect 24344 8374 24371 8434
rect 25821 8374 25848 8434
rect 25849 8374 25876 8434
rect 27326 8374 27353 8434
rect 27354 8374 27381 8434
rect 28831 8374 28858 8434
rect 28859 8374 28886 8434
rect 22811 7446 22838 7506
rect 22839 7446 22866 7506
rect 24316 7446 24343 7506
rect 24344 7446 24371 7506
rect 25821 7446 25848 7506
rect 25849 7446 25876 7506
rect 27326 7446 27353 7506
rect 27354 7446 27381 7506
rect 28831 7446 28858 7506
rect 28859 7446 28886 7506
rect 22811 7408 22838 7418
rect 22785 7348 22838 7408
rect 22811 7338 22838 7348
rect 22839 7408 22866 7418
rect 24316 7408 24343 7418
rect 22839 7348 22892 7408
rect 24290 7348 24343 7408
rect 22839 7338 22866 7348
rect 24316 7338 24343 7348
rect 24344 7408 24371 7418
rect 25821 7408 25848 7418
rect 24344 7348 24397 7408
rect 25795 7348 25848 7408
rect 24344 7338 24371 7348
rect 25821 7338 25848 7348
rect 25849 7408 25876 7418
rect 27326 7408 27353 7418
rect 25849 7348 25902 7408
rect 27300 7348 27353 7408
rect 25849 7338 25876 7348
rect 27326 7338 27353 7348
rect 27354 7408 27381 7418
rect 28831 7408 28858 7418
rect 27354 7348 27407 7408
rect 28805 7348 28858 7408
rect 27354 7338 27381 7348
rect 28831 7338 28858 7348
rect 28859 7408 28886 7418
rect 28859 7348 28912 7408
rect 28859 7338 28886 7348
rect 14782 1869 14878 2399
<< error_s >>
rect 21278 11869 21527 11896
rect 21304 11859 21527 11869
rect 21332 11815 21527 11852
rect 21409 9648 21527 9656
rect 21334 9596 21527 9648
rect 21332 9542 21527 9594
rect 21411 9534 21527 9542
<< error_ps >>
rect 21527 9622 21620 9656
rect 21796 9622 21996 9656
rect 22172 9622 22372 9656
rect 22548 9622 22748 9656
rect 21527 9534 21622 9568
rect 21798 9534 21998 9568
rect 22174 9534 22374 9568
rect 22550 9534 22750 9568
use cm_pcell_1_view  cm_pcell_1_view_0
timestamp 1749844197
transform 1 0 -1555 0 1 49033
box 1014 -5583 21819 5500
use cm_pcell_1_view  cm_pcell_1_view_1
timestamp 1749844197
transform 1 0 20187 0 1 12865
box 1014 -5583 21819 5500
use top_digital_cell  top_digital_cell_0
timestamp 1749834095
transform 1 0 -201 0 1 62
box -31 -831 19387 4119
use top_segment_1  top_segment_1_0
timestamp 1749633251
transform 0 1 -128 -1 0 21427
box -385 -49 14453 8429
use top_segment_2  top_segment_2_0
timestamp 1749580325
transform 0 -1 20281 1 0 11235
box -870 14 15704 7051
use top_segment_3  top_segment_3_0
timestamp 1749552768
transform 0 -1 20508 1 0 22318
box 5007 266 11251 6636
use top_segment_4  top_segment_4_1
timestamp 1749664768
transform 0 1 12179 -1 0 65606
box 29493 -12226 43322 -3773
<< end >>
