.subckt rseg_3_v3 v0 v1 v2 v3 v4 v5 v6 v7 v8 v9 v10 v11 v12 v13 v14 v15 v16 gnd
XR1 v0 v1 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.0665 mult=1 m=1
XR2 v1 v2 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.1033 mult=1 m=1
XR3 v2 v3 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.1217 mult=1 m=1
XR4 v3 v4 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.1400 mult=1 m=1
XR5 v4 v5 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.1951 mult=1 m=1
XR6 v5 v6 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.2134 mult=1 m=1
XR7 v6 v7 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.2501 mult=1 m=1
XR8 v7 v8 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.3052 mult=1 m=1
XR9 v8 v9 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.3419 mult=1 m=1
XR10 v9 v10 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.3970 mult=1 m=1
XR11 v10 v11 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.4338 mult=1 m=1
XR12 v11 v12 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.5255 mult=1 m=1
XR13 v12 v13 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.5806 mult=1 m=1
XR14 v13 v14 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6724 mult=1 m=1
XR15 v14 v15 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.7642 mult=1 m=1
XR16 v15 v16 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.8743 mult=1 m=1
.ends