magic
tech sky130A
magscale 1 2
timestamp 1749563245
<< pwell >>
rect 22810 -13247 39241 -9665
<< psubdiff >>
rect 22846 -9761 23106 -9701
rect 38945 -9761 39205 -9701
rect 22846 -9961 22906 -9761
rect 22846 -13151 22906 -12951
rect 39145 -9961 39205 -9761
rect 39145 -13151 39205 -12951
rect 22846 -13211 23105 -13151
rect 38944 -13211 39205 -13151
<< psubdiffcont >>
rect 23106 -9761 38945 -9701
rect 22846 -12951 22906 -9961
rect 39145 -12951 39205 -9961
rect 23105 -13211 38944 -13151
<< locali >>
rect 22846 -9761 23106 -9701
rect 38945 -9761 39205 -9701
rect 22846 -9961 22906 -9761
rect 23260 -9857 23692 -9761
rect 25974 -9857 26406 -9761
rect 27053 -9857 27485 -9761
rect 28487 -9857 28919 -9761
rect 29463 -9857 29895 -9761
rect 30887 -9857 31319 -9761
rect 31951 -9857 32383 -9761
rect 33293 -9857 33725 -9761
rect 34272 -9857 34704 -9761
rect 35624 -9857 36056 -9761
rect 36689 -9857 37121 -9761
rect 38359 -9857 38791 -9761
rect 22846 -13151 22906 -12951
rect 39145 -9961 39205 -9761
rect 23752 -13151 24184 -13055
rect 25482 -13151 25914 -13055
rect 26935 -13151 27367 -13055
rect 28605 -13151 29037 -13055
rect 29504 -13151 29936 -13055
rect 30846 -13151 31278 -13055
rect 31951 -13151 32383 -13055
rect 33293 -13151 33725 -13055
rect 34231 -13151 34663 -13055
rect 35665 -13151 36097 -13055
rect 36813 -13151 37245 -13055
rect 38257 -13151 38689 -13055
rect 39145 -13151 39205 -12951
rect 22846 -13211 23105 -13151
rect 38944 -13211 39205 -13151
<< metal1 >>
rect 36342 -10191 36343 -10042
<< via1 >>
rect 26334 -10453 26394 -10191
rect 28847 -10453 28907 -10191
rect 31247 -10453 31307 -10191
rect 33653 -10453 33713 -10191
rect 35984 -10453 36044 -10191
rect 38719 -10453 38779 -10191
rect 26686 -12721 26746 -12459
rect 28965 -12721 29025 -12459
rect 31599 -12721 31659 -12459
rect 33653 -12721 33713 -12459
rect 36336 -12721 36396 -12459
rect 38612 -12721 38672 -12459
<< metal2 >>
rect 22810 -10453 26334 -10191
rect 26394 -10453 26400 -10191
rect 28841 -10453 28847 -10191
rect 28907 -10453 31247 -10191
rect 31307 -10453 31313 -10191
rect 33647 -10453 33653 -10191
rect 33713 -10453 35984 -10191
rect 36044 -10453 36050 -10191
rect 38713 -10453 38719 -10191
rect 38779 -10453 39241 -10191
rect 26680 -12721 26686 -12459
rect 26746 -12721 28965 -12459
rect 29025 -12721 29031 -12459
rect 31593 -12721 31599 -12459
rect 31659 -12721 33653 -12459
rect 33713 -12721 33719 -12459
rect 36330 -12721 36336 -12459
rect 36396 -12721 38612 -12459
rect 38672 -12721 38678 -12459
use rseg_1_pin_4  rseg_1_pin_4_0
timestamp 1749560624
transform 1 0 21462 0 1 12573
box 1540 -22764 1864 -22616
use rseg_1_pin_4  rseg_1_pin_4_1
timestamp 1749560624
transform 1 0 24800 0 1 12573
box 1540 -22764 1864 -22616
use rseg_1_pin_4  rseg_1_pin_4_2
timestamp 1749560624
transform 1 0 27313 0 1 12573
box 1540 -22764 1864 -22616
use rseg_1_pin_4  rseg_1_pin_4_3
timestamp 1749560624
transform 1 0 27665 0 1 12573
box 1540 -22764 1864 -22616
use rseg_1_pin_4  rseg_1_pin_4_4
timestamp 1749560624
transform 1 0 29713 0 1 12573
box 1540 -22764 1864 -22616
use rseg_1_pin_4  rseg_1_pin_4_5
timestamp 1749560624
transform 1 0 32119 0 1 12573
box 1540 -22764 1864 -22616
use rseg_1_pin_4  rseg_1_pin_4_6
timestamp 1749560624
transform 1 0 32474 0 1 12573
box 1540 -22764 1864 -22616
use rseg_1_pin_4  rseg_1_pin_4_7
timestamp 1749560624
transform 1 0 34450 0 1 12573
box 1540 -22764 1864 -22616
use rseg_1_pin_4  rseg_1_pin_4_8
timestamp 1749560624
transform 1 0 37185 0 1 12573
box 1540 -22764 1864 -22616
use rseg_1_pin_5  rseg_1_pin_5_0
timestamp 1749563217
transform 1 0 25152 0 1 12573
box 1540 -22764 1952 -22615
use rseg_1_pin_5  rseg_1_pin_5_1
timestamp 1749563217
transform 1 0 30065 0 1 12573
box 1540 -22764 1952 -22615
use rseg_1_pin_5  rseg_1_pin_5_2
timestamp 1749563217
transform 1 0 34803 0 1 12573
box 1540 -22764 1952 -22615
use rseg_2_1  rseg_2_1_0
timestamp 1749485587
transform 1 0 18217 0 1 4094
box 4785 -17149 8535 -13951
use rseg_2_2  rseg_2_2_0
timestamp 1749485587
transform 1 0 16823 0 1 4958
box 9957 -18013 12354 -14815
use rseg_2_3  rseg_2_3_0
timestamp 1749485587
transform 1 0 15455 0 1 5171
box 13750 -18226 16210 -15028
use rseg_2_4  rseg_2_4_0
timestamp 1749369846
transform 1 0 18270 0 1 9878
box 13423 -22933 15713 -19735
use rseg_2_5  rseg_2_5_0
timestamp 1749369846
transform 1 0 16350 0 1 9986
box 17664 -23041 20052 -19843
use rseg_2_6  rseg_2_6_0
timestamp 1749369846
transform 1 0 14903 0 1 10179
box 21528 -23234 24146 -20036
<< labels >>
flabel metal2 s 22810 -10318 22810 -10318 0 FreeSans 1600 0 0 0 v0
port 0 nsew
flabel locali s 22846 -13211 22846 -13211 2 FreeSans 1600 0 0 0 gnd
port 49 ne
flabel metal1 s 23266 -10191 23266 -10191 2 FreeSans 480 0 0 0 v1
port 1 ne
flabel metal1 s 26428 -10191 26428 -10191 2 FreeSans 480 0 0 0 v2
port 2 ne
flabel metal1 s 23178 -10191 23178 -10191 2 FreeSans 320 0 0 0 v3
port 3 ne
flabel metal1 s 26516 -10191 26516 -10191 2 FreeSans 320 0 0 0 v4
port 4 ne
flabel metal1 s 23090 -10191 23090 -10191 2 FreeSans 320 0 0 0 v5
port 5 ne
flabel metal1 s 26604 -10191 26604 -10191 2 FreeSans 320 0 0 0 v6
port 6 ne
flabel metal1 s 23002 -10191 23002 -10191 2 FreeSans 320 0 0 0 v7
port 7 ne
flabel metal1 s 26692 -10191 26692 -10191 2 FreeSans 320 0 0 0 v8
port 8 ne
flabel metal1 s 26780 -10191 26780 -10191 2 FreeSans 320 0 0 0 v9
port 9 ne
flabel metal1 s 29117 -10191 29117 -10191 2 FreeSans 320 0 0 0 v10
port 10 ne
flabel metal1 s 26868 -10191 26868 -10191 2 FreeSans 320 0 0 0 v11
port 11 ne
flabel metal1 s 29029 -10191 29029 -10191 2 FreeSans 320 0 0 0 v12
port 12 ne
flabel metal1 s 26956 -10191 26956 -10191 2 FreeSans 320 0 0 0 v13
port 13 ne
flabel metal1 s 27044 -10191 27044 -10191 2 FreeSans 320 0 0 0 v15
port 15 ne
flabel metal1 s 28941 -10191 28941 -10191 2 FreeSans 320 0 0 0 v14
port 14 ne
flabel metal1 s 28853 -10191 28853 -10191 2 FreeSans 320 0 0 0 v16
port 16 ne
flabel metal1 s 29469 -10191 29469 -10191 2 FreeSans 160 0 0 0 v17
port 17 ne
flabel metal1 s 31341 -10191 31341 -10191 2 FreeSans 160 0 0 0 v18
port 18 ne
flabel metal1 s 29381 -10191 29381 -10191 2 FreeSans 240 0 0 0 v19
port 19 ne
flabel metal1 s 31429 -10191 31429 -10191 2 FreeSans 240 0 0 0 v20
port 20 ne
flabel metal1 s 29293 -10191 29293 -10191 2 FreeSans 240 0 0 0 v21
port 21 ne
flabel metal1 s 31517 -10191 31517 -10191 2 FreeSans 240 0 0 0 v22
port 22 ne
flabel metal1 s 29205 -10191 29205 -10191 2 FreeSans 240 0 0 0 v23
port 23 ne
flabel metal1 s 31605 -10191 31605 -10191 2 FreeSans 240 0 0 0 v24
port 24 ne
flabel metal1 s 31693 -10191 31693 -10191 2 FreeSans 240 0 0 0 v25
port 25 ne
flabel metal1 s 33923 -10191 33923 -10191 2 FreeSans 240 0 0 0 v26
port 26 ne
flabel metal1 s 31781 -10191 31781 -10191 2 FreeSans 240 0 0 0 v27
port 27 ne
flabel metal1 s 33835 -10191 33835 -10191 2 FreeSans 240 0 0 0 v28
port 28 ne
flabel metal1 s 31869 -10191 31869 -10191 2 FreeSans 240 0 0 0 v29
port 29 ne
flabel metal1 s 33747 -10191 33747 -10191 2 FreeSans 240 0 0 0 v30
port 30 ne
flabel metal1 s 31957 -10191 31957 -10191 2 FreeSans 240 0 0 0 v31
port 31 ne
flabel metal1 s 33659 -10191 33659 -10191 2 FreeSans 240 0 0 0 v32
port 32 ne
flabel metal1 s 34278 -10191 34278 -10191 2 FreeSans 240 0 0 0 v33
port 33 ne
flabel metal1 s 36078 -10191 36078 -10191 2 FreeSans 240 0 0 0 v34
port 34 ne
flabel metal1 s 34190 -10191 34190 -10191 2 FreeSans 240 0 0 0 v35
port 35 ne
flabel metal1 s 36166 -10191 36166 -10191 2 FreeSans 240 0 0 0 v36
port 36 ne
flabel metal1 s 34102 -10191 34102 -10191 2 FreeSans 240 0 0 0 v37
port 37 ne
flabel metal1 s 36254 -10191 36254 -10191 2 FreeSans 240 0 0 0 v38
port 38 ne
flabel metal1 s 34014 -10191 34014 -10191 2 FreeSans 240 0 0 0 v39
port 39 ne
flabel metal1 s 36342 -10191 36342 -10191 2 FreeSans 240 0 0 0 v40
port 40 ne
flabel metal1 s 36431 -10191 36431 -10191 2 FreeSans 240 0 0 0 v41
port 41 ne
flabel metal1 s 38989 -10191 38989 -10191 2 FreeSans 240 0 0 0 v42
port 42 ne
flabel metal1 s 36519 -10191 36519 -10191 2 FreeSans 240 0 0 0 v43
port 43 ne
flabel metal1 s 38901 -10191 38901 -10191 2 FreeSans 240 0 0 0 v44
port 44 ne
flabel metal1 s 36607 -10191 36607 -10191 2 FreeSans 240 0 0 0 v45
port 45 ne
flabel metal1 s 38813 -10191 38813 -10191 2 FreeSans 240 0 0 0 v46
port 46 ne
flabel metal1 s 36695 -10191 36695 -10191 2 FreeSans 240 0 0 0 v47
port 47 ne
flabel metal1 s 38725 -10191 38725 -10191 2 FreeSans 240 0 0 0 v48
port 48 ne
<< end >>
