magic
tech sky130A
magscale 1 2
timestamp 1750197143
<< pwell >>
rect -758 -287 758 287
<< mvnmos >>
rect -530 -91 530 29
<< mvndiff >>
rect -588 17 -530 29
rect -588 -79 -576 17
rect -542 -79 -530 17
rect -588 -91 -530 -79
rect 530 17 588 29
rect 530 -79 542 17
rect 576 -79 588 17
rect 530 -91 588 -79
<< mvndiffc >>
rect -576 -79 -542 17
rect 542 -79 576 17
<< mvpsubdiff >>
rect -722 239 722 251
rect -722 205 -614 239
rect 614 205 722 239
rect -722 193 722 205
rect -722 143 -664 193
rect -722 -143 -710 143
rect -676 -143 -664 143
rect 664 143 722 193
rect -722 -193 -664 -143
rect 664 -143 676 143
rect 710 -143 722 143
rect 664 -193 722 -143
rect -722 -205 722 -193
rect -722 -239 -614 -205
rect 614 -239 722 -205
rect -722 -251 722 -239
<< mvpsubdiffcont >>
rect -614 205 614 239
rect -710 -143 -676 143
rect 676 -143 710 143
rect -614 -239 614 -205
<< poly >>
rect -530 101 530 117
rect -530 67 -514 101
rect 514 67 530 101
rect -530 29 530 67
rect -530 -117 530 -91
<< polycont >>
rect -514 67 514 101
<< locali >>
rect -710 205 -614 239
rect 614 205 710 239
rect -710 143 -676 205
rect 676 143 710 205
rect -530 67 -514 101
rect 514 67 530 101
rect -576 17 -542 33
rect -576 -95 -542 -79
rect 542 17 576 33
rect 542 -95 576 -79
rect -710 -205 -676 -143
rect 676 -205 710 -143
rect -710 -239 -614 -205
rect 614 -239 710 -205
<< viali >>
rect -386 67 386 101
rect -576 -79 -542 17
rect 542 -79 576 17
<< metal1 >>
rect -398 101 398 107
rect -398 67 -386 101
rect 386 67 398 101
rect -398 61 398 67
rect -582 17 -536 29
rect -582 -79 -576 17
rect -542 -79 -536 17
rect -582 -91 -536 -79
rect 536 17 582 29
rect 536 -79 542 17
rect 576 -79 582 17
rect 536 -91 582 -79
<< properties >>
string FIXED_BBOX -693 -222 693 222
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.6 l 5.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
