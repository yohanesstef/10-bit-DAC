magic
tech sky130A
magscale 1 2
timestamp 1749057406
<< pwell >>
rect -307 -940 307 940
<< psubdiff >>
rect -271 870 -175 904
rect 175 870 271 904
rect -271 808 -237 870
rect 237 808 271 870
rect -271 -870 -237 -808
rect 237 -870 271 -808
rect -271 -904 -175 -870
rect 175 -904 271 -870
<< psubdiffcont >>
rect -175 870 175 904
rect -271 -808 -237 808
rect 237 -808 271 808
rect -175 -904 175 -870
<< xpolycontact >>
rect -141 342 141 774
rect -141 -774 141 -342
<< xpolyres >>
rect -141 -342 141 342
<< locali >>
rect -271 870 -175 904
rect 175 870 271 904
rect -271 808 -237 870
rect 237 808 271 870
rect -271 -870 -237 -808
rect 237 -870 271 -808
rect -271 -904 -175 -870
rect 175 -904 271 -870
<< viali >>
rect -125 359 125 756
rect -125 -756 125 -359
<< metal1 >>
rect -131 756 131 768
rect -131 359 -125 756
rect 125 359 131 756
rect -131 347 131 359
rect -131 -359 131 -347
rect -131 -756 -125 -359
rect 125 -756 131 -359
rect -131 -768 131 -756
<< properties >>
string FIXED_BBOX -254 -887 254 887
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 3.578 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 5.342k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
