magic
tech sky130A
magscale 1 2
timestamp 1750156376
<< error_s >>
rect -4651 4964 4758 5030
rect -4651 3650 -4585 4964
rect -4525 4885 4632 4904
rect -4525 4505 -4446 4885
rect -4410 4505 -4380 4785
rect 4486 4505 4516 4785
rect 4552 4505 4632 4885
rect -4525 4359 4632 4505
rect -4525 4255 -4459 4359
rect 4566 4255 4632 4359
rect -4525 4251 4632 4255
rect -4525 3729 -4446 4251
rect -4410 4185 -4094 4189
rect -4034 4185 4140 4189
rect 4200 4185 4516 4189
rect -4410 3829 -4380 4185
rect 4486 3829 4516 4185
rect 4552 3729 4632 4251
rect -4525 3710 4632 3729
rect 4692 3650 4758 4964
rect -4651 3584 4758 3650
<< metal1 >>
rect -4497 4397 -4437 4872
rect 4544 4866 4604 4872
rect -217 4425 -211 4485
rect -151 4425 -4 4485
rect 111 4425 258 4485
rect 318 4425 324 4485
rect -4028 4397 -3982 4425
rect 4088 4397 4134 4425
rect 4544 4397 4604 4806
rect -4497 4337 -91 4397
rect 198 4337 4604 4397
rect -4028 4217 -91 4277
rect 198 4217 4134 4277
rect -4028 4189 -3982 4217
rect 4088 4189 4134 4217
rect -217 4129 -211 4189
rect -151 4129 258 4189
rect 318 4129 324 4189
rect 4544 3808 4604 4337
rect 4544 3742 4604 3748
<< via1 >>
rect 4544 4806 4604 4866
rect -211 4425 -151 4485
rect 258 4425 318 4485
rect -211 4129 -151 4189
rect 258 4129 318 4189
rect 4544 3748 4604 3808
<< metal2 >>
rect 4604 4806 4610 4866
rect -211 4485 -151 4491
rect -211 4189 -151 4425
rect -211 4123 -151 4129
rect 258 4485 318 4491
rect 258 4189 318 4425
rect 258 4123 318 4129
rect 4604 3748 4610 3808
use cm_pcell3_2  cm_pcell3_2_0
timestamp 1750156376
transform 1 0 -4083 0 1 4367
box -568 -126 8841 663
use cm_pcell3_2  cm_pcell3_2_1
timestamp 1750156376
transform 1 0 -4083 0 -1 4247
box -568 -126 8841 663
use cross_pair  cross_pair_0
timestamp 1750150351
transform 1 0 -36205 0 1 2362
box 36114 1855 36403 2035
<< end >>
