magic
tech sky130A
magscale 1 2
timestamp 1750847318
<< error_p >>
rect -144 446 144 480
rect -174 231 174 446
rect -144 197 144 231
rect -174 -18 174 197
rect -144 -52 144 -18
rect -174 -267 174 -52
rect -174 -513 -144 -301
rect -108 -447 -78 -367
rect 78 -447 108 -367
rect -108 -451 108 -447
rect 144 -513 174 -301
rect -174 -517 174 -513
<< nwell >>
rect -144 234 144 480
rect -144 -15 144 231
rect -144 -264 144 -18
rect -144 -513 144 -267
<< mvpmos >>
rect -50 296 50 380
rect -50 47 50 131
rect -50 -202 50 -118
rect -50 -451 50 -367
<< mvpdiff >>
rect -108 368 -50 380
rect -108 308 -96 368
rect -62 308 -50 368
rect -108 296 -50 308
rect 50 368 108 380
rect 50 308 62 368
rect 96 308 108 368
rect 50 296 108 308
rect -108 119 -50 131
rect -108 59 -96 119
rect -62 59 -50 119
rect -108 47 -50 59
rect 50 119 108 131
rect 50 59 62 119
rect 96 59 108 119
rect 50 47 108 59
rect -108 -130 -50 -118
rect -108 -190 -96 -130
rect -62 -190 -50 -130
rect -108 -202 -50 -190
rect 50 -130 108 -118
rect 50 -190 62 -130
rect 96 -190 108 -130
rect 50 -202 108 -190
rect -108 -379 -50 -367
rect -108 -439 -96 -379
rect -62 -439 -50 -379
rect -108 -451 -50 -439
rect 50 -379 108 -367
rect 50 -439 62 -379
rect 96 -439 108 -379
rect 50 -451 108 -439
<< mvpdiffc >>
rect -96 308 -62 368
rect 62 308 96 368
rect -96 59 -62 119
rect 62 59 96 119
rect -96 -190 -62 -130
rect 62 -190 96 -130
rect -96 -439 -62 -379
rect 62 -439 96 -379
<< poly >>
rect -50 461 50 477
rect -50 427 -34 461
rect 34 427 50 461
rect -50 380 50 427
rect -50 270 50 296
rect -50 212 50 228
rect -50 178 -34 212
rect 34 178 50 212
rect -50 131 50 178
rect -50 21 50 47
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -228 50 -202
rect -50 -286 50 -270
rect -50 -320 -34 -286
rect 34 -320 50 -286
rect -50 -367 50 -320
rect -50 -477 50 -451
<< polycont >>
rect -34 427 34 461
rect -34 178 34 212
rect -34 -71 34 -37
rect -34 -320 34 -286
<< locali >>
rect -50 427 -34 461
rect 34 427 50 461
rect -96 368 -62 384
rect -96 292 -62 308
rect 62 368 96 384
rect 62 292 96 308
rect -50 178 -34 212
rect 34 178 50 212
rect -96 119 -62 135
rect -96 43 -62 59
rect 62 119 96 135
rect 62 43 96 59
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -206 -62 -190
rect 62 -130 96 -114
rect 62 -206 96 -190
rect -50 -320 -34 -286
rect 34 -320 50 -286
rect -96 -379 -62 -363
rect -96 -455 -62 -439
rect 62 -379 96 -363
rect 62 -455 96 -439
<< viali >>
rect -26 427 26 461
rect -96 308 -62 368
rect 62 308 96 368
rect -26 178 26 212
rect -96 59 -62 119
rect 62 59 96 119
rect -26 -71 26 -37
rect -96 -190 -62 -130
rect 62 -190 96 -130
rect -26 -320 26 -286
rect -96 -439 -62 -379
rect 62 -439 96 -379
<< metal1 >>
rect -38 461 38 467
rect -38 427 -26 461
rect 26 427 38 461
rect -38 421 38 427
rect -102 368 -56 380
rect -102 308 -96 368
rect -62 308 -56 368
rect -102 296 -56 308
rect 56 368 102 380
rect 56 308 62 368
rect 96 308 102 368
rect 56 296 102 308
rect -38 212 38 218
rect -38 178 -26 212
rect 26 178 38 212
rect -38 172 38 178
rect -102 119 -56 131
rect -102 59 -96 119
rect -62 59 -56 119
rect -102 47 -56 59
rect 56 119 102 131
rect 56 59 62 119
rect 96 59 102 119
rect 56 47 102 59
rect -38 -37 38 -31
rect -38 -71 -26 -37
rect 26 -71 38 -37
rect -38 -77 38 -71
rect -102 -130 -56 -118
rect -102 -190 -96 -130
rect -62 -190 -56 -130
rect -102 -202 -56 -190
rect 56 -130 102 -118
rect 56 -190 62 -130
rect 96 -190 102 -130
rect 56 -202 102 -190
rect -38 -286 38 -280
rect -38 -320 -26 -286
rect 26 -320 38 -286
rect -38 -326 38 -320
rect -102 -379 -56 -367
rect -102 -439 -96 -379
rect -62 -439 -56 -379
rect -102 -451 -56 -439
rect 56 -379 102 -367
rect 56 -439 62 -379
rect 96 -439 102 -379
rect 56 -451 102 -439
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 0.50 m 4 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
