magic
tech sky130A
magscale 1 2
timestamp 1750060524
<< error_s >>
rect 1159 868 1165 874
rect 1213 868 1219 874
rect 2663 868 2669 874
rect 2717 868 2723 874
rect 1153 862 1159 868
rect 1219 862 1225 868
rect 2657 862 2663 868
rect 2723 862 2729 868
rect 1153 808 1159 814
rect 1219 808 1225 814
rect 2657 808 2663 814
rect 2723 808 2729 814
rect 1159 802 1165 808
rect 1213 802 1219 808
rect 2663 802 2669 808
rect 2717 802 2723 808
rect 407 692 413 698
rect 461 692 467 698
rect 1911 692 1917 698
rect 1965 692 1971 698
rect 401 686 407 692
rect 467 686 473 692
rect 1905 686 1911 692
rect 1971 686 1977 692
rect 401 632 407 638
rect 467 632 473 638
rect 1905 632 1911 638
rect 1971 632 1977 638
rect 407 626 413 632
rect 461 626 467 632
rect 1911 626 1917 632
rect 1965 626 1971 632
rect 783 516 789 522
rect 837 516 843 522
rect 777 510 783 516
rect 843 510 849 516
rect 777 456 783 462
rect 843 456 849 462
rect 783 450 789 456
rect 837 450 843 456
rect 1535 428 1541 434
rect 1589 428 1595 434
rect 1529 422 1535 428
rect 1595 422 1601 428
rect 1529 368 1535 374
rect 1595 368 1601 374
rect 1535 362 1541 368
rect 1589 362 1595 368
<< metal1 >>
rect 1153 808 1159 868
rect 1219 808 1225 868
rect 2657 808 2663 868
rect 2723 808 2729 868
rect 1159 702 1219 808
rect 2663 632 2723 808
rect 2491 604 2775 632
rect 777 456 783 516
rect 843 456 849 516
rect 2491 456 2519 604
rect 2663 582 2723 604
rect 2235 428 2519 456
<< via1 >>
rect 1159 808 1219 868
rect 2663 808 2723 868
rect 407 632 467 692
rect 1911 632 1971 692
rect 783 456 843 516
rect 1535 368 1595 428
use cm_ncell1_cell  cm_ncell1_cell_0
timestamp 1750060524
transform 1 0 -9 0 1 0
box -12 -4 3580 1064
<< end >>
