magic
tech sky130A
magscale 1 2
timestamp 1751021419
<< metal1 >>
rect 13975 16863 14035 17640
rect 15217 16951 15277 17632
rect 15217 16885 15277 16891
rect 16314 16951 16374 16957
rect 13975 16797 14035 16803
rect 16072 16863 16132 16869
rect 16072 13025 16132 16803
rect 16072 12959 16132 12965
rect 16187 13377 16247 13383
rect 16187 6636 16247 13317
rect 16314 13113 16374 16891
rect 16314 13047 16374 13053
rect 16471 12937 16531 17646
rect 16471 12871 16531 12877
rect 16787 13465 16847 13471
rect 16787 8083 16847 13405
rect 17327 12849 17387 17646
rect 17327 12783 17387 12789
rect 17467 12761 17527 12767
rect 16781 8031 16787 8083
rect 16847 8031 16853 8083
rect 17467 8060 17527 12701
rect 18173 12761 18233 17645
rect 18173 12695 18233 12701
rect 18764 12673 18824 17646
rect 20660 13993 20720 17092
rect 20660 13927 20720 13933
rect 21240 13905 21300 17092
rect 21240 13839 21300 13845
rect 21820 13817 21880 17092
rect 21820 13751 21880 13757
rect 22400 13729 22460 17092
rect 23654 14081 23714 17092
rect 25062 14345 25122 17092
rect 25062 14279 25122 14285
rect 26470 14257 26530 17092
rect 26470 14191 26530 14197
rect 27878 14169 27938 17092
rect 31892 14433 31952 19133
rect 31892 14367 31952 14373
rect 27878 14103 27938 14109
rect 23654 14015 23714 14021
rect 22400 13663 22460 13669
rect 31468 13817 31528 13823
rect 18764 12607 18824 12613
rect 22995 12673 23055 12679
rect 19967 12585 20027 12591
rect 19122 12409 19182 12415
rect 18543 12321 18603 12327
rect 18239 12233 18299 12239
rect 17938 12145 17998 12151
rect 17938 9141 17998 12085
rect 18239 9141 18299 12173
rect 18543 9142 18603 12261
rect 19122 9144 19182 12349
rect 19967 9143 20027 12525
rect 21112 12497 21172 12503
rect 21112 9141 21172 12437
rect 22995 8062 23055 12613
rect 31468 8086 31528 13757
rect 37333 12761 37393 12767
rect 32093 12673 32153 12679
rect 31462 8026 31468 8086
rect 31528 8026 31534 8086
rect 32093 8056 32153 12613
rect 36213 12585 36273 12591
rect 35068 12497 35128 12503
rect 33644 12409 33704 12415
rect 33039 12233 33099 12239
rect 33039 9132 33099 12173
rect 33340 12145 33400 12151
rect 33340 9132 33400 12085
rect 33644 9133 33704 12349
rect 34223 12321 34283 12327
rect 34223 9136 34283 12261
rect 35068 9134 35128 12437
rect 36213 9132 36273 12525
rect 37333 8071 37393 12701
rect 16781 7587 16787 7639
rect 16847 7587 16853 7639
rect 16187 6578 16247 6584
rect 16787 6636 16847 7587
rect 31462 7586 31468 7646
rect 31528 7586 31534 7646
rect 31468 6645 31528 7586
rect 31468 6593 31763 6645
rect 16787 6578 16847 6584
<< via1 >>
rect 15217 16891 15277 16951
rect 16314 16891 16374 16951
rect 13975 16803 14035 16863
rect 16072 16803 16132 16863
rect 16072 12965 16132 13025
rect 16187 13317 16247 13377
rect 16314 13053 16374 13113
rect 16471 12877 16531 12937
rect 16787 13405 16847 13465
rect 17327 12789 17387 12849
rect 17467 12701 17527 12761
rect 16787 8031 16847 8083
rect 18173 12701 18233 12761
rect 20660 13933 20720 13993
rect 21240 13845 21300 13905
rect 21820 13757 21880 13817
rect 25062 14285 25122 14345
rect 26470 14197 26530 14257
rect 31892 14373 31952 14433
rect 27878 14109 27938 14169
rect 23654 14021 23714 14081
rect 22400 13669 22460 13729
rect 31468 13757 31528 13817
rect 18764 12613 18824 12673
rect 22995 12613 23055 12673
rect 19967 12525 20027 12585
rect 19122 12349 19182 12409
rect 18543 12261 18603 12321
rect 18239 12173 18299 12233
rect 17938 12085 17998 12145
rect 21112 12437 21172 12497
rect 37333 12701 37393 12761
rect 32093 12613 32153 12673
rect 31468 8026 31528 8086
rect 36213 12525 36273 12585
rect 35068 12437 35128 12497
rect 33644 12349 33704 12409
rect 33039 12173 33099 12233
rect 33340 12085 33400 12145
rect 34223 12261 34283 12321
rect 16787 7587 16847 7639
rect 16187 6584 16247 6636
rect 31468 7586 31528 7646
rect 16787 6584 16847 6636
<< metal2 >>
rect -1386 25030 49223 25630
rect -1386 24330 48523 24930
rect -1386 23630 47823 24230
rect 18478 20374 18616 20636
rect 21430 19079 21440 19135
rect 21496 19079 21506 19135
rect 26262 19079 26272 19135
rect 26328 19079 26338 19135
rect 15886 18762 15896 18818
rect 15952 18762 15962 18818
rect 18405 18762 18415 18818
rect 18471 18762 18481 18818
rect 15211 16891 15217 16951
rect 15277 16891 16314 16951
rect 16374 16891 16380 16951
rect 13969 16803 13975 16863
rect 14035 16803 16072 16863
rect 16132 16803 16138 16863
rect 21430 14551 21440 14607
rect 21496 14551 21506 14607
rect 26263 14463 26273 14519
rect 26329 14463 26339 14519
rect 38148 13936 38158 13992
rect 38214 13936 38224 13992
rect 34815 13845 34825 13901
rect 34881 13845 34891 13901
rect 23482 13583 23492 13639
rect 23548 13583 23558 13639
rect 20149 13495 20159 13551
rect 20215 13495 20225 13551
rect 15886 13231 15896 13287
rect 15952 13231 15962 13287
rect 18405 13143 18415 13199
rect 18471 13143 18481 13199
rect 12084 11997 15856 12057
rect 12084 11909 15856 11969
rect 12084 11821 15856 11881
rect 12084 11733 15856 11793
rect 16781 8031 16787 8083
rect 16847 8031 16853 8083
rect 16787 7639 16847 8031
rect 31462 8026 31468 8086
rect 31528 8026 31534 8086
rect 31468 7646 31528 8026
rect 16781 7587 16787 7639
rect 16847 7587 16853 7639
rect 31462 7586 31468 7646
rect 31528 7586 31534 7646
rect 16078 6584 16187 6636
rect 16247 6584 16253 6636
rect 16781 6584 16787 6636
rect 16847 6584 17024 6636
rect 20147 6584 20157 6640
rect 20213 6584 20223 6640
rect 23482 6584 23492 6640
rect 23548 6584 23558 6640
rect 34818 6591 34828 6647
rect 34884 6645 34894 6647
rect 34884 6593 35057 6645
rect 34884 6591 34894 6593
rect 38151 6591 38161 6647
rect 38217 6591 38227 6647
rect 47223 987 47823 23630
rect -916 387 47823 987
rect 47923 287 48523 24330
rect -916 -313 48523 287
rect 48623 -413 49223 25030
rect -916 -1013 49223 -413
<< via2 >>
rect 13850 20385 14009 20626
rect 34162 20383 34535 20626
rect 21440 19079 21496 19135
rect 26272 19079 26328 19135
rect 15896 18762 15952 18818
rect 18415 18762 18471 18818
rect 21440 14551 21496 14607
rect 26273 14463 26329 14519
rect 38158 13936 38214 13992
rect 34825 13845 34881 13901
rect 23492 13583 23548 13639
rect 20159 13495 20215 13551
rect 15896 13231 15952 13287
rect 18415 13143 18471 13199
rect 20157 6584 20213 6640
rect 23492 6584 23548 6640
rect 34828 6591 34884 6647
rect 38161 6591 38217 6647
rect 13764 3987 13895 4236
rect 39860 3981 39997 4234
<< metal3 >>
rect 13838 20626 17211 20636
rect 13838 20385 13850 20626
rect 14009 20385 17211 20626
rect 13838 20374 17211 20385
rect 15891 18818 15957 18828
rect 15891 18762 15896 18818
rect 15952 18762 15957 18818
rect 15891 18752 15957 18762
rect 15894 13297 15954 18752
rect 15891 13287 15957 13297
rect 15891 13231 15896 13287
rect 15952 13231 15957 13287
rect 15891 13221 15957 13231
rect 16811 4242 17211 20374
rect 34150 20626 34550 20636
rect 34150 20383 34162 20626
rect 34535 20383 34550 20626
rect 21435 19135 21501 19145
rect 21435 19079 21440 19135
rect 21496 19079 21501 19135
rect 21435 19069 21501 19079
rect 26267 19135 26333 19145
rect 26267 19079 26272 19135
rect 26328 19079 26333 19135
rect 26267 19069 26333 19079
rect 18410 18818 18476 18828
rect 18410 18762 18415 18818
rect 18471 18762 18476 18818
rect 18410 18752 18476 18762
rect 18413 17617 18473 18752
rect 18413 14343 18474 17617
rect 21438 14617 21498 19069
rect 21435 14607 21501 14617
rect 21435 14551 21440 14607
rect 21496 14551 21501 14607
rect 21435 14541 21501 14551
rect 26271 14529 26331 19069
rect 26268 14519 26334 14529
rect 26268 14463 26273 14519
rect 26329 14463 26334 14519
rect 26268 14453 26334 14463
rect 18413 13209 18473 14343
rect 23487 13639 23553 13649
rect 23487 13583 23492 13639
rect 23548 13583 23553 13639
rect 23487 13573 23553 13583
rect 20154 13551 20220 13561
rect 20154 13495 20159 13551
rect 20215 13495 20220 13551
rect 20154 13485 20220 13495
rect 18410 13199 18476 13209
rect 18410 13143 18415 13199
rect 18471 13143 18476 13199
rect 18410 13133 18476 13143
rect 20157 6650 20217 13485
rect 23490 6650 23550 13573
rect 20152 6640 20218 6650
rect 20152 6584 20157 6640
rect 20213 6584 20218 6640
rect 20152 6574 20218 6584
rect 23487 6640 23553 6650
rect 23487 6584 23492 6640
rect 23548 6584 23553 6640
rect 23487 6574 23553 6584
rect 13756 4236 17211 4242
rect 13756 3987 13764 4236
rect 13895 3987 17211 4236
rect 13756 3980 17211 3987
rect 34150 4242 34550 20383
rect 38153 13992 38219 14002
rect 38153 13936 38158 13992
rect 38214 13936 38219 13992
rect 38153 13926 38219 13936
rect 34820 13901 34886 13911
rect 34820 13845 34825 13901
rect 34881 13845 34886 13901
rect 34820 13835 34886 13845
rect 34823 6657 34883 13835
rect 38156 6657 38216 13926
rect 34823 6647 34889 6657
rect 34823 6591 34828 6647
rect 34884 6591 34889 6647
rect 34823 6581 34889 6591
rect 38156 6647 38222 6657
rect 38156 6591 38161 6647
rect 38217 6591 38222 6647
rect 38156 6581 38222 6591
rect 34150 4234 40015 4242
rect 34150 3981 39860 4234
rect 39997 3981 40015 4234
rect 34150 3970 40015 3981
<< comment >>
rect -916 1083 -816 1087
use grid_ys_0p14_yr_0p3  grid_ys_0p14_yr_0p3_0
timestamp 1749886903
transform 1 0 36789 0 1 5069
box 1801 3053 3589 4841
use top_dcell_routing  top_dcell_routing_0
timestamp 1750900893
transform 1 0 0 0 1 0
box 15856 1202 46831 23447
use top_opamp_n_final_switch  top_opamp_n_final_switch_0
timestamp 1751021419
transform 1 0 1407 0 1 401
box -2676 876 13894 23072
use top_segment_1  top_segment_1_0
timestamp 1750900893
transform 1 0 26106 0 1 1210
box -385 -24 14453 8429
use top_segment_2  top_segment_2_0
timestamp 1750900893
transform -1 0 34310 0 -1 23469
box -727 39 15704 7051
use top_segment_3  top_segment_3_0
timestamp 1749552768
transform -1 0 24112 0 -1 23696
box 5007 266 11251 6636
use top_segment_4  top_segment_4_1
timestamp 1749664768
transform 1 0 -17367 0 1 13412
box 29493 -12226 43322 -3773
<< end >>
