magic
tech sky130A
magscale 1 2
timestamp 1750060524
<< metal1 >>
rect -98 24 66 426
rect 278 24 442 144
rect 654 24 818 426
rect 1030 24 1194 144
rect 1406 24 1570 144
rect 278 -482 442 -80
rect 654 -200 818 -80
rect 1030 -482 1194 -80
rect 1406 -200 1570 -80
use cm_ncell1_4  cm_ncell1_4_0
timestamp 1750060524
transform 1 0 -5 0 1 -57
box -11 55 1493 563
use cm_ncell1_4  cm_ncell1_4_1
timestamp 1750060524
transform 1 0 -5 0 -1 1
box -11 55 1493 563
<< end >>
