magic
tech sky130A
magscale 1 2
timestamp 1749896124
<< error_s >>
rect 912 1711 918 1717
rect 966 1711 972 1717
rect 1554 1711 1560 1717
rect 1608 1711 1614 1717
rect 2416 1711 2422 1717
rect 2470 1711 2476 1717
rect 3058 1711 3064 1717
rect 3112 1711 3118 1717
rect 3920 1711 3926 1717
rect 3974 1711 3980 1717
rect 4562 1711 4568 1717
rect 4616 1711 4622 1717
rect 906 1705 912 1711
rect 972 1705 978 1711
rect 1548 1705 1554 1711
rect 1614 1705 1620 1711
rect 2410 1705 2416 1711
rect 2476 1705 2482 1711
rect 3052 1705 3058 1711
rect 3118 1705 3124 1711
rect 3914 1705 3920 1711
rect 3980 1705 3986 1711
rect 4556 1705 4562 1711
rect 4622 1705 4628 1711
rect 906 1651 912 1657
rect 972 1651 978 1657
rect 1548 1651 1554 1657
rect 1614 1651 1620 1657
rect 2410 1651 2416 1657
rect 2476 1651 2482 1657
rect 3052 1651 3058 1657
rect 3118 1651 3124 1657
rect 3914 1651 3920 1657
rect 3980 1651 3986 1657
rect 4556 1651 4562 1657
rect 4622 1651 4628 1657
rect 912 1645 918 1651
rect 966 1645 972 1651
rect 1554 1645 1560 1651
rect 1608 1645 1614 1651
rect 2416 1645 2422 1651
rect 2470 1645 2476 1651
rect 3058 1645 3064 1651
rect 3112 1645 3118 1651
rect 3920 1645 3926 1651
rect 3974 1645 3980 1651
rect 4562 1645 4568 1651
rect 4616 1645 4622 1651
rect 1664 1623 1670 1629
rect 1718 1623 1724 1629
rect 2306 1623 2312 1629
rect 2360 1623 2366 1629
rect 3168 1623 3174 1629
rect 3222 1623 3228 1629
rect 3810 1623 3816 1629
rect 3864 1623 3870 1629
rect 1658 1617 1664 1623
rect 1724 1617 1730 1623
rect 2300 1617 2306 1623
rect 2366 1617 2372 1623
rect 3162 1617 3168 1623
rect 3228 1617 3234 1623
rect 3804 1617 3810 1623
rect 3870 1617 3876 1623
rect 1658 1563 1664 1569
rect 1724 1563 1730 1569
rect 2300 1563 2306 1569
rect 2366 1563 2372 1569
rect 3162 1563 3168 1569
rect 3228 1563 3234 1569
rect 3804 1563 3810 1569
rect 3870 1563 3876 1569
rect 1664 1557 1670 1563
rect 1718 1557 1724 1563
rect 2306 1557 2312 1563
rect 2360 1557 2366 1563
rect 3168 1557 3174 1563
rect 3222 1557 3228 1563
rect 3810 1557 3816 1563
rect 3864 1557 3870 1563
rect 1233 1447 1239 1453
rect 1287 1447 1293 1453
rect 2737 1447 2743 1453
rect 2791 1447 2797 1453
rect 4241 1447 4247 1453
rect 4295 1447 4301 1453
rect 1227 1441 1233 1447
rect 1293 1441 1299 1447
rect 2731 1441 2737 1447
rect 2797 1441 2803 1447
rect 4235 1441 4241 1447
rect 4301 1441 4307 1447
rect 1227 1387 1233 1393
rect 1293 1387 1299 1393
rect 2731 1387 2737 1393
rect 2797 1387 2803 1393
rect 4235 1387 4241 1393
rect 4301 1387 4307 1393
rect 1233 1381 1239 1387
rect 1287 1381 1293 1387
rect 2737 1381 2743 1387
rect 2791 1381 2797 1387
rect 4241 1381 4247 1387
rect 4295 1381 4301 1387
rect 1985 1359 1991 1365
rect 2039 1359 2045 1365
rect 3489 1359 3495 1365
rect 3543 1359 3549 1365
rect 1979 1353 1985 1359
rect 2045 1353 2051 1359
rect 3483 1353 3489 1359
rect 3549 1353 3555 1359
rect 1979 1299 1985 1305
rect 2045 1299 2051 1305
rect 3483 1299 3489 1305
rect 3549 1299 3555 1305
rect 1985 1293 1991 1299
rect 2039 1293 2045 1299
rect 3489 1293 3495 1299
rect 3543 1293 3549 1299
rect 4387 1183 4393 1189
rect 4441 1183 4447 1189
rect 4381 1177 4387 1183
rect 4447 1177 4453 1183
rect 4381 1123 4387 1129
rect 4447 1123 4453 1129
rect 4387 1117 4393 1123
rect 4441 1117 4447 1123
rect 4558 1007 4564 1013
rect 4612 1007 4618 1013
rect 4552 1001 4558 1007
rect 4618 1001 4624 1007
rect 4552 947 4558 953
rect 4618 947 4624 953
rect 4558 941 4564 947
rect 4612 941 4618 947
rect 2044 831 2050 837
rect 2098 831 2104 837
rect 2678 831 2684 837
rect 2732 831 2738 837
rect 2038 825 2044 831
rect 2104 825 2110 831
rect 2672 825 2678 831
rect 2738 825 2744 831
rect 2038 771 2044 777
rect 2104 771 2110 777
rect 2672 771 2678 777
rect 2738 771 2744 777
rect 2044 765 2050 771
rect 2098 765 2104 771
rect 2678 765 2684 771
rect 2732 765 2738 771
rect 2361 655 2367 661
rect 2415 655 2421 661
rect 2355 649 2361 655
rect 2421 649 2427 655
rect 2355 595 2361 601
rect 2421 595 2427 601
rect 2361 589 2367 595
rect 2415 589 2421 595
rect 3865 567 3871 573
rect 3919 567 3925 573
rect 3859 561 3865 567
rect 3925 561 3931 567
rect 3859 507 3865 513
rect 3925 507 3931 513
rect 3865 501 3871 507
rect 3919 501 3925 507
rect 916 479 922 485
rect 970 479 976 485
rect 1609 479 1615 485
rect 1663 479 1669 485
rect 3113 479 3119 485
rect 3167 479 3173 485
rect 910 473 916 479
rect 976 473 982 479
rect 1603 473 1609 479
rect 1669 473 1675 479
rect 3107 473 3113 479
rect 3173 473 3179 479
rect 910 419 916 425
rect 976 419 982 425
rect 1603 419 1609 425
rect 1669 419 1675 425
rect 3107 419 3113 425
rect 3173 419 3179 425
rect 916 413 922 419
rect 970 413 976 419
rect 1609 413 1615 419
rect 1663 413 1669 419
rect 3113 413 3119 419
rect 3167 413 3173 419
rect 1178 303 1184 309
rect 1232 303 1238 309
rect 1288 303 1294 309
rect 1342 303 1348 309
rect 1930 303 1936 309
rect 1984 303 1990 309
rect 2792 303 2798 309
rect 2846 303 2852 309
rect 3434 303 3440 309
rect 3488 303 3494 309
rect 1172 297 1178 303
rect 1238 297 1244 303
rect 1282 297 1288 303
rect 1348 297 1354 303
rect 1924 297 1930 303
rect 1990 297 1996 303
rect 2786 297 2792 303
rect 2852 297 2858 303
rect 3428 297 3434 303
rect 3494 297 3500 303
rect 1172 243 1178 249
rect 1238 243 1244 249
rect 1282 243 1288 249
rect 1348 243 1354 249
rect 1924 243 1930 249
rect 1990 243 1996 249
rect 2786 243 2792 249
rect 2852 243 2858 249
rect 3428 243 3434 249
rect 3494 243 3500 249
rect 1178 237 1184 243
rect 1232 237 1238 243
rect 1288 237 1294 243
rect 1342 237 1348 243
rect 1930 237 1936 243
rect 1984 237 1990 243
rect 2792 237 2798 243
rect 2846 237 2852 243
rect 3434 237 3440 243
rect 3488 237 3494 243
rect 3544 215 3550 221
rect 3598 215 3604 221
rect 4186 215 4192 221
rect 4240 215 4246 221
rect 3538 209 3544 215
rect 3604 209 3610 215
rect 4180 209 4186 215
rect 4246 209 4252 215
rect 3538 155 3544 161
rect 3604 155 3610 161
rect 4180 155 4186 161
rect 4246 155 4252 161
rect 3544 149 3550 155
rect 3598 149 3604 155
rect 4186 149 4192 155
rect 4240 149 4246 155
<< metal1 >>
rect 906 1651 912 1711
rect 972 1651 978 1711
rect 1548 1651 1554 1711
rect 1614 1651 1620 1711
rect 2410 1651 2416 1711
rect 2476 1651 2482 1711
rect 3052 1651 3058 1711
rect 3118 1651 3124 1711
rect 3914 1651 3920 1711
rect 3980 1651 3986 1711
rect 4556 1651 4562 1711
rect 4622 1651 4628 1711
rect 912 1130 972 1651
rect 1181 1387 1233 1447
rect 1293 1387 1345 1447
rect 1554 1130 1614 1651
rect 1658 1563 1664 1623
rect 1724 1563 1730 1623
rect 2300 1563 2306 1623
rect 2366 1563 2372 1623
rect 1664 1130 1724 1563
rect 2306 1130 2366 1563
rect 2416 1130 2476 1651
rect 3058 1130 3118 1651
rect 3162 1563 3168 1623
rect 3228 1563 3234 1623
rect 3804 1563 3810 1623
rect 3870 1563 3876 1623
rect 3168 1130 3228 1563
rect 3810 1130 3870 1563
rect 3920 1130 3980 1651
rect 4381 1123 4387 1183
rect 4447 1123 4453 1183
rect 4562 1130 4622 1651
rect 2038 771 2044 831
rect 2104 771 2110 831
rect 2672 772 2678 831
rect 2738 772 2744 831
rect 910 419 916 479
rect 976 419 982 479
rect 1178 303 1238 736
rect 1288 303 1348 736
rect 1930 303 1990 736
rect 2044 460 2104 771
rect 2678 460 2738 771
rect 4387 736 4447 1123
rect 4552 947 4558 1007
rect 4618 947 4624 1007
rect 2792 303 2852 736
rect 3434 303 3494 736
rect 1172 243 1178 303
rect 1238 243 1288 303
rect 1348 243 1354 303
rect 1924 243 1930 303
rect 1990 243 1996 303
rect 2786 243 2792 303
rect 2852 243 2858 303
rect 3428 243 3434 303
rect 3494 243 3500 303
rect 3544 215 3604 736
rect 4186 215 4246 736
rect 4353 676 4447 736
rect 4558 460 4618 947
rect 3538 155 3544 215
rect 3604 155 3610 215
rect 4180 155 4186 215
rect 4246 155 4252 215
<< via1 >>
rect 912 1651 972 1711
rect 1554 1651 1614 1711
rect 2416 1651 2476 1711
rect 3058 1651 3118 1711
rect 3920 1651 3980 1711
rect 4562 1651 4622 1711
rect 1233 1387 1293 1447
rect 1664 1563 1724 1623
rect 2306 1563 2366 1623
rect 1985 1299 2045 1359
rect 2737 1387 2797 1447
rect 3168 1563 3228 1623
rect 3810 1563 3870 1623
rect 3489 1299 3549 1359
rect 4241 1387 4301 1447
rect 4387 1123 4447 1183
rect 2044 771 2104 831
rect 2678 771 2738 831
rect 916 419 976 479
rect 1609 419 1669 479
rect 2361 595 2421 655
rect 4558 947 4618 1007
rect 3113 419 3173 479
rect 1178 243 1238 303
rect 1288 243 1348 303
rect 1930 243 1990 303
rect 2792 243 2852 303
rect 3434 243 3494 303
rect 3865 507 3925 567
rect 3544 155 3604 215
rect 4186 155 4246 215
use cm_pcell2_cell  cm_pcell2_cell_0
timestamp 1749896124
transform -1 0 8137 0 1 -1741
box 3424 1732 8172 3616
<< end >>
