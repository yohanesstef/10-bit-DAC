magic
tech sky130A
magscale 1 2
timestamp 1749415301
<< error_s >>
rect 31807 -7208 31813 -7202
rect 31861 -7208 31867 -7202
rect 31801 -7214 31807 -7208
rect 31867 -7214 31873 -7208
rect 31801 -7268 31807 -7262
rect 31867 -7268 31873 -7262
rect 31807 -7274 31813 -7268
rect 31861 -7274 31867 -7268
rect 31531 -7296 31537 -7290
rect 31585 -7296 31591 -7290
rect 31525 -7302 31531 -7296
rect 31591 -7302 31597 -7296
rect 31525 -7356 31531 -7350
rect 31591 -7356 31597 -7350
rect 31531 -7362 31537 -7356
rect 31585 -7362 31591 -7356
rect 31255 -7384 31261 -7378
rect 31309 -7384 31315 -7378
rect 31249 -7390 31255 -7384
rect 31315 -7390 31321 -7384
rect 31249 -7444 31255 -7438
rect 31315 -7444 31321 -7438
rect 31255 -7450 31261 -7444
rect 31309 -7450 31315 -7444
rect 30979 -7472 30985 -7466
rect 31033 -7472 31039 -7466
rect 30973 -7478 30979 -7472
rect 31039 -7478 31045 -7472
rect 30973 -7532 30979 -7526
rect 31039 -7532 31045 -7526
rect 30979 -7538 30985 -7532
rect 31033 -7538 31039 -7532
rect 30495 -7560 30501 -7554
rect 30549 -7560 30555 -7554
rect 30489 -7566 30495 -7560
rect 30555 -7566 30561 -7560
rect 30489 -7620 30495 -7614
rect 30555 -7620 30561 -7614
rect 30495 -7626 30501 -7620
rect 30549 -7626 30555 -7620
rect 30219 -7648 30225 -7642
rect 30273 -7648 30279 -7642
rect 30213 -7654 30219 -7648
rect 30279 -7654 30285 -7648
rect 30213 -7708 30219 -7702
rect 30279 -7708 30285 -7702
rect 30219 -7714 30225 -7708
rect 30273 -7714 30279 -7708
rect 29943 -7736 29949 -7730
rect 29997 -7736 30003 -7730
rect 29937 -7742 29943 -7736
rect 30003 -7742 30009 -7736
rect 29937 -7796 29943 -7790
rect 30003 -7796 30009 -7790
rect 29943 -7802 29949 -7796
rect 29997 -7802 30003 -7796
rect 29667 -7824 29673 -7818
rect 29721 -7824 29727 -7818
rect 29661 -7830 29667 -7824
rect 29727 -7830 29733 -7824
rect 29661 -7884 29667 -7878
rect 29727 -7884 29733 -7878
rect 29667 -7890 29673 -7884
rect 29721 -7890 29727 -7884
<< metal1 >>
rect 31807 -7208 31867 -7202
rect 31531 -7296 31591 -7290
rect 31255 -7384 31315 -7378
rect 30979 -7472 31039 -7466
rect 30495 -7560 30555 -7554
rect 30219 -7648 30279 -7642
rect 29943 -7736 30003 -7730
rect 29667 -7824 29727 -7818
rect 29667 -8174 29727 -7884
rect 29943 -8174 30003 -7796
rect 30219 -8174 30279 -7708
rect 30495 -8174 30555 -7620
rect 29857 -8378 29903 -8174
rect 30133 -8290 30179 -8174
rect 30409 -8202 30455 -8174
rect 30409 -8262 30665 -8202
rect 30133 -8350 30577 -8290
rect 29857 -8438 30489 -8378
rect 30429 -8466 30489 -8438
rect 30517 -8466 30577 -8350
rect 30605 -8466 30665 -8262
rect 30693 -8466 30753 -8090
rect 30781 -8466 30841 -8090
rect 30979 -8174 31039 -7532
rect 31255 -8174 31315 -7444
rect 31358 -8170 31401 -8162
rect 31079 -8202 31125 -8174
rect 30869 -8262 31125 -8202
rect 30869 -8466 30929 -8262
rect 31355 -8290 31401 -8170
rect 31531 -8174 31591 -7356
rect 30957 -8350 31401 -8290
rect 30957 -8466 31017 -8350
rect 31631 -8378 31677 -8162
rect 31807 -8174 31867 -7268
rect 31045 -8438 31677 -8378
rect 31045 -8466 31105 -8438
<< via1 >>
rect 31807 -7268 31867 -7208
rect 31531 -7356 31591 -7296
rect 31255 -7444 31315 -7384
rect 30979 -7532 31039 -7472
rect 30495 -7620 30555 -7560
rect 30219 -7708 30279 -7648
rect 29943 -7796 30003 -7736
rect 29667 -7884 29727 -7824
use hpmos_8  hpmos_8_8
timestamp 1749415301
transform 1 0 29266 0 1 -8228
box 227 -172 2775 436
<< end >>
