magic
tech sky130A
magscale 1 2
timestamp 1749057406
<< pwell >>
rect -307 -1094 307 1094
<< psubdiff >>
rect -271 1024 -175 1058
rect 175 1024 271 1058
rect -271 962 -237 1024
rect 237 962 271 1024
rect -271 -1024 -237 -962
rect 237 -1024 271 -962
rect -271 -1058 -175 -1024
rect 175 -1058 271 -1024
<< psubdiffcont >>
rect -175 1024 175 1058
rect -271 -962 -237 962
rect 237 -962 271 962
rect -175 -1058 175 -1024
<< xpolycontact >>
rect -141 496 141 928
rect -141 -928 141 -496
<< xpolyres >>
rect -141 -496 141 496
<< locali >>
rect -271 1024 -175 1058
rect 175 1024 271 1058
rect -271 962 -237 1024
rect 237 962 271 1024
rect -271 -1024 -237 -962
rect 237 -1024 271 -962
rect -271 -1058 -175 -1024
rect 175 -1058 271 -1024
<< viali >>
rect -125 513 125 910
rect -125 -910 125 -513
<< metal1 >>
rect -131 910 131 922
rect -131 513 -125 910
rect 125 513 131 910
rect -131 501 131 513
rect -131 -513 131 -501
rect -131 -910 -125 -513
rect 125 -910 131 -513
rect -131 -922 131 -910
<< properties >>
string FIXED_BBOX -254 -1041 254 1041
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 5.115 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 7.522k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
