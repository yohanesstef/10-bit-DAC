* PEX produced on Wed Jun 11 16:28:55 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from lvsf.ext - technology: sky130A

.subckt lvsf_posim VPBIAS VNBIAS IN INB OUTP VDDH GND
X0 a_2725_n218.t1 OUTP.t2 a_3321_n121.t0 VDDH.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X1 VDDH.t1 VPBIAS.t0 a_2885_n121.t0 VDDH.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X2 a_2725_n218.t0 VNBIAS.t0 a_3191_n1615.t0 GND.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_3191_n1615.t1 IN.t0 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X4 a_2885_n121.t1 a_2725_n218.t2 OUTP.t0 VDDH.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X5 a_2925_n631.t0 VNBIAS.t1 OUTP.t1 GND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X6 a_3321_n121.t1 VPBIAS.t1 VDDH.t5 VDDH.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X7 GND.t5 INB.t0 a_2925_n631.t1 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
R0 OUTP.n0 OUTP.t0 227.856
R1 OUTP.n1 OUTP.t2 139.375
R2 OUTP.n0 OUTP.t1 83.3993
R3 OUTP.n1 OUTP.n0 6.09008
R4 OUTP OUTP.n1 0.0755
R5 a_3321_n121.t0 a_3321_n121.t1 55.3905
R6 a_2725_n218.n0 a_2725_n218.t1 228.04
R7 a_2725_n218.n0 a_2725_n218.t2 145.648
R8 a_2725_n218.t0 a_2725_n218.n0 83.2159
R9 VDDH.t4 VDDH.t3 378.611
R10 VDDH.t0 VDDH.t2 378.611
R11 VDDH.n2 VDDH.n0 200.111
R12 VDDH.n1 VDDH.t4 189.305
R13 VDDH.n1 VDDH.t0 189.305
R14 VDDH.n2 VDDH.n1 31.6793
R15 VDDH.n0 VDDH.t5 27.6955
R16 VDDH.n0 VDDH.t1 27.6955
R17 VDDH VDDH.n2 1.03175
R18 VPBIAS.n0 VPBIAS.t1 139.66
R19 VPBIAS.n0 VPBIAS.t0 139.206
R20 VPBIAS VPBIAS.n0 0.804667
R21 a_2885_n121.t0 a_2885_n121.t1 55.3905
R22 VNBIAS.n0 VNBIAS.t0 126.178
R23 VNBIAS.n0 VNBIAS.t1 124.9
R24 VNBIAS VNBIAS.n0 0.391454
R25 a_3191_n1615.t0 a_3191_n1615.t1 114.206
R26 GND.t2 GND.t1 749.482
R27 GND.t4 GND.t0 749.482
R28 GND.n1 GND.t2 125.389
R29 GND.n1 GND.t4 125.389
R30 GND.n2 GND.n1 90.7159
R31 GND.n2 GND.n0 25.0255
R32 GND.n0 GND.t3 5.8005
R33 GND.n0 GND.t5 5.8005
R34 GND GND.n2 1.03175
R35 IN IN.t0 713.933
R36 a_2925_n631.t0 a_2925_n631.t1 114.206
R37 INB INB.t0 713.749
C0 IN INB 0.07211f
C1 VDDH OUTP 0.24956f
C2 VNBIAS OUTP 0.10828f
C3 OUTP VPBIAS 0.17336f
C4 IN VNBIAS 0.0219f
C5 VNBIAS INB 0.01377f
C6 VDDH VNBIAS 0.01579f
C7 VDDH VPBIAS 0.89256f
C8 IN GND 0.22059f
C9 INB GND 0.21722f
C10 VNBIAS GND 1.25173f
C11 OUTP GND 0.54264f
C12 VPBIAS GND 0.54942f
C13 VDDH GND 2.28556f
.ends

