* PEX produced on Wed Jun 11 01:32:27 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from top_segment_1.ext - technology: sky130A

.subckt top_segment_1_posim V0 V64 DEC[0] DEC[1] DEC[2] DEC[3] b[0] b[1] b[2] b[3] bb[0]
+ bb[1] bb[2] bb[3] VOUT GND
X0 a_1875_4028.t4 DEC[0].t0 rseg_1_v3_1.v7.t2 GND.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1 GND.t45 GND.t46 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=2.5
X2 rseg_1_v3_1.v11.t2 rseg_1_v3_1.v10.t2 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=2.09
X3 rseg_1_v3_1.v34.t1 DEC[2].t0 a_337_4028.t2 GND.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X4 rseg_1_v3_1.v11.t1 DEC[0].t1 a_3049_5464.t4 GND.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X5 a_1323_4028.t3 DEC[2].t1 rseg_1_v3_1.v37.t2 GND.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X6 a_5799_6728.t2 bb[3].t0 a_n215_4028.t3 GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X7 rseg_1_v3_1.v10.t1 DEC[0].t2 a_2773_5464.t4 GND.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X8 a_3483_5464.t1 DEC[2].t2 rseg_1_v3_1.v44.t0 GND.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 rseg_1_v3_1.v61.t1 rseg_1_v3_1.v60.t1 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X10 rseg_1_v3_1.v13.t0 rseg_1_v3_1.v12.t0 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=1.89
X11 a_1599_4028.t1 DEC[3].t0 rseg_1_v3_1.v54.t0 GND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X12 a_7618_7809.t2 b[2].t0 a_7573_6728.t1 GND.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X13 GND.t54 GND.t55 GND.t47 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X14 rseg_1_v3_1.v39.t0 rseg_1_v3_1.v40.t0 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X15 rseg_1_v3_1.v3.t1 rseg_1_v3_1.v4.t0 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=3.37
X16 rseg_1_v3_1.v15.t0 rseg_1_v3_1.v16.t1 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=1.68
X17 a_4035_5464.t3 DEC[2].t3 rseg_1_v3_1.v46.t1 GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X18 a_8198_7809.t1 bb[1].t0 a_7010_7809.t2 GND.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X19 rseg_1_v3_1.v59.t1 DEC[3].t1 a_3049_5464.t0 GND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X20 GND.t97 GND.t98 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X21 GND.t85 GND.t86 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=2.35
X22 rseg_1_v3_1.v49.t0 rseg_1_v3_1.v50.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X23 a_7314_7809.t2 bb[0].t0 VOUT.t1 GND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X24 a_8198_7809.t0 bb[2].t0 a_6075_6728.t1 GND.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X25 a_1599_4028.t3 DEC[0].t3 rseg_1_v3_1.v6.t2 GND.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X26 rseg_1_v3_1.v7.t1 rseg_1_v3_1.v8.t1 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=2.5
X27 a_1875_4028.t1 DEC[2].t4 rseg_1_v3_1.v39.t1 GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X28 rseg_1_v3_1.v50.t1 DEC[3].t2 a_337_4028.t1 GND.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X29 rseg_1_v3_1.v9.t2 DEC[0].t4 a_2497_5464.t3 GND.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X30 a_3483_5464.t2 DEC[0].t5 rseg_1_v3_1.v12.t2 GND.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X31 a_6351_6728.t2 bb[3].t1 a_337_4028.t0 GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X32 V0.t1 DEC[0].t6 a_n215_4028.t2 GND.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X33 rseg_1_v3_1.v57.t2 rseg_1_v3_1.v58.t2 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X34 rseg_1_v3_1.v49.t1 DEC[3].t3 a_61_4028.t0 GND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X35 GND.t99 GND.t100 GND.t47 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X36 a_1047_4028.t0 DEC[3].t4 rseg_1_v3_1.v52.t2 GND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X37 rseg_1_v3_1.v47.t0 rseg_1_v3_1.v48.t1 GND.t47 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X38 a_7573_6728.t0 b[3].t0 a_4311_5464.t3 GND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X39 rseg_1_v3_1.v15.t1 rseg_1_v3_1.v14.t0 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X40 rseg_1_v3_1.v23.t0 rseg_1_v3_1.v24.t1 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X41 rseg_1_v3_1.v9.t1 rseg_1_v3_1.v8.t0 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=2.35
X42 rseg_1_v3_1.v59.t2 rseg_1_v3_1.v60.t0 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X43 a_8474_7809.t1 bb[2].t1 a_5799_6728.t0 GND.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X44 rseg_1_v3_1.v27.t1 rseg_1_v3_1.v28.t1 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X45 a_1323_4028.t4 DEC[0].t7 rseg_1_v3_1.v5.t2 GND.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X46 rseg_1_v3_1.v43.t0 DEC[2].t5 a_3049_5464.t2 GND.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X47 rseg_1_v3_1.v19.t0 DEC[1].t0 a_613_4028.t0 GND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X48 a_1599_4028.t2 DEC[2].t6 rseg_1_v3_1.v38.t1 GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X49 rseg_1_v3_1.v8.t2 DEC[0].t8 a_2221_5464.t4 GND.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X50 a_1599_4028.t0 DEC[1].t1 rseg_1_v3_1.v22.t0 GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X51 rseg_1_v3_1.v25.t2 rseg_1_v3_1.v26.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X52 rseg_1_v3_1.v21.t0 rseg_1_v3_1.v20.t0 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X53 rseg_1_v3_1.v51.t2 rseg_1_v3_1.v50.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X54 rseg_1_v3_1.v1.t0 rseg_1_v3_1.v2.t0 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=4.24
X55 rseg_1_v3_1.v48.t0 DEC[3].t5 a_n215_4028.t4 GND.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X56 rseg_1_v3_1.v51.t1 DEC[3].t6 a_613_4028.t1 GND.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X57 rseg_1_v3_1.v27.t2 DEC[1].t2 a_3049_5464.t3 GND.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X58 rseg_1_v3_1.v41.t2 rseg_1_v3_1.v40.t2 GND.t47 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X59 a_4035_5464.t1 DEC[1].t3 rseg_1_v3_1.v30.t0 GND.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X60 rseg_1_v3_1.v35.t0 rseg_1_v3_1.v36.t0 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X61 a_7297_6728.t0 b[3].t1 a_4035_5464.t2 GND.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X62 rseg_1_v3_1.v56.t0 DEC[3].t7 a_2221_5464.t1 GND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X63 a_7894_7809.t1 bb[2].t2 a_6351_6728.t1 GND.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X64 rseg_1_v3_1.v18.t1 DEC[1].t4 a_337_4028.t3 GND.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X65 rseg_1_v3_1.v51.t0 rseg_1_v3_1.v52.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X66 rseg_1_v3_1.v47.t2 rseg_1_v3_1.v46.t2 GND.t47 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X67 a_7618_7809.t0 b[1].t0 a_7010_7809.t0 GND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X68 rseg_1_v3_1.v42.t0 DEC[2].t7 a_2773_5464.t3 GND.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X69 a_1047_4028.t3 DEC[0].t9 rseg_1_v3_1.v4.t2 GND.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X70 a_1323_4028.t0 DEC[1].t5 rseg_1_v3_1.v21.t1 GND.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X71 GND.t128 GND.t129 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X72 rseg_1_v3_1.v33.t1 DEC[2].t8 a_61_4028.t2 GND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X73 a_1047_4028.t1 DEC[2].t9 rseg_1_v3_1.v36.t2 GND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X74 rseg_1_v3_1.v55.t1 rseg_1_v3_1.v54.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X75 rseg_1_v3_1.v26.t1 DEC[1].t6 a_2773_5464.t2 GND.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X76 rseg_1_v3_1.v59.t0 rseg_1_v3_1.v58.t0 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X77 rseg_1_v3_1.v27.t0 rseg_1_v3_1.v26.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X78 a_3759_5464.t0 DEC[1].t7 rseg_1_v3_1.v29.t0 GND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X79 a_7894_7809.t2 b[2].t1 a_7297_6728.t1 GND.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X80 a_7021_6728.t0 b[3].t2 a_3759_5464.t3 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X81 a_2497_5464.t0 b[3].t3 a_6075_6728.t0 GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X82 a_3483_5464.t0 DEC[1].t8 rseg_1_v3_1.v28.t0 GND.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X83 a_6745_6728.t0 b[3].t4 a_3483_5464.t3 GND.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X84 rseg_1_v3_1.v21.t2 rseg_1_v3_1.v22.t1 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X85 rseg_1_v3_1.v37.t1 rseg_1_v3_1.v36.t1 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X86 rseg_1_v3_1.v41.t0 DEC[2].t10 a_2497_5464.t2 GND.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X87 a_1047_4028.t2 DEC[1].t9 rseg_1_v3_1.v20.t1 GND.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X88 GND.t71 GND.t72 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X89 rseg_1_v3_1.v32.t2 DEC[2].t11 a_n215_4028.t1 GND.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X90 a_8474_7809.t2 b[2].t2 a_6745_6728.t1 GND.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X91 rseg_1_v3_1.v16.t0 DEC[1].t10 a_n215_4028.t0 GND.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X92 rseg_1_v3_1.v31.t2 rseg_1_v3_1.v30.t1 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X93 rseg_1_v3_1.v49.t2 rseg_1_v3_1.v48.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X94 rseg_1_v3_1.v35.t2 DEC[2].t12 a_613_4028.t2 GND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X95 a_7894_7809.t0 b[1].t1 a_7314_7809.t0 GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X96 a_4035_5464.t0 DEC[3].t8 rseg_1_v3_1.v62.t1 GND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X97 rseg_1_v3_1.v53.t0 rseg_1_v3_1.v52.t1 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X98 a_7010_7809.t1 b[0].t0 VOUT.t0 GND.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X99 rseg_1_v3_1.v11.t0 rseg_1_v3_1.v12.t1 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=1.99
X100 a_8198_7809.t2 b[2].t3 a_7021_6728.t1 GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X101 rseg_1_v3_1.v45.t0 rseg_1_v3_1.v46.t0 GND.t47 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X102 rseg_1_v3_1.v24.t0 DEC[1].t11 a_2221_5464.t0 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X103 a_2221_5464.t3 b[3].t5 a_5799_6728.t1 GND.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X104 a_3049_5464.t1 b[3].t6 a_6627_6728.t1 GND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X105 GND.t39 GND.t40 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X106 GND.t37 GND.t38 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X107 rseg_1_v3_1.v19.t2 rseg_1_v3_1.v18.t2 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X108 GND.t74 GND.t75 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X109 rseg_1_v3_1.v40.t1 DEC[2].t13 a_2221_5464.t2 GND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X110 GND.t95 GND.t96 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X111 rseg_1_v3_1.v33.t2 rseg_1_v3_1.v34.t2 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X112 rseg_1_v3_1.v45.t2 rseg_1_v3_1.v44.t1 GND.t47 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X113 rseg_1_v3_1.v9.t0 rseg_1_v3_1.v10.t0 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=2.19
X114 rseg_1_v3_1.v31.t1 rseg_1_v3_1.v32.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X115 rseg_1_v3_1.v5.t1 rseg_1_v3_1.v4.t1 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=3.12
X116 rseg_1_v3_1.v19.t1 rseg_1_v3_1.v20.t2 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X117 rseg_1_v3_1.v37.t0 rseg_1_v3_1.v38.t0 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X118 GND.t2 GND.t3 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X119 a_2773_5464.t0 b[3].t7 a_6351_6728.t0 GND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X120 rseg_1_v3_1.v5.t0 rseg_1_v3_1.v6.t1 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=2.86
X121 rseg_1_v3_1.v25.t1 rseg_1_v3_1.v24.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X122 rseg_1_v3_1.v17.t0 rseg_1_v3_1.v18.t0 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X123 a_1047_4028.t4 bb[3].t2 a_6745_6728.t2 GND.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X124 a_4035_5464.t4 DEC[0].t10 rseg_1_v3_1.v14.t1 GND.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X125 rseg_1_v3_1.v1.t1 V0.t0 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X126 a_1875_4028.t2 bb[3].t3 a_7573_6728.t2 GND.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X127 rseg_1_v3_1.v1.t2 DEC[0].t11 a_61_4028.t3 GND.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X128 GND.t87 GND.t88 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X129 rseg_1_v3_1.v53.t2 rseg_1_v3_1.v54.t1 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X130 rseg_1_v3_1.v29.t1 rseg_1_v3_1.v30.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X131 rseg_1_v3_1.v3.t0 rseg_1_v3_1.v2.t1 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=3.73
X132 a_4311_5464.t2 DEC[2].t14 rseg_1_v3_1.v47.t1 GND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X133 rseg_1_v3_1.v57.t1 rseg_1_v3_1.v56.t1 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X134 rseg_1_v3_1.v33.t0 rseg_1_v3_1.v32.t1 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X135 rseg_1_v3_1.v17.t1 DEC[1].t12 a_61_4028.t1 GND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X136 rseg_1_v3_1.v3.t2 DEC[0].t12 a_613_4028.t3 GND.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X137 a_4311_5464.t1 DEC[3].t9 rseg_1_v3_1.v63.t0 GND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X138 rseg_1_v3_1.v39.t2 rseg_1_v3_1.v38.t2 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X139 GND.t93 GND.t94 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X140 rseg_1_v3_1.v25.t0 DEC[1].t13 a_2497_5464.t4 GND.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X141 rseg_1_v3_1.v41.t1 rseg_1_v3_1.v42.t1 GND.t47 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X142 rseg_1_v3_1.v29.t2 rseg_1_v3_1.v28.t2 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X143 rseg_1_v3_1.v35.t1 rseg_1_v3_1.v34.t0 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X144 rseg_1_v3_1.v63.t2 rseg_1_v3_1.v62.t2 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X145 a_3759_5464.t4 DEC[0].t13 rseg_1_v3_1.v13.t1 GND.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X146 a_6627_6728.t2 bb[3].t4 a_613_4028.t4 GND.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X147 rseg_1_v3_1.v23.t2 rseg_1_v3_1.v22.t2 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X148 rseg_1_v3_1.v17.t2 rseg_1_v3_1.v16.t2 GND.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X149 a_1599_4028.t4 bb[3].t5 a_7297_6728.t2 GND.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X150 rseg_1_v3_1.v43.t2 rseg_1_v3_1.v44.t2 GND.t47 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X151 rseg_1_v3_1.v55.t2 rseg_1_v3_1.v56.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X152 a_1323_4028.t2 DEC[3].t10 rseg_1_v3_1.v53.t1 GND.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X153 rseg_1_v3_1.v2.t2 DEC[0].t14 a_337_4028.t4 GND.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X154 rseg_1_v3_1.v58.t1 DEC[3].t11 a_2773_5464.t1 GND.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X155 a_3759_5464.t1 DEC[3].t12 rseg_1_v3_1.v61.t2 GND.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X156 rseg_1_v3_1.v63.t1 V64.t0 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X157 a_1875_4028.t3 DEC[1].t14 rseg_1_v3_1.v23.t1 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X158 a_1323_4028.t1 bb[3].t6 a_7021_6728.t2 GND.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X159 a_4311_5464.t4 DEC[0].t15 rseg_1_v3_1.v15.t2 GND.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X160 a_6075_6728.t2 bb[3].t7 a_61_4028.t4 GND.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X161 a_3759_5464.t2 DEC[2].t15 rseg_1_v3_1.v45.t1 GND.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X162 rseg_1_v3_1.v7.t0 rseg_1_v3_1.v6.t0 GND.t6 sky130_fd_pr__res_xhigh_po_1p41 l=2.66
X163 GND.t67 GND.t68 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=1.68
X164 a_1875_4028.t0 DEC[3].t13 rseg_1_v3_1.v55.t0 GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X165 a_4311_5464.t0 DEC[1].t15 rseg_1_v3_1.v31.t0 GND.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X166 GND.t65 GND.t66 GND.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X167 rseg_1_v3_1.v13.t2 rseg_1_v3_1.v14.t2 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=1.84
X168 rseg_1_v3_1.v57.t0 DEC[3].t14 a_2497_5464.t1 GND.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X169 rseg_1_v3_1.v43.t1 rseg_1_v3_1.v42.t2 GND.t47 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X170 rseg_1_v3_1.v61.t0 rseg_1_v3_1.v62.t0 GND.t20 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X171 a_8474_7809.t0 bb[1].t1 a_7314_7809.t1 GND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X172 a_3483_5464.t4 DEC[3].t15 rseg_1_v3_1.v60.t2 GND.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X173 a_7618_7809.t1 bb[2].t3 a_6627_6728.t0 GND.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
R0 DEC[0].n10 DEC[0].t6 213.218
R1 DEC[0].n7 DEC[0].t0 213.218
R2 DEC[0].n0 DEC[0].t15 213.218
R3 DEC[0].n10 DEC[0].t11 212.554
R4 DEC[0].n11 DEC[0].t14 212.554
R5 DEC[0].n12 DEC[0].t12 212.554
R6 DEC[0].n9 DEC[0].t9 212.554
R7 DEC[0].n8 DEC[0].t7 212.554
R8 DEC[0].n7 DEC[0].t3 212.554
R9 DEC[0].n6 DEC[0].t8 212.554
R10 DEC[0].n5 DEC[0].t4 212.554
R11 DEC[0].n4 DEC[0].t2 212.554
R12 DEC[0].n3 DEC[0].t1 212.554
R13 DEC[0].n2 DEC[0].t5 212.554
R14 DEC[0].n1 DEC[0].t13 212.554
R15 DEC[0].n0 DEC[0].t10 212.554
R16 DEC[0] DEC[0].n13 14.3922
R17 DEC[0].n12 DEC[0].n11 0.663962
R18 DEC[0].n11 DEC[0].n10 0.663962
R19 DEC[0].n8 DEC[0].n7 0.663962
R20 DEC[0].n9 DEC[0].n8 0.663962
R21 DEC[0].n1 DEC[0].n0 0.663962
R22 DEC[0].n2 DEC[0].n1 0.663962
R23 DEC[0].n3 DEC[0].n2 0.663962
R24 DEC[0].n4 DEC[0].n3 0.663962
R25 DEC[0].n5 DEC[0].n4 0.663962
R26 DEC[0].n6 DEC[0].n5 0.663962
R27 DEC[0].n13 DEC[0].n12 0.312199
R28 DEC[0].n13 DEC[0].n9 0.312199
R29 DEC[0] DEC[0].n6 0.254667
R30 rseg_1_v3_1.v7 rseg_1_v3_1.v7.t2 248.075
R31 rseg_1_v3_1.v7.n0 rseg_1_v3_1.v7.t1 10.5773
R32 rseg_1_v3_1.v7.n0 rseg_1_v3_1.v7.t0 10.5739
R33 rseg_1_v3_1.v7 rseg_1_v3_1.v7.n0 4.31612
R34 a_1875_4028.n0 a_1875_4028.t4 248.653
R35 a_1875_4028.t0 a_1875_4028.n2 246.668
R36 a_1875_4028.n1 a_1875_4028.t2 243.488
R37 a_1875_4028.n0 a_1875_4028.t3 240
R38 a_1875_4028.n2 a_1875_4028.t1 240
R39 a_1875_4028.n1 a_1875_4028.n0 5.15258
R40 a_1875_4028.n2 a_1875_4028.n1 1.86925
R41 GND.n117 GND.n71 28676.6
R42 GND.n156 GND.n117 28676.6
R43 GND.n160 GND.n71 28673.3
R44 GND.n160 GND.n156 28673.3
R45 GND.n102 GND.n97 7416.07
R46 GND.n102 GND.n98 7416.07
R47 GND.n98 GND.n92 7416.07
R48 GND.n97 GND.n92 7416.07
R49 GND.n206 GND.n4 4458.86
R50 GND.n206 GND.n5 4458.86
R51 GND.n208 GND.n5 4458.86
R52 GND.n208 GND.n4 4458.86
R53 GND.n176 GND.n35 4458.86
R54 GND.n178 GND.n35 4458.86
R55 GND.n178 GND.n34 4458.86
R56 GND.n176 GND.n34 4458.86
R57 GND.n58 GND.n26 4458.86
R58 GND.n58 GND.n27 4458.86
R59 GND.n185 GND.n27 4458.86
R60 GND.n185 GND.n26 4458.86
R61 GND.n107 GND.n88 4458.86
R62 GND.n90 GND.n88 4458.86
R63 GND.n90 GND.n86 4458.86
R64 GND.n107 GND.n86 4458.86
R65 GND.n114 GND.n77 4458.86
R66 GND.n77 GND.n72 4458.86
R67 GND.n73 GND.n72 4458.86
R68 GND.n114 GND.n73 4458.86
R69 GND.n158 GND.n36 4458.86
R70 GND.n158 GND.n37 4458.86
R71 GND.n167 GND.n37 4458.86
R72 GND.n167 GND.n36 4458.86
R73 GND.n64 GND.n43 4458.86
R74 GND.n64 GND.n44 4458.86
R75 GND.n56 GND.n44 4458.86
R76 GND.n56 GND.n43 4458.86
R77 GND.n188 GND.n24 4458.86
R78 GND.n25 GND.n24 4458.86
R79 GND.n25 GND.n23 4458.86
R80 GND.n188 GND.n23 4458.86
R81 GND.n195 GND.n16 4458.86
R82 GND.n16 GND.n14 4458.86
R83 GND.n15 GND.n14 4458.86
R84 GND.n195 GND.n15 4458.86
R85 GND.n198 GND.n11 4458.86
R86 GND.n198 GND.n12 4458.86
R87 GND.n13 GND.n12 4458.86
R88 GND.n13 GND.n11 4458.86
R89 GND.n202 GND.n201 982.966
R90 GND.n101 GND.n99 852.33
R91 GND.n101 GND.n100 852.33
R92 GND.n91 GND.n9 781.929
R93 GND.n91 GND.n7 781.929
R94 GND.n165 GND.n66 669.365
R95 GND.n41 GND.n40 646.4
R96 GND GND.n0 583.907
R97 GND.n175 GND.n174 514.26
R98 GND.n113 GND.n78 514.26
R99 GND.n81 GND.n78 514.26
R100 GND.n68 GND.n67 514.26
R101 GND.n49 GND.n48 514.26
R102 GND.n199 GND.n10 514.26
R103 GND.n205 GND.n204 514.26
R104 GND.n161 GND.n70 511.591
R105 GND.n135 GND.n134 461.243
R106 GND.n136 GND.n135 459.111
R107 GND.n108 GND.n85 443.86
R108 GND.n171 GND.n170 443.86
R109 GND.n175 GND.n173 443.86
R110 GND.n82 GND.n81 443.86
R111 GND.n89 GND.n18 443.86
R112 GND.n89 GND.n21 443.86
R113 GND.n183 GND.n182 443.86
R114 GND.n182 GND.n181 443.86
R115 GND.n180 GND.n179 443.86
R116 GND.n179 GND.n33 443.86
R117 GND.n165 GND.n164 443.86
R118 GND.n50 GND.n49 443.86
R119 GND.n52 GND.n51 443.86
R120 GND.n53 GND.n52 443.86
R121 GND.n54 GND.n39 443.86
R122 GND.n67 GND.n38 443.86
R123 GND.n80 GND.n79 443.86
R124 GND.n79 GND.n0 443.86
R125 GND.n210 GND.n209 443.86
R126 GND.n209 GND.n3 443.86
R127 GND.n203 GND.n202 431.812
R128 GND.n181 GND.n180 428.8
R129 GND.n66 GND.n39 427.671
R130 GND.n170 GND.n2 414.872
R131 GND.n173 GND.n172 399.812
R132 GND GND.n210 399.06
R133 GND.n54 GND.n53 380.988
R134 GND.n46 GND.n45 380.988
R135 GND.n162 GND.n161 361.601
R136 GND.n82 GND.n17 350.872
R137 GND.n193 GND.n18 350.872
R138 GND.n190 GND.n21 350.872
R139 GND.n183 GND.n22 350.872
R140 GND.n181 GND.n29 350.872
R141 GND.n180 GND.n32 350.872
R142 GND.n40 GND.n33 350.872
R143 GND.n48 GND.n17 345.976
R144 GND.n85 GND.n28 338.825
R145 GND.n183 GND.n21 338.825
R146 GND.n112 GND.n80 332.8
R147 GND.n109 GND.n0 332.8
R148 GND.n210 GND.n2 332.8
R149 GND.n172 GND.n3 332.8
R150 GND.n51 GND.n50 317.365
R151 GND.n192 GND.n191 317.365
R152 GND.n112 GND.n111 313.601
R153 GND.n193 GND.n192 310.589
R154 GND.n111 GND.n110 301.553
R155 GND.n82 GND.n18 301.553
R156 GND.n164 GND.n163 295.906
R157 GND.n200 GND.n199 294.776
R158 GND.n46 GND.n22 289.13
R159 GND.n110 GND.n109 272.565
R160 GND.n191 GND.n190 259.765
R161 GND.n73 GND.t34 257.123
R162 GND.t114 GND.n158 257.123
R163 GND.n41 GND.n32 241.319
R164 GND.n200 GND.n9 240.565
R165 GND.n203 GND.n7 240.565
R166 GND.n118 GND.n69 235.98
R167 GND.n42 GND.n29 226.26
R168 GND.n45 GND.n29 217.601
R169 GND.n146 GND.n145 207.393
R170 GND.n42 GND.n32 202.542
R171 GND.n163 GND.n68 195.766
R172 GND.n190 GND.n189 184.095
R173 GND.n150 GND.n149 172.619
R174 GND.n142 GND.n141 171.554
R175 GND.n119 GND.n118 171.339
R176 GND.n129 GND.n128 171.339
R177 GND.n133 GND.n132 171.339
R178 GND.n138 GND.n137 171.339
R179 GND.n109 GND.n108 171.294
R180 GND.n124 GND.n123 170.274
R181 GND.n194 GND.n17 168.282
R182 GND.n189 GND.n22 154.73
R183 GND.n144 GND.n143 151.714
R184 GND.n127 GND.n126 151.5
R185 GND.n131 GND.n130 151.5
R186 GND.n140 GND.n139 150.434
R187 GND.n122 GND.n121 149.367
R188 GND.n201 GND.n200 149.083
R189 GND.n48 GND.n15 146.25
R190 GND.n75 GND.n15 146.25
R191 GND.n19 GND.n16 146.25
R192 GND.n94 GND.n16 146.25
R193 GND.n23 GND.n20 146.25
R194 GND.n105 GND.n23 146.25
R195 GND.n47 GND.n24 146.25
R196 GND.n153 GND.n24 146.25
R197 GND.n56 GND.n55 146.25
R198 GND.n57 GND.n56 146.25
R199 GND.n65 GND.n64 146.25
R200 GND.n64 GND.n63 146.25
R201 GND.n167 GND.n166 146.25
R202 GND.n168 GND.n167 146.25
R203 GND.n158 GND.n68 146.25
R204 GND.n78 GND.n73 146.25
R205 GND.n83 GND.n77 146.25
R206 GND.n77 GND.n76 146.25
R207 GND.n86 GND.n84 146.25
R208 GND.n93 GND.n86 146.25
R209 GND.n88 GND.n87 146.25
R210 GND.n104 GND.n88 146.25
R211 GND.n185 GND.n184 146.25
R212 GND.n186 GND.n185 146.25
R213 GND.n58 GND.n30 146.25
R214 GND.n59 GND.n58 146.25
R215 GND.n34 GND.n31 146.25
R216 GND.n62 GND.n34 146.25
R217 GND.n174 GND.n35 146.25
R218 GND.n169 GND.n35 146.25
R219 GND.n4 GND.n1 146.25
R220 GND.n152 GND.n4 146.25
R221 GND.n99 GND.n97 146.25
R222 GND.n97 GND.n96 146.25
R223 GND.n100 GND.n98 146.25
R224 GND.n98 GND.n6 146.25
R225 GND.n12 GND.n8 146.25
R226 GND.n95 GND.n12 146.25
R227 GND.n11 GND.n10 146.25
R228 GND.n74 GND.n11 146.25
R229 GND.n204 GND.n5 146.25
R230 GND.n60 GND.n5 146.25
R231 GND.t90 GND.t89 143.666
R232 GND.t89 GND.t131 143.666
R233 GND.t103 GND.t35 143.666
R234 GND.t119 GND.t118 143.666
R235 GND.t118 GND.t116 143.666
R236 GND.t116 GND.t112 143.666
R237 GND.t117 GND.t120 143.666
R238 GND.t111 GND.t113 143.666
R239 GND.t106 GND.t108 143.666
R240 GND.t109 GND.t106 143.666
R241 GND.n148 GND.n147 142.754
R242 GND.t1 GND.t19 141.583
R243 GND.n145 GND.n70 135.286
R244 GND.t107 GND.t53 133.775
R245 GND.n194 GND.n193 133.272
R246 GND.n113 GND.n112 130.26
R247 GND.n147 GND.n146 128.887
R248 GND.t29 GND.t130 116.599
R249 GND.n116 GND.t90 115.037
R250 GND.t6 GND.t117 114.516
R251 GND.n94 GND.t77 112.433
R252 GND.t10 GND.t105 111.913
R253 GND.t112 GND.n169 110.873
R254 GND.n168 GND.t120 110.873
R255 GND.n74 GND.t8 108.269
R256 GND.t16 GND.t50 108.269
R257 GND.t79 GND.t82 103.585
R258 GND.t57 GND.t123 102.023
R259 GND.t125 GND.t49 102.023
R260 GND.n120 GND.n119 100.299
R261 GND.n162 GND.n69 99.6436
R262 GND.n123 GND.n122 96.0333
R263 GND.t126 GND.n186 92.1335
R264 GND.t69 GND.t127 91.0924
R265 GND.t14 GND.t91 91.0924
R266 GND.n149 GND.n148 84.94
R267 GND.n163 GND.n162 80.0005
R268 GND.n121 GND.n66 80.0005
R269 GND.t23 GND.t48 79.6409
R270 GND.t92 GND.t62 79.6409
R271 GND.t28 GND.t73 79.1203
R272 GND.t44 GND.n62 79.1203
R273 GND.n63 GND.t110 79.1203
R274 GND.n159 GND.t114 78.0793
R275 GND.t80 GND.t26 75.4767
R276 GND.t36 GND.t70 75.4767
R277 GND.n66 GND.n65 74.0272
R278 GND.t17 GND.t124 73.3946
R279 GND.n128 GND.n127 72.14
R280 GND.n115 GND.t8 71.833
R281 GND.n106 GND.t81 71.833
R282 GND.n187 GND.t84 71.833
R283 GND.n61 GND.t101 71.833
R284 GND.t35 GND.n61 71.833
R285 GND.n177 GND.t115 71.833
R286 GND.n177 GND.t119 71.833
R287 GND.n157 GND.t111 71.833
R288 GND.t108 GND.n157 71.833
R289 GND.n151 GND.n150 70.499
R290 GND.n100 GND.n7 70.4005
R291 GND.n99 GND.n9 70.4005
R292 GND.n202 GND.n1 70.4005
R293 GND.n210 GND.n1 70.4005
R294 GND.n174 GND.n33 70.4005
R295 GND.n171 GND.n30 70.4005
R296 GND.n181 GND.n30 70.4005
R297 GND.n184 GND.n28 70.4005
R298 GND.n184 GND.n183 70.4005
R299 GND.n87 GND.n85 70.4005
R300 GND.n87 GND.n21 70.4005
R301 GND.n110 GND.n84 70.4005
R302 GND.n84 GND.n18 70.4005
R303 GND.n111 GND.n83 70.4005
R304 GND.n83 GND.n82 70.4005
R305 GND.n173 GND.n31 70.4005
R306 GND.n180 GND.n31 70.4005
R307 GND.n166 GND.n38 70.4005
R308 GND.n166 GND.n165 70.4005
R309 GND.n192 GND.n19 70.4005
R310 GND.n50 GND.n19 70.4005
R311 GND.n191 GND.n20 70.4005
R312 GND.n51 GND.n20 70.4005
R313 GND.n47 GND.n46 70.4005
R314 GND.n53 GND.n47 70.4005
R315 GND.n55 GND.n45 70.4005
R316 GND.n55 GND.n54 70.4005
R317 GND.n65 GND.n41 70.4005
R318 GND.n201 GND.n8 70.4005
R319 GND.n8 GND.n0 70.4005
R320 GND.n80 GND.n10 70.4005
R321 GND.n204 GND.n3 70.4005
R322 GND.t13 GND.n104 69.2304
R323 GND.n141 GND.n140 67.4467
R324 GND.n159 GND.t109 65.5867
R325 GND.n125 GND.n124 65.3297
R326 GND.n143 GND.n142 65.3133
R327 GND.n62 GND.t103 64.5456
R328 GND.n63 GND.t107 64.5456
R329 GND.n132 GND.n131 63.18
R330 GND.n155 GND.t33 62.9841
R331 GND.n130 GND.n129 61.0467
R332 GND.n137 GND.n136 58.9133
R333 GND.n139 GND.n138 58.9133
R334 GND.t12 GND.t42 58.8199
R335 GND.t9 GND.n75 58.2993
R336 GND.t132 GND.n95 58.2993
R337 GND.n57 GND.t25 57.2583
R338 GND.t19 GND.n60 57.2583
R339 GND.n134 GND.n133 54.6467
R340 GND.t30 GND.t9 52.5736
R341 GND.t63 GND.t80 52.5736
R342 GND.t127 GND.t27 52.5736
R343 GND.t91 GND.t52 52.5736
R344 GND.t84 GND.t126 49.9709
R345 GND.n96 GND.t22 48.4093
R346 GND.t133 GND.n57 46.3272
R347 GND.n59 GND.t32 46.3272
R348 GND.t131 GND.t20 45.8067
R349 GND.t18 GND.t7 44.7657
R350 GND.t76 GND.t12 44.7657
R351 GND.n169 GND.n168 40.6015
R352 GND.t82 GND.t104 40.0809
R353 GND.t25 GND.t79 40.0809
R354 GND.t51 GND.t133 40.0809
R355 GND.t83 GND.t28 40.0809
R356 GND.n60 GND.n59 40.0809
R357 GND.n119 GND.t68 39.3159
R358 GND.n118 GND.t39 39.3159
R359 GND.n69 GND.t40 39.3159
R360 GND.n120 GND.t67 39.3159
R361 GND.n122 GND.t3 39.3159
R362 GND.n123 GND.t2 39.3159
R363 GND.n124 GND.t72 39.3159
R364 GND.n126 GND.t71 39.3159
R365 GND.n127 GND.t75 39.3159
R366 GND.n128 GND.t74 39.3159
R367 GND.n129 GND.t55 39.3159
R368 GND.n130 GND.t54 39.3159
R369 GND.n131 GND.t129 39.3159
R370 GND.n132 GND.t128 39.3159
R371 GND.n133 GND.t94 39.3159
R372 GND.n134 GND.t93 39.3159
R373 GND.n136 GND.t95 39.3159
R374 GND.n137 GND.t96 39.3159
R375 GND.n138 GND.t87 39.3159
R376 GND.n139 GND.t88 39.3159
R377 GND.n140 GND.t99 39.3159
R378 GND.n141 GND.t100 39.3159
R379 GND.n142 GND.t65 39.3159
R380 GND.n143 GND.t66 39.3159
R381 GND.n144 GND.t37 39.3159
R382 GND.n150 GND.t38 39.3159
R383 GND.n149 GND.t97 39.3159
R384 GND.n148 GND.t98 39.3159
R385 GND.n147 GND.t85 39.3159
R386 GND.n146 GND.t86 39.3159
R387 GND.n145 GND.t45 39.3159
R388 GND.n70 GND.t46 39.3159
R389 GND.t130 GND.n105 39.0399
R390 GND.n152 GND.t122 38.5194
R391 GND.t56 GND.n153 38.5194
R392 GND.t64 GND.t132 36.9578
R393 GND.t31 GND.n74 35.3962
R394 GND.n76 GND.t36 35.3962
R395 GND.t41 GND.t125 35.3962
R396 GND.t24 GND.t13 35.3962
R397 GND.t15 GND.t16 35.3962
R398 GND.t61 GND.t18 34.3552
R399 GND.t121 GND.t76 34.3552
R400 GND.t4 GND.n196 33.8346
R401 GND.n106 GND.t47 33.8346
R402 GND.t78 GND.n154 31.7525
R403 GND.n207 GND.t104 31.7525
R404 GND.t105 GND.t44 31.7525
R405 GND.t110 GND.t10 31.7525
R406 GND.t48 GND.n93 31.232
R407 GND.t58 GND.t17 30.191
R408 GND.n40 GND.n38 29.3652
R409 GND.t113 GND.t6 29.1499
R410 GND.n28 GND.n2 28.9887
R411 GND.n172 GND.n171 28.9887
R412 GND.n116 GND.t34 28.6294
R413 GND.t60 GND.t11 27.0678
R414 GND.t77 GND.t43 27.0678
R415 GND.t81 GND.t29 27.0678
R416 GND.t50 GND.t5 27.0678
R417 GND.t20 GND.n115 26.0268
R418 GND.t7 GND.n152 26.0268
R419 GND.n155 GND.t56 24.9857
R420 GND.n104 GND.n103 24.4652
R421 GND.t59 GND.t0 24.4652
R422 GND.t73 GND.t51 24.4652
R423 GND.t32 GND.t83 24.4652
R424 GND.n154 GND.n6 23.4241
R425 GND.t5 GND.t21 22.9036
R426 GND.n187 GND.t21 21.8626
R427 GND.n93 GND.t14 21.342
R428 GND.n95 GND.t60 21.342
R429 GND.n197 GND.t27 19.2599
R430 GND.n196 GND.t52 19.2599
R431 GND.n197 GND.t4 18.7394
R432 GND.n195 GND.n194 18.2817
R433 GND.n196 GND.n195 18.2817
R434 GND.n49 GND.n14 18.2817
R435 GND.n196 GND.n14 18.2817
R436 GND.n189 GND.n188 18.2817
R437 GND.n188 GND.n187 18.2817
R438 GND.n52 GND.n25 18.2817
R439 GND.n187 GND.n25 18.2817
R440 GND.n43 GND.n42 18.2817
R441 GND.n61 GND.n43 18.2817
R442 GND.n44 GND.n39 18.2817
R443 GND.n61 GND.n44 18.2817
R444 GND.n67 GND.n36 18.2817
R445 GND.n157 GND.n36 18.2817
R446 GND.n164 GND.n37 18.2817
R447 GND.n157 GND.n37 18.2817
R448 GND.n114 GND.n113 18.2817
R449 GND.n115 GND.n114 18.2817
R450 GND.n81 GND.n72 18.2817
R451 GND.n115 GND.n72 18.2817
R452 GND.n108 GND.n107 18.2817
R453 GND.n107 GND.n106 18.2817
R454 GND.n90 GND.n89 18.2817
R455 GND.n106 GND.n90 18.2817
R456 GND.n170 GND.n26 18.2817
R457 GND.n154 GND.n26 18.2817
R458 GND.n182 GND.n27 18.2817
R459 GND.n154 GND.n27 18.2817
R460 GND.n176 GND.n175 18.2817
R461 GND.n177 GND.n176 18.2817
R462 GND.n179 GND.n178 18.2817
R463 GND.n178 GND.n177 18.2817
R464 GND.n199 GND.n198 18.2817
R465 GND.n198 GND.n197 18.2817
R466 GND.n206 GND.n205 18.2817
R467 GND.n207 GND.n206 18.2817
R468 GND.n79 GND.n13 18.2817
R469 GND.n197 GND.n13 18.2817
R470 GND.n209 GND.n208 18.2817
R471 GND.n208 GND.n207 18.2817
R472 GND.n75 GND.t31 17.1778
R473 GND.n76 GND.t69 17.1778
R474 GND.n207 GND.n6 16.6573
R475 GND.t26 GND.t30 15.6163
R476 GND.t70 GND.t63 15.6163
R477 GND.t102 GND.t64 15.6163
R478 GND.t33 GND.t59 15.6163
R479 GND.t0 GND.t78 15.6163
R480 GND.n103 GND.t15 14.5752
R481 GND.n161 GND.n160 13.296
R482 GND.n160 GND.n159 13.296
R483 GND.n135 GND.n117 13.296
R484 GND.n117 GND.n116 13.296
R485 GND.n205 GND.n203 12.0476
R486 GND.t22 GND.t23 11.4521
R487 GND.t62 GND.t102 11.4521
R488 GND.t43 GND.t47 10.9315
R489 GND.n151 GND.n144 10.1749
R490 GND.n92 GND.n91 9.91575
R491 GND.n103 GND.n92 9.91575
R492 GND.n102 GND.n101 9.91575
R493 GND.n103 GND.n102 9.91575
R494 GND.t53 GND.t115 9.89048
R495 GND.n126 GND.n125 8.94409
R496 GND.t123 GND.t41 6.2468
R497 GND.t49 GND.t24 6.2468
R498 GND.t42 GND.t61 5.72628
R499 GND.t124 GND.t121 5.72628
R500 GND.n96 GND.t92 4.1647
R501 GND.t11 GND.n94 4.1647
R502 GND.n156 GND.n151 2.9255
R503 GND.n156 GND.n155 2.9255
R504 GND.n125 GND.n71 2.9255
R505 GND.n155 GND.n71 2.9255
R506 GND.n105 GND.t57 2.60313
R507 GND.n121 GND.n120 2.13383
R508 GND.t101 GND.t1 2.0826
R509 GND.n186 GND.t122 1.56208
R510 GND.n153 GND.t58 1.56208
R511 rseg_1_v3_1.v11 rseg_1_v3_1.v11.t1 248.95
R512 rseg_1_v3_1.v11.n0 rseg_1_v3_1.v11.t0 10.5761
R513 rseg_1_v3_1.v11.n0 rseg_1_v3_1.v11.t2 10.5739
R514 rseg_1_v3_1.v11 rseg_1_v3_1.v11.n0 2.84608
R515 rseg_1_v3_1.v10 rseg_1_v3_1.v10.t1 250.332
R516 rseg_1_v3_1.v10.n0 rseg_1_v3_1.v10.t2 10.5307
R517 rseg_1_v3_1.v10.n0 rseg_1_v3_1.v10.t0 10.5295
R518 rseg_1_v3_1.v10 rseg_1_v3_1.v10.n0 3.51046
R519 DEC[2].n6 DEC[2].t11 213.218
R520 DEC[2].n11 DEC[2].t4 213.218
R521 DEC[2].n0 DEC[2].t14 213.218
R522 DEC[2].n6 DEC[2].t8 212.554
R523 DEC[2].n7 DEC[2].t0 212.554
R524 DEC[2].n8 DEC[2].t12 212.554
R525 DEC[2].n9 DEC[2].t9 212.554
R526 DEC[2].n10 DEC[2].t1 212.554
R527 DEC[2].n5 DEC[2].t10 212.554
R528 DEC[2].n4 DEC[2].t7 212.554
R529 DEC[2].n3 DEC[2].t5 212.554
R530 DEC[2].n2 DEC[2].t2 212.554
R531 DEC[2].n1 DEC[2].t15 212.554
R532 DEC[2].n0 DEC[2].t3 212.554
R533 DEC[2].n13 DEC[2].t13 208.054
R534 DEC[2].n12 DEC[2].t6 208.054
R535 DEC[2].n12 DEC[2].n11 4.5005
R536 DEC[2].n14 DEC[2].n13 4.5005
R537 DEC[2].n13 DEC[2].n12 2.59281
R538 DEC[2].n11 DEC[2].n10 0.663962
R539 DEC[2].n10 DEC[2].n9 0.663962
R540 DEC[2].n9 DEC[2].n8 0.663962
R541 DEC[2].n8 DEC[2].n7 0.663962
R542 DEC[2].n7 DEC[2].n6 0.663962
R543 DEC[2].n1 DEC[2].n0 0.663962
R544 DEC[2].n2 DEC[2].n1 0.663962
R545 DEC[2].n3 DEC[2].n2 0.663962
R546 DEC[2].n4 DEC[2].n3 0.663962
R547 DEC[2].n5 DEC[2].n4 0.663962
R548 DEC[2].n14 DEC[2].n5 0.663962
R549 DEC[2] DEC[2].n14 0.291365
R550 a_337_4028.n1 a_337_4028.t4 247.736
R551 a_337_4028.n0 a_337_4028.t1 245.752
R552 a_337_4028.t0 a_337_4028.n2 245.172
R553 a_337_4028.n1 a_337_4028.t3 239.083
R554 a_337_4028.n0 a_337_4028.t2 239.083
R555 a_337_4028.n2 a_337_4028.n0 5.85467
R556 a_337_4028.n2 a_337_4028.n1 1.16717
R557 rseg_1_v3_1.v34 rseg_1_v3_1.v34.t1 246.804
R558 rseg_1_v3_1.v34.n0 rseg_1_v3_1.v34.t0 10.6257
R559 rseg_1_v3_1.v34.n0 rseg_1_v3_1.v34.t2 10.5285
R560 rseg_1_v3_1.v34 rseg_1_v3_1.v34.n0 0.86158
R561 a_3049_5464.n0 a_3049_5464.t4 246.429
R562 a_3049_5464.t0 a_3049_5464.n2 241.959
R563 a_3049_5464.n2 a_3049_5464.t1 239.822
R564 a_3049_5464.n0 a_3049_5464.t3 239.143
R565 a_3049_5464.n1 a_3049_5464.t2 239.143
R566 a_3049_5464.n1 a_3049_5464.n0 6.788
R567 a_3049_5464.n2 a_3049_5464.n1 3.76508
R568 rseg_1_v3_1.v37 rseg_1_v3_1.v37.t2 246.63
R569 rseg_1_v3_1.v37.n0 rseg_1_v3_1.v37.t1 10.575
R570 rseg_1_v3_1.v37.n0 rseg_1_v3_1.v37.t0 10.5739
R571 rseg_1_v3_1.v37 rseg_1_v3_1.v37.n0 2.81913
R572 a_1323_4028.n2 a_1323_4028.t4 248.286
R573 a_1323_4028.n0 a_1323_4028.t2 246.303
R574 a_1323_4028.n1 a_1323_4028.t1 244.629
R575 a_1323_4028.n0 a_1323_4028.t3 239.633
R576 a_1323_4028.t0 a_1323_4028.n2 239.633
R577 a_1323_4028.n2 a_1323_4028.n1 5.93592
R578 a_1323_4028.n1 a_1323_4028.n0 1.08592
R579 bb[3].n2 bb[3].t0 213.218
R580 bb[3].n0 bb[3].t3 213.218
R581 bb[3].n2 bb[3].t7 212.554
R582 bb[3].n3 bb[3].t1 212.554
R583 bb[3].n4 bb[3].t4 212.554
R584 bb[3].n5 bb[3].t2 212.554
R585 bb[3].n1 bb[3].t6 212.554
R586 bb[3].n0 bb[3].t5 212.554
R587 bb[3].n1 bb[3].n0 0.663962
R588 bb[3].n5 bb[3].n4 0.663962
R589 bb[3].n4 bb[3].n3 0.663962
R590 bb[3].n3 bb[3].n2 0.663962
R591 bb[3] bb[3].n5 0.541365
R592 bb[3] bb[3].n1 0.123096
R593 a_n215_4028.n2 a_n215_4028.t2 247.369
R594 a_n215_4028.n0 a_n215_4028.t4 245.386
R595 a_n215_4028.n1 a_n215_4028.t3 244.766
R596 a_n215_4028.n0 a_n215_4028.t1 238.716
R597 a_n215_4028.t0 a_n215_4028.n2 238.716
R598 a_n215_4028.n1 a_n215_4028.n0 5.07133
R599 a_n215_4028.n2 a_n215_4028.n1 1.9505
R600 a_5799_6728.n0 a_5799_6728.t2 244.542
R601 a_5799_6728.n0 a_5799_6728.t1 242.81
R602 a_5799_6728.t0 a_5799_6728.n0 239.857
R603 a_2773_5464.n0 a_2773_5464.t4 246.244
R604 a_2773_5464.n2 a_2773_5464.t1 241.385
R605 a_2773_5464.t0 a_2773_5464.n2 240.358
R606 a_2773_5464.n0 a_2773_5464.t2 238.959
R607 a_2773_5464.n1 a_2773_5464.t3 238.959
R608 a_2773_5464.n1 a_2773_5464.n0 6.788
R609 a_2773_5464.n2 a_2773_5464.n1 4.15675
R610 rseg_1_v3_1.v44 rseg_1_v3_1.v44.t0 249.209
R611 rseg_1_v3_1.v44.n0 rseg_1_v3_1.v44.t1 10.5296
R612 rseg_1_v3_1.v44.n0 rseg_1_v3_1.v44.t2 10.5285
R613 rseg_1_v3_1.v44 rseg_1_v3_1.v44.n0 2.13671
R614 a_3483_5464.n2 a_3483_5464.t2 246.612
R615 a_3483_5464.n0 a_3483_5464.t4 242.863
R616 a_3483_5464.n0 a_3483_5464.t3 239.639
R617 a_3483_5464.n1 a_3483_5464.t1 239.326
R618 a_3483_5464.t0 a_3483_5464.n2 239.326
R619 a_3483_5464.n2 a_3483_5464.n1 6.788
R620 a_3483_5464.n1 a_3483_5464.n0 3.04425
R621 rseg_1_v3_1.v61 rseg_1_v3_1.v61.t2 249.321
R622 rseg_1_v3_1.v61.n0 rseg_1_v3_1.v61.t1 10.6701
R623 rseg_1_v3_1.v61.n0 rseg_1_v3_1.v61.t0 10.5739
R624 rseg_1_v3_1.v61 rseg_1_v3_1.v61.n0 1.53658
R625 rseg_1_v3_1.v60 rseg_1_v3_1.v60.t2 249.148
R626 rseg_1_v3_1.v60.n0 rseg_1_v3_1.v60.t0 10.6257
R627 rseg_1_v3_1.v60.n0 rseg_1_v3_1.v60.t1 10.5285
R628 rseg_1_v3_1.v60 rseg_1_v3_1.v60.n0 2.09277
R629 rseg_1_v3_1.v13 rseg_1_v3_1.v13.t1 249.321
R630 rseg_1_v3_1.v13.n0 rseg_1_v3_1.v13.t2 10.575
R631 rseg_1_v3_1.v13.n0 rseg_1_v3_1.v13.t0 10.5739
R632 rseg_1_v3_1.v13 rseg_1_v3_1.v13.n0 1.60689
R633 rseg_1_v3_1.v12 rseg_1_v3_1.v12.t2 249.594
R634 rseg_1_v3_1.v12.n0 rseg_1_v3_1.v12.t0 10.5317
R635 rseg_1_v3_1.v12.n0 rseg_1_v3_1.v12.t1 10.5285
R636 rseg_1_v3_1.v12 rseg_1_v3_1.v12.n0 2.17402
R637 DEC[3].n6 DEC[3].t5 213.218
R638 DEC[3].n11 DEC[3].t13 213.218
R639 DEC[3].n0 DEC[3].t9 213.218
R640 DEC[3].n6 DEC[3].t3 212.554
R641 DEC[3].n7 DEC[3].t2 212.554
R642 DEC[3].n8 DEC[3].t6 212.554
R643 DEC[3].n9 DEC[3].t4 212.554
R644 DEC[3].n10 DEC[3].t10 212.554
R645 DEC[3].n5 DEC[3].t14 212.554
R646 DEC[3].n4 DEC[3].t11 212.554
R647 DEC[3].n3 DEC[3].t1 212.554
R648 DEC[3].n2 DEC[3].t15 212.554
R649 DEC[3].n1 DEC[3].t12 212.554
R650 DEC[3].n0 DEC[3].t8 212.554
R651 DEC[3].n13 DEC[3].t7 208.054
R652 DEC[3].n12 DEC[3].t0 208.054
R653 DEC[3].n12 DEC[3].n11 4.5005
R654 DEC[3].n14 DEC[3].n13 4.5005
R655 DEC[3].n13 DEC[3].n12 2.588
R656 DEC[3].n11 DEC[3].n10 0.663962
R657 DEC[3].n10 DEC[3].n9 0.663962
R658 DEC[3].n9 DEC[3].n8 0.663962
R659 DEC[3].n8 DEC[3].n7 0.663962
R660 DEC[3].n7 DEC[3].n6 0.663962
R661 DEC[3].n1 DEC[3].n0 0.663962
R662 DEC[3].n2 DEC[3].n1 0.663962
R663 DEC[3].n3 DEC[3].n2 0.663962
R664 DEC[3].n4 DEC[3].n3 0.663962
R665 DEC[3].n5 DEC[3].n4 0.663962
R666 DEC[3].n14 DEC[3].n5 0.663962
R667 DEC[3] DEC[3].n14 0.313
R668 rseg_1_v3_1.v54 rseg_1_v3_1.v54.t0 246.798
R669 rseg_1_v3_1.v54.n0 rseg_1_v3_1.v54.t2 10.6247
R670 rseg_1_v3_1.v54.n0 rseg_1_v3_1.v54.t1 10.5285
R671 rseg_1_v3_1.v54 rseg_1_v3_1.v54.n0 3.49191
R672 a_1599_4028.n2 a_1599_4028.t3 248.469
R673 a_1599_4028.n0 a_1599_4028.t1 246.486
R674 a_1599_4028.n1 a_1599_4028.t4 244.054
R675 a_1599_4028.n0 a_1599_4028.t2 239.816
R676 a_1599_4028.t0 a_1599_4028.n2 239.816
R677 a_1599_4028.n2 a_1599_4028.n1 5.54425
R678 a_1599_4028.n1 a_1599_4028.n0 1.47758
R679 b[2].n1 b[2].t2 213.218
R680 b[2].n0 b[2].t0 213.218
R681 b[2].n1 b[2].t3 212.554
R682 b[2].n0 b[2].t1 212.554
R683 b[2] b[2].n1 0.380308
R684 b[2] b[2].n0 0.284154
R685 a_7573_6728.n0 a_7573_6728.t2 246.316
R686 a_7573_6728.t0 a_7573_6728.n0 244.469
R687 a_7573_6728.n0 a_7573_6728.t1 238.573
R688 a_7618_7809.t0 a_7618_7809.n0 243.633
R689 a_7618_7809.n0 a_7618_7809.t2 241.625
R690 a_7618_7809.n0 a_7618_7809.t1 239.267
R691 rseg_1_v3_1.v39 rseg_1_v3_1.v39.t1 248.075
R692 rseg_1_v3_1.v39.n0 rseg_1_v3_1.v39.t0 10.575
R693 rseg_1_v3_1.v39.n0 rseg_1_v3_1.v39.t2 10.5739
R694 rseg_1_v3_1.v39 rseg_1_v3_1.v39.n0 4.2135
R695 rseg_1_v3_1.v40 rseg_1_v3_1.v40.t1 249.738
R696 rseg_1_v3_1.v40.n0 rseg_1_v3_1.v40.t2 13.4746
R697 rseg_1_v3_1.v40.n0 rseg_1_v3_1.v40.t0 10.7886
R698 rseg_1_v3_1.v40 rseg_1_v3_1.v40.n0 4.72836
R699 rseg_1_v3_1.v3 rseg_1_v3_1.v3.t2 245.726
R700 rseg_1_v3_1.v3.n0 rseg_1_v3_1.v3.t1 10.5816
R701 rseg_1_v3_1.v3.n0 rseg_1_v3_1.v3.t0 10.5739
R702 rseg_1_v3_1.v3 rseg_1_v3_1.v3.n0 1.48638
R703 rseg_1_v3_1.v4 rseg_1_v3_1.v4.t2 247.869
R704 rseg_1_v3_1.v4.n0 rseg_1_v3_1.v4.t1 10.5339
R705 rseg_1_v3_1.v4.n0 rseg_1_v3_1.v4.t0 10.5295
R706 rseg_1_v3_1.v4 rseg_1_v3_1.v4.n0 2.21785
R707 rseg_1_v3_1.v15.n0 rseg_1_v3_1.v15.t2 240.469
R708 rseg_1_v3_1.v15.n0 rseg_1_v3_1.v15.t1 10.6713
R709 rseg_1_v3_1.v15.t0 rseg_1_v3_1.v15.n0 10.5739
R710 rseg_1_v3_1.v16.t0 rseg_1_v3_1.v16.n0 241.547
R711 rseg_1_v3_1.v16.n0 rseg_1_v3_1.v16.t2 12.2056
R712 rseg_1_v3_1.v16.n0 rseg_1_v3_1.v16.t1 12.0758
R713 rseg_1_v3_1.v46 rseg_1_v3_1.v46.t1 249.239
R714 rseg_1_v3_1.v46.n0 rseg_1_v3_1.v46.t0 10.6257
R715 rseg_1_v3_1.v46.n0 rseg_1_v3_1.v46.t2 10.5285
R716 rseg_1_v3_1.v46 rseg_1_v3_1.v46.n0 0.872789
R717 a_4035_5464.n0 a_4035_5464.t4 246.978
R718 a_4035_5464.t0 a_4035_5464.n2 244.013
R719 a_4035_5464.n2 a_4035_5464.t2 240.072
R720 a_4035_5464.n0 a_4035_5464.t1 239.692
R721 a_4035_5464.n1 a_4035_5464.t3 239.692
R722 a_4035_5464.n1 a_4035_5464.n0 6.788
R723 a_4035_5464.n2 a_4035_5464.n1 2.26092
R724 bb[1] bb[1].t1 213.042
R725 bb[1] bb[1].t0 212.73
R726 a_7010_7809.n0 a_7010_7809.t2 240.108
R727 a_7010_7809.n0 a_7010_7809.t1 239.733
R728 a_7010_7809.t0 a_7010_7809.n0 238.899
R729 a_8198_7809.n0 a_8198_7809.t2 241.258
R730 a_8198_7809.n0 a_8198_7809.t1 240.909
R731 a_8198_7809.t0 a_8198_7809.n0 238.899
R732 rseg_1_v3_1.v59 rseg_1_v3_1.v59.t1 248.95
R733 rseg_1_v3_1.v59.n0 rseg_1_v3_1.v59.t0 10.6701
R734 rseg_1_v3_1.v59.n0 rseg_1_v3_1.v59.t2 10.5739
R735 rseg_1_v3_1.v59 rseg_1_v3_1.v59.n0 2.77016
R736 rseg_1_v3_1.v49.n0 rseg_1_v3_1.v49.t1 236.649
R737 rseg_1_v3_1.v49.t0 rseg_1_v3_1.v49.n0 10.6713
R738 rseg_1_v3_1.v49.n0 rseg_1_v3_1.v49.t2 10.5739
R739 rseg_1_v3_1.v50 rseg_1_v3_1.v50.t1 246.716
R740 rseg_1_v3_1.v50.n0 rseg_1_v3_1.v50.t2 10.5296
R741 rseg_1_v3_1.v50.n0 rseg_1_v3_1.v50.t0 10.5295
R742 rseg_1_v3_1.v50 rseg_1_v3_1.v50.n0 0.886534
R743 bb[0] bb[0].t0 212.614
R744 VOUT VOUT.t1 239.155
R745 VOUT VOUT.t0 238.912
R746 a_7314_7809.n0 a_7314_7809.t1 240.13
R747 a_7314_7809.n0 a_7314_7809.t2 239.512
R748 a_7314_7809.t0 a_7314_7809.n0 238.921
R749 bb[2].n1 bb[2].t1 213.218
R750 bb[2].n0 bb[2].t3 213.218
R751 bb[2].n1 bb[2].t0 212.554
R752 bb[2].n0 bb[2].t2 212.554
R753 bb[2] bb[2].n0 0.445212
R754 bb[2] bb[2].n1 0.21925
R755 a_6075_6728.n0 a_6075_6728.t2 244.725
R756 a_6075_6728.t0 a_6075_6728.n0 242.994
R757 a_6075_6728.n0 a_6075_6728.t1 239.673
R758 rseg_1_v3_1.v6 rseg_1_v3_1.v6.t2 248.484
R759 rseg_1_v3_1.v6.n0 rseg_1_v3_1.v6.t0 10.5338
R760 rseg_1_v3_1.v6.n0 rseg_1_v3_1.v6.t1 10.5285
R761 rseg_1_v3_1.v6 rseg_1_v3_1.v6.n0 3.63285
R762 rseg_1_v3_1.v8 rseg_1_v3_1.v8.t2 249.738
R763 rseg_1_v3_1.v8.n0 rseg_1_v3_1.v8.t0 13.5854
R764 rseg_1_v3_1.v8.n0 rseg_1_v3_1.v8.t1 10.8954
R765 rseg_1_v3_1.v8 rseg_1_v3_1.v8.n0 4.7255
R766 a_2497_5464.n0 a_2497_5464.t3 246.061
R767 a_2497_5464.t0 a_2497_5464.n2 240.989
R768 a_2497_5464.n2 a_2497_5464.t1 240.81
R769 a_2497_5464.n0 a_2497_5464.t4 238.775
R770 a_2497_5464.n1 a_2497_5464.t2 238.775
R771 a_2497_5464.n1 a_2497_5464.n0 6.788
R772 a_2497_5464.n2 a_2497_5464.n1 4.54842
R773 rseg_1_v3_1.v9 rseg_1_v3_1.v9.t2 249.345
R774 rseg_1_v3_1.v9.n0 rseg_1_v3_1.v9.t0 10.5773
R775 rseg_1_v3_1.v9.n0 rseg_1_v3_1.v9.t1 10.5739
R776 rseg_1_v3_1.v9 rseg_1_v3_1.v9.n0 4.18158
R777 a_6351_6728.n0 a_6351_6728.t2 244.909
R778 a_6351_6728.t0 a_6351_6728.n0 243.178
R779 a_6351_6728.n0 a_6351_6728.t1 239.489
R780 V0.n0 V0.t1 241.547
R781 V0.n0 V0.t0 12.5185
R782 V0 V0.n0 0.274355
R783 rseg_1_v3_1.v57 rseg_1_v3_1.v57.t0 249.345
R784 rseg_1_v3_1.v57.n0 rseg_1_v3_1.v57.t2 10.575
R785 rseg_1_v3_1.v57.n0 rseg_1_v3_1.v57.t1 10.5739
R786 rseg_1_v3_1.v57 rseg_1_v3_1.v57.n0 4.20587
R787 rseg_1_v3_1.v58 rseg_1_v3_1.v58.t1 249.886
R788 rseg_1_v3_1.v58.n0 rseg_1_v3_1.v58.t2 10.6247
R789 rseg_1_v3_1.v58.n0 rseg_1_v3_1.v58.t0 10.5295
R790 rseg_1_v3_1.v58 rseg_1_v3_1.v58.n0 3.48476
R791 a_61_4028.n0 a_61_4028.t3 247.553
R792 a_61_4028.t0 a_61_4028.n2 245.569
R793 a_61_4028.n1 a_61_4028.t4 244.964
R794 a_61_4028.n0 a_61_4028.t1 238.899
R795 a_61_4028.n2 a_61_4028.t2 238.899
R796 a_61_4028.n2 a_61_4028.n1 5.463
R797 a_61_4028.n1 a_61_4028.n0 1.55883
R798 rseg_1_v3_1.v52 rseg_1_v3_1.v52.t2 246.18
R799 rseg_1_v3_1.v52.n0 rseg_1_v3_1.v52.t1 10.5296
R800 rseg_1_v3_1.v52.n0 rseg_1_v3_1.v52.t0 10.5295
R801 rseg_1_v3_1.v52 rseg_1_v3_1.v52.n0 2.14387
R802 a_1047_4028.n0 a_1047_4028.t3 248.102
R803 a_1047_4028.t0 a_1047_4028.n2 246.119
R804 a_1047_4028.n1 a_1047_4028.t4 245.203
R805 a_1047_4028.n0 a_1047_4028.t2 239.45
R806 a_1047_4028.n2 a_1047_4028.t1 239.45
R807 a_1047_4028.n1 a_1047_4028.n0 6.32758
R808 a_1047_4028.n2 a_1047_4028.n1 0.69425
R809 rseg_1_v3_1.v47.n0 rseg_1_v3_1.v47.t1 240.469
R810 rseg_1_v3_1.v47.n0 rseg_1_v3_1.v47.t2 10.6713
R811 rseg_1_v3_1.v47.t0 rseg_1_v3_1.v47.n0 10.5739
R812 rseg_1_v3_1.v48.t0 rseg_1_v3_1.v48.n0 241.547
R813 rseg_1_v3_1.v48.n0 rseg_1_v3_1.v48.t2 12.1321
R814 rseg_1_v3_1.v48.n0 rseg_1_v3_1.v48.t1 12.0758
R815 b[3].n0 b[3].t0 213.218
R816 b[3] b[3].t5 212.77
R817 b[3].n5 b[3].t3 212.554
R818 b[3].n4 b[3].t7 212.554
R819 b[3].n3 b[3].t6 212.554
R820 b[3].n2 b[3].t4 212.554
R821 b[3].n1 b[3].t2 212.554
R822 b[3].n0 b[3].t1 212.554
R823 b[3].n1 b[3].n0 0.663962
R824 b[3].n2 b[3].n1 0.663962
R825 b[3].n3 b[3].n2 0.663962
R826 b[3].n4 b[3].n3 0.663962
R827 b[3].n5 b[3].n4 0.663962
R828 b[3] b[3].n5 0.447615
R829 a_4311_5464.n2 a_4311_5464.t4 247.161
R830 a_4311_5464.n0 a_4311_5464.t1 244.589
R831 a_4311_5464.n0 a_4311_5464.t3 240.337
R832 a_4311_5464.n1 a_4311_5464.t2 239.875
R833 a_4311_5464.t0 a_4311_5464.n2 239.875
R834 a_4311_5464.n2 a_4311_5464.n1 6.788
R835 a_4311_5464.n1 a_4311_5464.n0 1.86925
R836 rseg_1_v3_1.v14 rseg_1_v3_1.v14.t1 249.623
R837 rseg_1_v3_1.v14.n0 rseg_1_v3_1.v14.t0 10.5319
R838 rseg_1_v3_1.v14.n0 rseg_1_v3_1.v14.t2 10.5285
R839 rseg_1_v3_1.v14 rseg_1_v3_1.v14.n0 0.915451
R840 rseg_1_v3_1.v23 rseg_1_v3_1.v23.t1 248.075
R841 rseg_1_v3_1.v23.n0 rseg_1_v3_1.v23.t0 10.6701
R842 rseg_1_v3_1.v23.n0 rseg_1_v3_1.v23.t2 10.5739
R843 rseg_1_v3_1.v23 rseg_1_v3_1.v23.n0 4.17455
R844 rseg_1_v3_1.v24 rseg_1_v3_1.v24.t0 249.738
R845 rseg_1_v3_1.v24.n0 rseg_1_v3_1.v24.t2 13.5018
R846 rseg_1_v3_1.v24.n0 rseg_1_v3_1.v24.t1 10.7924
R847 rseg_1_v3_1.v24 rseg_1_v3_1.v24.n0 4.72836
R848 a_8474_7809.n0 a_8474_7809.t2 241.075
R849 a_8474_7809.t0 a_8474_7809.n0 239.35
R850 a_8474_7809.n0 a_8474_7809.t1 238.716
R851 rseg_1_v3_1.v27 rseg_1_v3_1.v27.t2 248.95
R852 rseg_1_v3_1.v27.n0 rseg_1_v3_1.v27.t0 10.6701
R853 rseg_1_v3_1.v27.n0 rseg_1_v3_1.v27.t1 10.5739
R854 rseg_1_v3_1.v27 rseg_1_v3_1.v27.n0 2.76539
R855 rseg_1_v3_1.v28 rseg_1_v3_1.v28.t0 249.328
R856 rseg_1_v3_1.v28.n0 rseg_1_v3_1.v28.t2 10.5296
R857 rseg_1_v3_1.v28.n0 rseg_1_v3_1.v28.t1 10.5285
R858 rseg_1_v3_1.v28 rseg_1_v3_1.v28.n0 2.13671
R859 rseg_1_v3_1.v5 rseg_1_v3_1.v5.t2 246.63
R860 rseg_1_v3_1.v5.n0 rseg_1_v3_1.v5.t0 10.5795
R861 rseg_1_v3_1.v5.n0 rseg_1_v3_1.v5.t1 10.5739
R862 rseg_1_v3_1.v5 rseg_1_v3_1.v5.n0 2.90483
R863 rseg_1_v3_1.v43 rseg_1_v3_1.v43.t0 248.95
R864 rseg_1_v3_1.v43.n0 rseg_1_v3_1.v43.t1 10.575
R865 rseg_1_v3_1.v43.n0 rseg_1_v3_1.v43.t2 10.5739
R866 rseg_1_v3_1.v43 rseg_1_v3_1.v43.n0 2.81389
R867 DEC[1].n6 DEC[1].t10 213.218
R868 DEC[1].n11 DEC[1].t14 213.218
R869 DEC[1].n0 DEC[1].t15 213.218
R870 DEC[1].n6 DEC[1].t12 212.554
R871 DEC[1].n7 DEC[1].t4 212.554
R872 DEC[1].n8 DEC[1].t0 212.554
R873 DEC[1].n9 DEC[1].t9 212.554
R874 DEC[1].n10 DEC[1].t5 212.554
R875 DEC[1].n5 DEC[1].t13 212.554
R876 DEC[1].n4 DEC[1].t6 212.554
R877 DEC[1].n3 DEC[1].t2 212.554
R878 DEC[1].n2 DEC[1].t8 212.554
R879 DEC[1].n1 DEC[1].t7 212.554
R880 DEC[1].n0 DEC[1].t3 212.554
R881 DEC[1].n13 DEC[1].t11 208.054
R882 DEC[1].n12 DEC[1].t1 208.054
R883 DEC[1].n12 DEC[1].n11 4.5005
R884 DEC[1].n14 DEC[1].n13 4.5005
R885 DEC[1].n13 DEC[1].n12 2.97742
R886 DEC[1].n11 DEC[1].n10 0.663962
R887 DEC[1].n10 DEC[1].n9 0.663962
R888 DEC[1].n9 DEC[1].n8 0.663962
R889 DEC[1].n8 DEC[1].n7 0.663962
R890 DEC[1].n7 DEC[1].n6 0.663962
R891 DEC[1].n1 DEC[1].n0 0.663962
R892 DEC[1].n2 DEC[1].n1 0.663962
R893 DEC[1].n3 DEC[1].n2 0.663962
R894 DEC[1].n4 DEC[1].n3 0.663962
R895 DEC[1].n5 DEC[1].n4 0.663962
R896 DEC[1].n14 DEC[1].n5 0.663962
R897 DEC[1] DEC[1].n14 0.269731
R898 a_613_4028.n2 a_613_4028.t3 247.918
R899 a_613_4028.n0 a_613_4028.t1 245.935
R900 a_613_4028.n1 a_613_4028.t4 245.381
R901 a_613_4028.n0 a_613_4028.t2 239.267
R902 a_613_4028.t0 a_613_4028.n2 239.267
R903 a_613_4028.n1 a_613_4028.n0 6.24633
R904 a_613_4028.n2 a_613_4028.n1 0.7755
R905 rseg_1_v3_1.v19 rseg_1_v3_1.v19.t0 245.726
R906 rseg_1_v3_1.v19.n0 rseg_1_v3_1.v19.t1 10.6701
R907 rseg_1_v3_1.v19.n0 rseg_1_v3_1.v19.t2 10.5739
R908 rseg_1_v3_1.v19 rseg_1_v3_1.v19.n0 1.51759
R909 rseg_1_v3_1.v38 rseg_1_v3_1.v38.t1 246.885
R910 rseg_1_v3_1.v38.n0 rseg_1_v3_1.v38.t2 10.5296
R911 rseg_1_v3_1.v38.n0 rseg_1_v3_1.v38.t0 10.5295
R912 rseg_1_v3_1.v38 rseg_1_v3_1.v38.n0 3.53633
R913 a_2221_5464.n2 a_2221_5464.t4 245.879
R914 a_2221_5464.n0 a_2221_5464.t3 241.619
R915 a_2221_5464.n0 a_2221_5464.t1 240.234
R916 a_2221_5464.n1 a_2221_5464.t2 238.593
R917 a_2221_5464.t0 a_2221_5464.n2 238.593
R918 a_2221_5464.n2 a_2221_5464.n1 6.788
R919 a_2221_5464.n1 a_2221_5464.n0 4.94008
R920 rseg_1_v3_1.v22 rseg_1_v3_1.v22.t0 247.119
R921 rseg_1_v3_1.v22.n0 rseg_1_v3_1.v22.t2 10.5296
R922 rseg_1_v3_1.v22.n0 rseg_1_v3_1.v22.t1 10.5285
R923 rseg_1_v3_1.v22 rseg_1_v3_1.v22.n0 3.54349
R924 rseg_1_v3_1.v25 rseg_1_v3_1.v25.t0 249.345
R925 rseg_1_v3_1.v25.n0 rseg_1_v3_1.v25.t1 10.6701
R926 rseg_1_v3_1.v25.n0 rseg_1_v3_1.v25.t2 10.5739
R927 rseg_1_v3_1.v25 rseg_1_v3_1.v25.n0 4.15498
R928 rseg_1_v3_1.v26 rseg_1_v3_1.v26.t1 250.066
R929 rseg_1_v3_1.v26.n0 rseg_1_v3_1.v26.t0 10.5306
R930 rseg_1_v3_1.v26.n0 rseg_1_v3_1.v26.t2 10.5285
R931 rseg_1_v3_1.v26 rseg_1_v3_1.v26.n0 3.52631
R932 rseg_1_v3_1.v21 rseg_1_v3_1.v21.t1 246.63
R933 rseg_1_v3_1.v21.n0 rseg_1_v3_1.v21.t2 10.6701
R934 rseg_1_v3_1.v21.n0 rseg_1_v3_1.v21.t0 10.5739
R935 rseg_1_v3_1.v21 rseg_1_v3_1.v21.n0 2.78018
R936 rseg_1_v3_1.v20 rseg_1_v3_1.v20.t1 246.501
R937 rseg_1_v3_1.v20.n0 rseg_1_v3_1.v20.t0 10.5319
R938 rseg_1_v3_1.v20.n0 rseg_1_v3_1.v20.t2 10.5285
R939 rseg_1_v3_1.v20 rseg_1_v3_1.v20.n0 2.14784
R940 rseg_1_v3_1.v51 rseg_1_v3_1.v51.t1 245.726
R941 rseg_1_v3_1.v51.n0 rseg_1_v3_1.v51.t2 10.575
R942 rseg_1_v3_1.v51.n0 rseg_1_v3_1.v51.t0 10.5739
R943 rseg_1_v3_1.v51 rseg_1_v3_1.v51.n0 1.5626
R944 rseg_1_v3_1.v1.n0 rseg_1_v3_1.v1.t2 236.657
R945 rseg_1_v3_1.v1.t0 rseg_1_v3_1.v1.n0 10.6906
R946 rseg_1_v3_1.v1.n0 rseg_1_v3_1.v1.t1 10.5739
R947 rseg_1_v3_1.v2 rseg_1_v3_1.v2.t2 248.405
R948 rseg_1_v3_1.v2.n0 rseg_1_v3_1.v2.t1 10.5394
R949 rseg_1_v3_1.v2.n0 rseg_1_v3_1.v2.t0 10.5295
R950 rseg_1_v3_1.v2 rseg_1_v3_1.v2.n0 0.791214
R951 rseg_1_v3_1.v41 rseg_1_v3_1.v41.t0 249.345
R952 rseg_1_v3_1.v41.n0 rseg_1_v3_1.v41.t1 10.575
R953 rseg_1_v3_1.v41.n0 rseg_1_v3_1.v41.t2 10.5739
R954 rseg_1_v3_1.v41 rseg_1_v3_1.v41.n0 4.20348
R955 rseg_1_v3_1.v30 rseg_1_v3_1.v30.t0 249.358
R956 rseg_1_v3_1.v30.n0 rseg_1_v3_1.v30.t1 10.5296
R957 rseg_1_v3_1.v30.n0 rseg_1_v3_1.v30.t2 10.5285
R958 rseg_1_v3_1.v30 rseg_1_v3_1.v30.n0 0.905521
R959 rseg_1_v3_1.v35 rseg_1_v3_1.v35.t2 245.728
R960 rseg_1_v3_1.v35.n0 rseg_1_v3_1.v35.t0 10.5752
R961 rseg_1_v3_1.v35.n0 rseg_1_v3_1.v35.t1 10.5739
R962 rseg_1_v3_1.v35 rseg_1_v3_1.v35.n0 1.55257
R963 rseg_1_v3_1.v36 rseg_1_v3_1.v36.t2 246.268
R964 rseg_1_v3_1.v36.n0 rseg_1_v3_1.v36.t1 10.5296
R965 rseg_1_v3_1.v36.n0 rseg_1_v3_1.v36.t0 10.5295
R966 rseg_1_v3_1.v36 rseg_1_v3_1.v36.n0 2.15701
R967 a_7297_6728.n0 a_7297_6728.t2 246.133
R968 a_7297_6728.t0 a_7297_6728.n0 244.286
R969 a_7297_6728.n0 a_7297_6728.t1 238.756
R970 rseg_1_v3_1.v56 rseg_1_v3_1.v56.t0 249.738
R971 rseg_1_v3_1.v56.n0 rseg_1_v3_1.v56.t1 13.4579
R972 rseg_1_v3_1.v56.n0 rseg_1_v3_1.v56.t2 10.7848
R973 rseg_1_v3_1.v56 rseg_1_v3_1.v56.n0 4.72836
R974 a_7894_7809.t0 a_7894_7809.n0 242.075
R975 a_7894_7809.n0 a_7894_7809.t2 241.441
R976 a_7894_7809.n0 a_7894_7809.t1 239.083
R977 rseg_1_v3_1.v18 rseg_1_v3_1.v18.t1 247.037
R978 rseg_1_v3_1.v18.n0 rseg_1_v3_1.v18.t2 10.5307
R979 rseg_1_v3_1.v18.n0 rseg_1_v3_1.v18.t0 10.5295
R980 rseg_1_v3_1.v18 rseg_1_v3_1.v18.n0 0.885467
R981 b[1] b[1].t1 212.911
R982 b[1] b[1].t0 212.863
R983 rseg_1_v3_1.v42 rseg_1_v3_1.v42.t0 249.947
R984 rseg_1_v3_1.v42.n0 rseg_1_v3_1.v42.t2 10.5296
R985 rseg_1_v3_1.v42.n0 rseg_1_v3_1.v42.t1 10.5285
R986 rseg_1_v3_1.v42 rseg_1_v3_1.v42.n0 3.5287
R987 rseg_1_v3_1.v33.n0 rseg_1_v3_1.v33.t1 236.65
R988 rseg_1_v3_1.v33.n0 rseg_1_v3_1.v33.t2 10.6732
R989 rseg_1_v3_1.v33.t0 rseg_1_v3_1.v33.n0 10.5739
R990 rseg_1_v3_1.v55 rseg_1_v3_1.v55.t0 248.075
R991 rseg_1_v3_1.v55.n0 rseg_1_v3_1.v55.t2 10.6701
R992 rseg_1_v3_1.v55.n0 rseg_1_v3_1.v55.t1 10.5739
R993 rseg_1_v3_1.v55 rseg_1_v3_1.v55.n0 4.16691
R994 rseg_1_v3_1.v29 rseg_1_v3_1.v29.t0 249.321
R995 rseg_1_v3_1.v29.n0 rseg_1_v3_1.v29.t2 10.6701
R996 rseg_1_v3_1.v29.n0 rseg_1_v3_1.v29.t1 10.5739
R997 rseg_1_v3_1.v29 rseg_1_v3_1.v29.n0 1.54779
R998 a_3759_5464.n2 a_3759_5464.t4 246.794
R999 a_3759_5464.n0 a_3759_5464.t1 243.439
R1000 a_3759_5464.n0 a_3759_5464.t3 239.809
R1001 a_3759_5464.n1 a_3759_5464.t2 239.51
R1002 a_3759_5464.t0 a_3759_5464.n2 239.51
R1003 a_3759_5464.n2 a_3759_5464.n1 6.788
R1004 a_3759_5464.n1 a_3759_5464.n0 2.65258
R1005 a_7021_6728.n0 a_7021_6728.t2 245.95
R1006 a_7021_6728.t0 a_7021_6728.n0 244.102
R1007 a_7021_6728.n0 a_7021_6728.t1 238.94
R1008 a_6745_6728.n0 a_6745_6728.t2 245.95
R1009 a_6745_6728.t0 a_6745_6728.n0 243.918
R1010 a_6745_6728.n0 a_6745_6728.t1 239.124
R1011 rseg_1_v3_1.v32.n0 rseg_1_v3_1.v32.t2 241.547
R1012 rseg_1_v3_1.v32.n0 rseg_1_v3_1.v32.t1 12.1521
R1013 rseg_1_v3_1.v32.t0 rseg_1_v3_1.v32.n0 12.0768
R1014 rseg_1_v3_1.v31.t0 rseg_1_v3_1.v31.n0 240.469
R1015 rseg_1_v3_1.v31.n0 rseg_1_v3_1.v31.t2 10.6701
R1016 rseg_1_v3_1.v31.n0 rseg_1_v3_1.v31.t1 10.5739
R1017 rseg_1_v3_1.v62 rseg_1_v3_1.v62.t1 249.178
R1018 rseg_1_v3_1.v62.n0 rseg_1_v3_1.v62.t0 10.6257
R1019 rseg_1_v3_1.v62.n0 rseg_1_v3_1.v62.t2 10.5285
R1020 rseg_1_v3_1.v62 rseg_1_v3_1.v62.n0 0.872789
R1021 rseg_1_v3_1.v53 rseg_1_v3_1.v53.t1 246.63
R1022 rseg_1_v3_1.v53.n0 rseg_1_v3_1.v53.t2 10.6701
R1023 rseg_1_v3_1.v53.n0 rseg_1_v3_1.v53.t0 10.5739
R1024 rseg_1_v3_1.v53 rseg_1_v3_1.v53.n0 2.77493
R1025 b[0] b[0].t0 212.767
R1026 rseg_1_v3_1.v45 rseg_1_v3_1.v45.t1 249.321
R1027 rseg_1_v3_1.v45.n0 rseg_1_v3_1.v45.t2 10.6671
R1028 rseg_1_v3_1.v45.n0 rseg_1_v3_1.v45.t0 10.5769
R1029 rseg_1_v3_1.v45 rseg_1_v3_1.v45.n0 1.55078
R1030 a_6627_6728.n0 a_6627_6728.t2 245.316
R1031 a_6627_6728.n0 a_6627_6728.t1 243.361
R1032 a_6627_6728.t0 a_6627_6728.n0 239.308
R1033 rseg_1_v3_1.v17.n0 rseg_1_v3_1.v17.t1 236.649
R1034 rseg_1_v3_1.v17.t0 rseg_1_v3_1.v17.n0 10.6701
R1035 rseg_1_v3_1.v17.n0 rseg_1_v3_1.v17.t2 10.5739
R1036 rseg_1_v3_1.v63.t0 rseg_1_v3_1.v63.n0 240.469
R1037 rseg_1_v3_1.v63.n0 rseg_1_v3_1.v63.t2 10.6713
R1038 rseg_1_v3_1.v63.n0 rseg_1_v3_1.v63.t1 10.5739
R1039 V64 V64.t0 11.9718
C0 DEC[1] rseg_1_v3_1.v27 0.09136f
C1 rseg_1_v3_1.v58 rseg_1_v3_1.v60 1.89956f
C2 rseg_1_v3_1.v41 DEC[2] 0.16384f
C3 rseg_1_v3_1.v18 rseg_1_v3_1.v20 1.26125f
C4 rseg_1_v3_1.v58 rseg_1_v3_1.v56 0.55355f
C5 rseg_1_v3_1.v59 rseg_1_v3_1.v54 0.05305f
C6 rseg_1_v3_1.v25 rseg_1_v3_1.v24 3.7974f
C7 rseg_1_v3_1.v9 rseg_1_v3_1.v8 3.76093f
C8 rseg_1_v3_1.v53 rseg_1_v3_1.v55 1.97838f
C9 rseg_1_v3_1.v26 rseg_1_v3_1.v28 1.94958f
C10 rseg_1_v3_1.v25 rseg_1_v3_1.v29 0.08427f
C11 rseg_1_v3_1.v62 rseg_1_v3_1.v60 1.15664f
C12 rseg_1_v3_1.v27 rseg_1_v3_1.v22 0.05302f
C13 rseg_1_v3_1.v42 DEC[2] 0.1787f
C14 rseg_1_v3_1.v50 rseg_1_v3_1.v53 0.04864f
C15 rseg_1_v3_1.v9 rseg_1_v3_1.v12 0.02715f
C16 rseg_1_v3_1.v21 rseg_1_v3_1.v18 0.04809f
C17 rseg_1_v3_1.v57 DEC[3] 0.16773f
C18 rseg_1_v3_1.v42 rseg_1_v3_1.v53 0.02726f
C19 rseg_1_v3_1.v45 rseg_1_v3_1.v41 0.08427f
C20 DEC[1] rseg_1_v3_1.v24 0.20487f
C21 rseg_1_v3_1.v27 rseg_1_v3_1.v30 0.0119f
C22 DEC[0] rseg_1_v3_1.v10 0.17828f
C23 rseg_1_v3_1.v7 rseg_1_v3_1.v4 0.05585f
C24 bb[0] b[1] 0.04277f
C25 rseg_1_v3_1.v36 DEC[2] 0.03176f
C26 rseg_1_v3_1.v55 DEC[3] 0.15096f
C27 rseg_1_v3_1.v39 DEC[2] 0.15051f
C28 DEC[1] rseg_1_v3_1.v29 0.17836f
C29 rseg_1_v3_1.v40 rseg_1_v3_1.v34 0.0119f
C30 rseg_1_v3_1.v40 rseg_1_v3_1.v38 1.73225f
C31 rseg_1_v3_1.v56 rseg_1_v3_1.v54 1.73519f
C32 rseg_1_v3_1.v11 DEC[0] 0.09117f
C33 rseg_1_v3_1.v52 rseg_1_v3_1.v55 0.06115f
C34 rseg_1_v3_1.v11 rseg_1_v3_1.v10 1.27692f
C35 rseg_1_v3_1.v37 DEC[2] 0.06044f
C36 rseg_1_v3_1.v50 DEC[3] 0.06054f
C37 rseg_1_v3_1.v42 rseg_1_v3_1.v45 0.09544f
C38 rseg_1_v3_1.v24 rseg_1_v3_1.v22 1.73509f
C39 rseg_1_v3_1.v61 DEC[3] 0.17877f
C40 rseg_1_v3_1.v42 DEC[3] 0.01149f
C41 b[1] bb[1] 0.04277f
C42 rseg_1_v3_1.v50 rseg_1_v3_1.v52 1.21429f
C43 rseg_1_v3_1.v22 rseg_1_v3_1.v29 0.02015f
C44 rseg_1_v3_1.v39 rseg_1_v3_1.v30 0.01647f
C45 DEC[1] rseg_1_v3_1.v10 0.01136f
C46 DEC[1] rseg_1_v3_1.v25 0.15742f
C47 rseg_1_v3_1.v52 rseg_1_v3_1.v61 0.02197f
C48 rseg_1_v3_1.v36 rseg_1_v3_1.v45 0.02194f
C49 rseg_1_v3_1.v46 rseg_1_v3_1.v43 0.0119f
C50 rseg_1_v3_1.v59 DEC[3] 0.09927f
C51 rseg_1_v3_1.v27 rseg_1_v3_1.v20 0.02198f
C52 rseg_1_v3_1.v30 rseg_1_v3_1.v29 1.19856f
C53 rseg_1_v3_1.v13 rseg_1_v3_1.v6 0.02015f
C54 rseg_1_v3_1.v3 rseg_1_v3_1.v7 0.05245f
C55 rseg_1_v3_1.v44 DEC[2] 0.09138f
C56 rseg_1_v3_1.v40 rseg_1_v3_1.v41 3.81788f
C57 rseg_1_v3_1.v40 rseg_1_v3_1.v55 0.0484f
C58 rseg_1_v3_1.v58 DEC[3] 0.17913f
C59 rseg_1_v3_1.v52 rseg_1_v3_1.v59 0.02201f
C60 rseg_1_v3_1.v25 rseg_1_v3_1.v22 0.04732f
C61 rseg_1_v3_1.v44 rseg_1_v3_1.v53 0.02615f
C62 rseg_1_v3_1.v53 rseg_1_v3_1.v54 0.48841f
C63 rseg_1_v3_1.v46 rseg_1_v3_1.v51 0.02493f
C64 rseg_1_v3_1.v27 rseg_1_v3_1.v26 1.31057f
C65 DEC[0] rseg_1_v3_1.v8 0.15248f
C66 rseg_1_v3_1.v62 DEC[3] 0.15788f
C67 rseg_1_v3_1.v42 rseg_1_v3_1.v40 0.55369f
C68 rseg_1_v3_1.v8 rseg_1_v3_1.v10 0.54398f
C69 rseg_1_v3_1.v60 DEC[3] 0.09325f
C70 rseg_1_v3_1.v38 rseg_1_v3_1.v43 0.05318f
C71 rseg_1_v3_1.v56 DEC[3] 0.29328f
C72 rseg_1_v3_1.v44 rseg_1_v3_1.v45 1.21986f
C73 V0 rseg_1_v3_1.v5 0.22753f
C74 V0 rseg_1_v3_1.v2 1.17753f
C75 DEC[1] rseg_1_v3_1.v22 0.12529f
C76 rseg_1_v3_1.v11 rseg_1_v3_1.v8 0.0981f
C77 DEC[0] rseg_1_v3_1.v12 0.09116f
C78 rseg_1_v3_1.v6 rseg_1_v3_1.v5 0.39192f
C79 rseg_1_v3_1.v20 rseg_1_v3_1.v29 0.02197f
C80 rseg_1_v3_1.v10 rseg_1_v3_1.v12 2.0142f
C81 rseg_1_v3_1.v40 rseg_1_v3_1.v39 0.14454f
C82 rseg_1_v3_1.v18 rseg_1_v3_1.v23 0.05838f
C83 rseg_1_v3_1.v54 DEC[3] 0.097f
C84 rseg_1_v3_1.v39 rseg_1_v3_1.v26 1.34056f
C85 DEC[0] rseg_1_v3_1.v7 0.1499f
C86 rseg_1_v3_1.v35 rseg_1_v3_1.v28 0.03392f
C87 rseg_1_v3_1.v11 rseg_1_v3_1.v12 1.2875f
C88 DEC[1] rseg_1_v3_1.v30 0.15598f
C89 rseg_1_v3_1.v24 rseg_1_v3_1.v26 0.55643f
C90 rseg_1_v3_1.v52 rseg_1_v3_1.v54 1.63811f
C91 rseg_1_v3_1.v26 rseg_1_v3_1.v37 0.02766f
C92 DEC[1] rseg_1_v3_1.v19 0.03135f
C93 rseg_1_v3_1.v26 rseg_1_v3_1.v29 0.0954f
C94 DEC[0] rseg_1_v3_1.v14 0.15587f
C95 rseg_1_v3_1.v10 rseg_1_v3_1.v14 0.43907f
C96 rseg_1_v3_1.v30 DEC[2] 0.02106f
C97 rseg_1_v3_1.v43 rseg_1_v3_1.v41 1.7882f
C98 rseg_1_v3_1.v45 DEC[2] 0.17841f
C99 rseg_1_v3_1.v11 rseg_1_v3_1.v14 0.0119f
C100 rseg_1_v3_1.v13 rseg_1_v3_1.v2 0.01887f
C101 rseg_1_v3_1.v9 rseg_1_v3_1.v6 0.04313f
C102 rseg_1_v3_1.v34 rseg_1_v3_1.v35 0.66352f
C103 DEC[3] DEC[2] 0.01053f
C104 V0 rseg_1_v3_1.v4 0.01904f
C105 rseg_1_v3_1.v6 rseg_1_v3_1.v4 1.8445f
C106 rseg_1_v3_1.v53 DEC[3] 0.06038f
C107 rseg_1_v3_1.v25 rseg_1_v3_1.v26 1.29067f
C108 rseg_1_v3_1.v21 rseg_1_v3_1.v10 0.02839f
C109 DEC[1] rseg_1_v3_1.v14 0.02042f
C110 DEC[1] rseg_1_v3_1.v20 0.03142f
C111 rseg_1_v3_1.v42 rseg_1_v3_1.v43 1.34308f
C112 rseg_1_v3_1.v52 rseg_1_v3_1.v53 0.60003f
C113 rseg_1_v3_1.v55 rseg_1_v3_1.v51 0.05244f
C114 bb[0] VOUT 0.10609f
C115 rseg_1_v3_1.v50 rseg_1_v3_1.v51 0.69962f
C116 rseg_1_v3_1.v43 rseg_1_v3_1.v36 0.02214f
C117 rseg_1_v3_1.v19 rseg_1_v3_1.v12 0.03446f
C118 rseg_1_v3_1.v13 rseg_1_v3_1.v9 0.08427f
C119 DEC[1] rseg_1_v3_1.v26 0.17853f
C120 rseg_1_v3_1.v5 rseg_1_v3_1.v2 0.0481f
C121 rseg_1_v3_1.v22 rseg_1_v3_1.v20 1.68068f
C122 rseg_1_v3_1.v8 rseg_1_v3_1.v7 0.04824f
C123 DEC[1] rseg_1_v3_1.v21 0.06044f
C124 rseg_1_v3_1.v13 rseg_1_v3_1.v4 0.01848f
C125 V0 rseg_1_v3_1.v3 0.32489f
C126 rseg_1_v3_1.v52 DEC[3] 0.03202f
C127 rseg_1_v3_1.v40 DEC[2] 0.258f
C128 rseg_1_v3_1.v26 DEC[2] 0.01144f
C129 rseg_1_v3_1.v19 rseg_1_v3_1.v14 0.02541f
C130 rseg_1_v3_1.v20 rseg_1_v3_1.v19 0.54711f
C131 rseg_1_v3_1.v21 rseg_1_v3_1.v22 0.42912f
C132 rseg_1_v3_1.v12 rseg_1_v3_1.v14 1.15763f
C133 V64 rseg_1_v3_1.v58 0.16537f
C134 rseg_1_v3_1.v46 rseg_1_v3_1.v55 0.01649f
C135 rseg_1_v3_1.v26 rseg_1_v3_1.v30 0.36625f
C136 rseg_1_v3_1.v44 rseg_1_v3_1.v43 1.34563f
C137 rseg_1_v3_1.v24 rseg_1_v3_1.v23 0.10072f
C138 rseg_1_v3_1.v40 rseg_1_v3_1.v45 0.21426f
C139 rseg_1_v3_1.v4 rseg_1_v3_1.v5 0.50407f
C140 rseg_1_v3_1.v4 rseg_1_v3_1.v2 1.40088f
C141 rseg_1_v3_1.v35 rseg_1_v3_1.v36 0.57986f
C142 rseg_1_v3_1.v39 rseg_1_v3_1.v35 0.05244f
C143 b[2] bb[2] 0.04353f
C144 rseg_1_v3_1.v21 rseg_1_v3_1.v19 1.44458f
C145 rseg_1_v3_1.v27 rseg_1_v3_1.v28 1.31906f
C146 V0 DEC[0] 0.05996f
C147 V64 rseg_1_v3_1.v62 0.76724f
C148 rseg_1_v3_1.v46 rseg_1_v3_1.v42 0.33336f
C149 V64 rseg_1_v3_1.v60 0.18355f
C150 rseg_1_v3_1.v35 rseg_1_v3_1.v37 1.45085f
C151 DEC[0] rseg_1_v3_1.v6 0.11835f
C152 rseg_1_v3_1.v21 rseg_1_v3_1.v12 0.0266f
C153 rseg_1_v3_1.v44 rseg_1_v3_1.v51 0.03397f
C154 rseg_1_v3_1.v11 rseg_1_v3_1.v6 0.04904f
C155 rseg_1_v3_1.v38 rseg_1_v3_1.v41 0.04748f
C156 rseg_1_v3_1.v10 rseg_1_v3_1.v23 1.34685f
C157 rseg_1_v3_1.v43 DEC[2] 0.0945f
C158 rseg_1_v3_1.v21 rseg_1_v3_1.v20 0.54188f
C159 rseg_1_v3_1.v3 rseg_1_v3_1.v5 1.41253f
C160 rseg_1_v3_1.v3 rseg_1_v3_1.v2 0.59845f
C161 rseg_1_v3_1.v37 rseg_1_v3_1.v28 0.02611f
C162 rseg_1_v3_1.v29 rseg_1_v3_1.v28 1.19056f
C163 rseg_1_v3_1.v13 DEC[0] 0.17825f
C164 rseg_1_v3_1.v24 rseg_1_v3_1.v18 0.0119f
C165 rseg_1_v3_1.v13 rseg_1_v3_1.v10 0.09535f
C166 DEC[1] rseg_1_v3_1.v23 0.15222f
C167 rseg_1_v3_1.v18 rseg_1_v3_1.v29 0.02163f
C168 rseg_1_v3_1.v13 rseg_1_v3_1.v11 1.72759f
C169 rseg_1_v3_1.v34 rseg_1_v3_1.v36 1.22987f
C170 rseg_1_v3_1.v38 rseg_1_v3_1.v36 1.64648f
C171 rseg_1_v3_1.v39 rseg_1_v3_1.v34 0.05777f
C172 rseg_1_v3_1.v39 rseg_1_v3_1.v38 0.62948f
C173 rseg_1_v3_1.v53 rseg_1_v3_1.v51 1.45197f
C174 rseg_1_v3_1.v43 rseg_1_v3_1.v45 1.73307f
C175 rseg_1_v3_1.v46 rseg_1_v3_1.v44 1.15703f
C176 rseg_1_v3_1.v25 rseg_1_v3_1.v28 0.02715f
C177 rseg_1_v3_1.v34 rseg_1_v3_1.v37 0.04811f
C178 rseg_1_v3_1.v37 rseg_1_v3_1.v38 0.4572f
C179 rseg_1_v3_1.v22 rseg_1_v3_1.v23 0.59336f
C180 rseg_1_v3_1.v57 rseg_1_v3_1.v61 0.08493f
C181 rseg_1_v3_1.v35 DEC[2] 0.03135f
C182 rseg_1_v3_1.v6 rseg_1_v3_1.v8 1.73087f
C183 rseg_1_v3_1.v50 rseg_1_v3_1.v55 0.05769f
C184 b[0] VOUT 0.16526f
C185 rseg_1_v3_1.v3 rseg_1_v3_1.v4 0.51079f
C186 DEC[0] rseg_1_v3_1.v5 0.06052f
C187 DEC[0] rseg_1_v3_1.v2 0.06158f
C188 rseg_1_v3_1.v42 rseg_1_v3_1.v41 1.32022f
C189 rseg_1_v3_1.v42 rseg_1_v3_1.v55 1.33973f
C190 rseg_1_v3_1.v51 DEC[3] 0.03135f
C191 rseg_1_v3_1.v8 rseg_1_v3_1.v23 0.05173f
C192 rseg_1_v3_1.v57 rseg_1_v3_1.v59 1.79255f
C193 rseg_1_v3_1.v23 rseg_1_v3_1.v19 0.05244f
C194 V0 rseg_1_v3_1.v7 0.27768f
C195 DEC[1] rseg_1_v3_1.v28 0.09131f
C196 rseg_1_v3_1.v52 rseg_1_v3_1.v51 0.60342f
C197 rseg_1_v3_1.v50 rseg_1_v3_1.v61 0.02147f
C198 rseg_1_v3_1.v6 rseg_1_v3_1.v7 0.55841f
C199 rseg_1_v3_1.v58 rseg_1_v3_1.v57 1.34945f
C200 rseg_1_v3_1.v35 rseg_1_v3_1.v30 0.02537f
C201 DEC[1] rseg_1_v3_1.v18 0.06065f
C202 rseg_1_v3_1.v46 DEC[2] 0.15602f
C203 rseg_1_v3_1.v40 rseg_1_v3_1.v43 0.09811f
C204 rseg_1_v3_1.v13 rseg_1_v3_1.v8 0.2143f
C205 rseg_1_v3_1.v27 rseg_1_v3_1.v24 0.09809f
C206 rseg_1_v3_1.v9 DEC[0] 0.15598f
C207 rseg_1_v3_1.v59 rseg_1_v3_1.v61 1.73155f
C208 rseg_1_v3_1.v9 rseg_1_v3_1.v10 1.25806f
C209 rseg_1_v3_1.v57 rseg_1_v3_1.v60 0.02715f
C210 bb[0] b[0] 0.04277f
C211 rseg_1_v3_1.v27 rseg_1_v3_1.v29 1.72824f
C212 DEC[0] rseg_1_v3_1.v4 0.03958f
C213 rseg_1_v3_1.v13 rseg_1_v3_1.v12 1.15809f
C214 rseg_1_v3_1.v56 rseg_1_v3_1.v57 3.83937f
C215 rseg_1_v3_1.v23 rseg_1_v3_1.v14 0.01643f
C216 rseg_1_v3_1.v20 rseg_1_v3_1.v23 0.06177f
C217 rseg_1_v3_1.v58 rseg_1_v3_1.v61 0.0961f
C218 rseg_1_v3_1.v30 rseg_1_v3_1.v28 1.1572f
C219 rseg_1_v3_1.v9 rseg_1_v3_1.v11 1.78725f
C220 rseg_1_v3_1.v46 rseg_1_v3_1.v45 1.22792f
C221 rseg_1_v3_1.v39 rseg_1_v3_1.v36 0.06132f
C222 rseg_1_v3_1.v56 rseg_1_v3_1.v55 0.17104f
C223 rseg_1_v3_1.v11 rseg_1_v3_1.v4 0.01835f
C224 rseg_1_v3_1.v57 rseg_1_v3_1.v54 0.04735f
C225 rseg_1_v3_1.v34 DEC[2] 0.06082f
C226 rseg_1_v3_1.v38 DEC[2] 0.09798f
C227 rseg_1_v3_1.v46 DEC[3] 0.02161f
C228 rseg_1_v3_1.v44 rseg_1_v3_1.v41 0.02715f
C229 rseg_1_v3_1.v39 rseg_1_v3_1.v24 0.04787f
C230 rseg_1_v3_1.v18 rseg_1_v3_1.v19 0.63647f
C231 rseg_1_v3_1.v58 rseg_1_v3_1.v59 1.36638f
C232 rseg_1_v3_1.v37 rseg_1_v3_1.v36 0.57403f
C233 rseg_1_v3_1.v39 rseg_1_v3_1.v37 1.97694f
C234 rseg_1_v3_1.v62 rseg_1_v3_1.v61 1.25122f
C235 rseg_1_v3_1.v54 rseg_1_v3_1.v55 0.65418f
C236 bb[1] bb[2] 0.04353f
C237 rseg_1_v3_1.v50 rseg_1_v3_1.v56 0.0119f
C238 rseg_1_v3_1.v13 rseg_1_v3_1.v14 1.16723f
C239 rseg_1_v3_1.v27 rseg_1_v3_1.v25 1.789f
C240 rseg_1_v3_1.v8 rseg_1_v3_1.v2 0.0119f
C241 rseg_1_v3_1.v61 rseg_1_v3_1.v60 1.24381f
C242 rseg_1_v3_1.v21 rseg_1_v3_1.v23 1.97444f
C243 rseg_1_v3_1.v56 rseg_1_v3_1.v61 0.21492f
C244 rseg_1_v3_1.v24 rseg_1_v3_1.v29 0.21425f
C245 rseg_1_v3_1.v42 rseg_1_v3_1.v44 1.916f
C246 rseg_1_v3_1.v59 rseg_1_v3_1.v62 0.0119f
C247 rseg_1_v3_1.v3 DEC[0] 0.03915f
C248 rseg_1_v3_1.v54 rseg_1_v3_1.v61 0.02015f
C249 rseg_1_v3_1.v34 rseg_1_v3_1.v45 0.02179f
C250 rseg_1_v3_1.v38 rseg_1_v3_1.v45 0.02015f
C251 rseg_1_v3_1.v59 rseg_1_v3_1.v60 1.37492f
C252 rseg_1_v3_1.v7 rseg_1_v3_1.v5 1.9603f
C253 rseg_1_v3_1.v7 rseg_1_v3_1.v2 0.0555f
C254 rseg_1_v3_1.v56 rseg_1_v3_1.v59 0.09809f
C255 rseg_1_v3_1.v58 rseg_1_v3_1.v62 0.31595f
C256 V64 GND 0.73424f
C257 V0 GND 1.62173f
C258 DEC[3] GND 5.17399f
C259 DEC[2] GND 4.78008f
C260 DEC[1] GND 4.92723f
C261 DEC[0] GND 5.51685f
C262 b[3] GND 2.3967f
C263 bb[3] GND 2.33896f
C264 VOUT GND 0.34261f
C265 b[2] GND 1.18209f
C266 bb[2] GND 1.14271f
C267 bb[1] GND 0.55895f
C268 b[1] GND 0.5536f
C269 bb[0] GND 0.28631f
C270 b[0] GND 0.31391f
C271 rseg_1_v3_1.v55 GND 1.58528f
C272 rseg_1_v3_1.v54 GND 1.01698f
C273 rseg_1_v3_1.v53 GND 0.83396f
C274 rseg_1_v3_1.v52 GND 0.84338f
C275 rseg_1_v3_1.v51 GND 0.72928f
C276 rseg_1_v3_1.v50 GND 0.81839f
C277 rseg_1_v3_1.v39 GND 1.60778f
C278 rseg_1_v3_1.v38 GND 1.05072f
C279 rseg_1_v3_1.v37 GND 0.85279f
C280 rseg_1_v3_1.v36 GND 0.85992f
C281 rseg_1_v3_1.v35 GND 0.74171f
C282 rseg_1_v3_1.v34 GND 0.83636f
C283 rseg_1_v3_1.v23 GND 1.64324f
C284 rseg_1_v3_1.v22 GND 1.10435f
C285 rseg_1_v3_1.v21 GND 0.88408f
C286 rseg_1_v3_1.v20 GND 0.90291f
C287 rseg_1_v3_1.v19 GND 0.77336f
C288 rseg_1_v3_1.v18 GND 0.88264f
C289 rseg_1_v3_1.v7 GND 2.55779f
C290 rseg_1_v3_1.v6 GND 1.42715f
C291 rseg_1_v3_1.v5 GND 1.11483f
C292 rseg_1_v3_1.v4 GND 1.14591f
C293 rseg_1_v3_1.v3 GND 1.00561f
C294 rseg_1_v3_1.v2 GND 1.11031f
C295 rseg_1_v3_1.v62 GND 1.01582f
C296 rseg_1_v3_1.v61 GND 0.9432f
C297 rseg_1_v3_1.v60 GND 0.93065f
C298 rseg_1_v3_1.v59 GND 0.86196f
C299 rseg_1_v3_1.v58 GND 1.65047f
C300 rseg_1_v3_1.v57 GND 2.41521f
C301 rseg_1_v3_1.v56 GND 3.42807f
C302 rseg_1_v3_1.v46 GND 0.999f
C303 rseg_1_v3_1.v45 GND 0.9622f
C304 rseg_1_v3_1.v44 GND 0.95203f
C305 rseg_1_v3_1.v43 GND 0.93445f
C306 rseg_1_v3_1.v42 GND 1.12363f
C307 rseg_1_v3_1.v41 GND 2.48425f
C308 rseg_1_v3_1.v40 GND 3.47892f
C309 rseg_1_v3_1.v30 GND 1.03387f
C310 rseg_1_v3_1.v29 GND 0.98141f
C311 rseg_1_v3_1.v28 GND 0.97038f
C312 rseg_1_v3_1.v27 GND 0.95434f
C313 rseg_1_v3_1.v26 GND 1.13851f
C314 rseg_1_v3_1.v25 GND 2.48829f
C315 rseg_1_v3_1.v24 GND 3.56548f
C316 rseg_1_v3_1.v14 GND 1.10656f
C317 rseg_1_v3_1.v13 GND 1.03923f
C318 rseg_1_v3_1.v12 GND 1.49966f
C319 rseg_1_v3_1.v11 GND 1.01681f
C320 rseg_1_v3_1.v10 GND 1.69216f
C321 rseg_1_v3_1.v9 GND 2.57353f
C322 rseg_1_v3_1.v8 GND 3.90298f
C323 a_6627_6728.t1 GND 0.10211f
C324 a_6627_6728.t2 GND 0.12012f
C325 a_6627_6728.n0 GND 5.90174f
C326 a_6627_6728.t0 GND 0.07604f
C327 a_6745_6728.t2 GND 0.12718f
C328 a_6745_6728.t1 GND 0.07284f
C329 a_6745_6728.n0 GND 6.19294f
C330 a_6745_6728.t0 GND 0.10705f
C331 a_7021_6728.t2 GND 0.12828f
C332 a_7021_6728.t1 GND 0.06882f
C333 a_7021_6728.n0 GND 6.09613f
C334 a_7021_6728.t0 GND 0.10677f
C335 a_3759_5464.t1 GND 0.10563f
C336 a_3759_5464.t3 GND 0.08474f
C337 a_3759_5464.n0 GND 3.77304f
C338 a_3759_5464.t2 GND 0.08064f
C339 a_3759_5464.n1 GND 2.70857f
C340 a_3759_5464.t4 GND 0.14779f
C341 a_3759_5464.n2 GND 5.91896f
C342 a_3759_5464.t0 GND 0.08064f
C343 rseg_1_v3_1.v56.t0 GND 0.03703f
C344 rseg_1_v3_1.v56.t2 GND 0.12366f
C345 rseg_1_v3_1.v56.t1 GND 0.36626f
C346 rseg_1_v3_1.v56.n0 GND 2.56502f
C347 a_7297_6728.t2 GND 0.13049f
C348 a_7297_6728.t1 GND 0.06644f
C349 a_7297_6728.n0 GND 6.09434f
C350 a_7297_6728.t0 GND 0.10872f
C351 rseg_1_v3_1.v41.t0 GND 0.04657f
C352 rseg_1_v3_1.v41.t1 GND 0.13984f
C353 rseg_1_v3_1.v41.t2 GND 0.13973f
C354 rseg_1_v3_1.v41.n0 GND 2.57846f
C355 rseg_1_v3_1.v25.t0 GND 0.04645f
C356 rseg_1_v3_1.v25.t2 GND 0.13937f
C357 rseg_1_v3_1.v25.t1 GND 0.14921f
C358 rseg_1_v3_1.v25.n0 GND 2.57872f
C359 a_2221_5464.t1 GND 0.04115f
C360 a_2221_5464.t3 GND 0.05703f
C361 a_2221_5464.n0 GND 1.94212f
C362 a_2221_5464.t2 GND 0.03868f
C363 a_2221_5464.n1 GND 1.52384f
C364 a_2221_5464.t4 GND 0.06894f
C365 a_2221_5464.n2 GND 2.78956f
C366 a_2221_5464.t0 GND 0.03868f
C367 a_613_4028.t1 GND 0.12364f
C368 a_613_4028.t2 GND 0.07206f
C369 a_613_4028.n0 GND 4.94854f
C370 a_613_4028.t4 GND 0.15859f
C371 a_613_4028.n1 GND 4.24803f
C372 a_613_4028.t3 GND 0.15202f
C373 a_613_4028.n2 GND 4.62506f
C374 a_613_4028.t0 GND 0.07206f
C375 rseg_1_v3_1.v24.t0 GND 0.03636f
C376 rseg_1_v3_1.v24.t1 GND 0.12209f
C377 rseg_1_v3_1.v24.t2 GND 0.36895f
C378 rseg_1_v3_1.v24.n0 GND 2.57743f
C379 a_4311_5464.t1 GND 0.05828f
C380 a_4311_5464.t3 GND 0.04276f
C381 a_4311_5464.n0 GND 2.03892f
C382 a_4311_5464.t2 GND 0.04087f
C383 a_4311_5464.n1 GND 1.29976f
C384 a_4311_5464.t4 GND 0.07543f
C385 a_4311_5464.n2 GND 3.00311f
C386 a_4311_5464.t0 GND 0.04087f
C387 a_1047_4028.t3 GND 0.15386f
C388 a_1047_4028.t2 GND 0.07275f
C389 a_1047_4028.n0 GND 5.76483f
C390 a_1047_4028.t4 GND 0.15297f
C391 a_1047_4028.n1 GND 4.11942f
C392 a_1047_4028.t1 GND 0.07275f
C393 a_1047_4028.n2 GND 3.93804f
C394 a_1047_4028.t0 GND 0.12539f
C395 a_61_4028.t3 GND 0.17054f
C396 a_61_4028.t1 GND 0.0814f
C397 a_61_4028.n0 GND 5.33946f
C398 a_61_4028.t4 GND 0.17912f
C399 a_61_4028.n1 GND 4.85263f
C400 a_61_4028.t2 GND 0.0814f
C401 a_61_4028.n2 GND 5.35733f
C402 a_61_4028.t0 GND 0.13813f
C403 rseg_1_v3_1.v57.t0 GND 0.04652f
C404 rseg_1_v3_1.v57.t2 GND 0.13968f
C405 rseg_1_v3_1.v57.t1 GND 0.13957f
C406 rseg_1_v3_1.v57.n0 GND 2.57959f
C407 a_6351_6728.t2 GND 0.11093f
C408 a_6351_6728.t1 GND 0.07357f
C409 a_6351_6728.n0 GND 5.52202f
C410 a_6351_6728.t0 GND 0.09348f
C411 rseg_1_v3_1.v9.t2 GND 0.04754f
C412 rseg_1_v3_1.v9.t0 GND 0.14298f
C413 rseg_1_v3_1.v9.t1 GND 0.14263f
C414 rseg_1_v3_1.v9.n0 GND 2.55569f
C415 a_2497_5464.t1 GND 0.0855f
C416 a_2497_5464.t3 GND 0.14007f
C417 a_2497_5464.t4 GND 0.07805f
C418 a_2497_5464.n0 GND 5.65951f
C419 a_2497_5464.t2 GND 0.07805f
C420 a_2497_5464.n1 GND 2.99489f
C421 a_2497_5464.n2 GND 3.75935f
C422 a_2497_5464.t0 GND 0.10458f
C423 rseg_1_v3_1.v8.t2 GND 0.0341f
C424 rseg_1_v3_1.v8.t1 GND 0.12376f
C425 rseg_1_v3_1.v8.t0 GND 0.363f
C426 rseg_1_v3_1.v8.n0 GND 2.62718f
C427 a_6075_6728.t2 GND 0.10894f
C428 a_6075_6728.t1 GND 0.07635f
C429 a_6075_6728.n0 GND 5.52296f
C430 a_6075_6728.t0 GND 0.09175f
C431 a_4035_5464.t4 GND 0.14987f
C432 a_4035_5464.t1 GND 0.08147f
C433 a_4035_5464.n0 GND 5.98504f
C434 a_4035_5464.t3 GND 0.08147f
C435 a_4035_5464.n1 GND 2.66272f
C436 a_4035_5464.t2 GND 0.08541f
C437 a_4035_5464.n2 GND 3.94271f
C438 a_4035_5464.t0 GND 0.11133f
C439 rseg_1_v3_1.v40.t1 GND 0.03678f
C440 rseg_1_v3_1.v40.t0 GND 0.12308f
C441 rseg_1_v3_1.v40.t2 GND 0.36729f
C442 rseg_1_v3_1.v40.n0 GND 2.56969f
C443 a_7573_6728.t2 GND 0.06636f
C444 a_7573_6728.t1 GND 0.03208f
C445 a_7573_6728.n0 GND 3.04622f
C446 a_7573_6728.t0 GND 0.05535f
C447 a_1599_4028.t1 GND 0.14531f
C448 a_1599_4028.t2 GND 0.08367f
C449 a_1599_4028.n0 GND 4.77562f
C450 a_1599_4028.t4 GND 0.14572f
C451 a_1599_4028.n1 GND 4.0453f
C452 a_1599_4028.t3 GND 0.17762f
C453 a_1599_4028.n2 GND 6.44309f
C454 a_1599_4028.t0 GND 0.08367f
C455 rseg_1_v3_1.v12.t2 GND 0.02587f
C456 rseg_1_v3_1.v12.t0 GND 0.07998f
C457 rseg_1_v3_1.v12.t1 GND 0.07984f
C458 rseg_1_v3_1.v12.n0 GND 1.3573f
C459 a_3483_5464.t4 GND 0.10032f
C460 a_3483_5464.t3 GND 0.08434f
C461 a_3483_5464.n0 GND 3.60497f
C462 a_3483_5464.t1 GND 0.07983f
C463 a_3483_5464.n1 GND 2.75522f
C464 a_3483_5464.t2 GND 0.14569f
C465 a_3483_5464.n2 GND 5.84981f
C466 a_3483_5464.t0 GND 0.07983f
C467 a_2773_5464.t1 GND 0.0892f
C468 a_2773_5464.t4 GND 0.14222f
C469 a_2773_5464.t2 GND 0.07875f
C470 a_2773_5464.n0 GND 5.73614f
C471 a_2773_5464.t3 GND 0.07875f
C472 a_2773_5464.n1 GND 2.9429f
C473 a_2773_5464.n2 GND 3.63616f
C474 a_2773_5464.t0 GND 0.09588f
C475 a_5799_6728.t1 GND 0.04502f
C476 a_5799_6728.t2 GND 0.05347f
C477 a_5799_6728.n0 GND 2.76188f
C478 a_5799_6728.t0 GND 0.03963f
C479 a_n215_4028.t4 GND 0.06897f
C480 a_n215_4028.t1 GND 0.04091f
C481 a_n215_4028.n0 GND 2.62657f
C482 a_n215_4028.t3 GND 0.08929f
C483 a_n215_4028.n1 GND 2.43648f
C484 a_n215_4028.t2 GND 0.08534f
C485 a_n215_4028.n2 GND 2.71152f
C486 a_n215_4028.t0 GND 0.04091f
C487 a_1323_4028.t2 GND 0.14276f
C488 a_1323_4028.t3 GND 0.08249f
C489 a_1323_4028.n0 GND 4.59159f
C490 a_1323_4028.t1 GND 0.15799f
C491 a_1323_4028.n1 GND 4.32313f
C492 a_1323_4028.t4 GND 0.17484f
C493 a_1323_4028.n2 GND 6.44471f
C494 a_1323_4028.t0 GND 0.08249f
C495 a_3049_5464.t4 GND 0.14424f
C496 a_3049_5464.t3 GND 0.07942f
C497 a_3049_5464.n0 GND 5.80531f
C498 a_3049_5464.t2 GND 0.07942f
C499 a_3049_5464.n1 GND 2.88984f
C500 a_3049_5464.t1 GND 0.08812f
C501 a_3049_5464.n2 GND 3.52034f
C502 a_3049_5464.t0 GND 0.0933f
C503 a_337_4028.t1 GND 0.13945f
C504 a_337_4028.t2 GND 0.0817f
C505 a_337_4028.n0 GND 5.49877f
C506 a_337_4028.t4 GND 0.17181f
C507 a_337_4028.t3 GND 0.0817f
C508 a_337_4028.n1 GND 5.30212f
C509 a_337_4028.n2 GND 4.84462f
C510 a_337_4028.t0 GND 0.17983f
C511 rseg_1_v3_1.v10.t1 GND 0.02638f
C512 rseg_1_v3_1.v10.t2 GND 0.07391f
C513 rseg_1_v3_1.v10.t0 GND 0.0738f
C514 rseg_1_v3_1.v10.n0 GND 1.32117f
C515 a_1875_4028.t4 GND 0.09262f
C516 a_1875_4028.t3 GND 0.04358f
C517 a_1875_4028.n0 GND 3.30724f
C518 a_1875_4028.t2 GND 0.06837f
C519 a_1875_4028.n1 GND 1.92423f
C520 a_1875_4028.t1 GND 0.04358f
C521 a_1875_4028.n2 GND 2.54446f
C522 a_1875_4028.t0 GND 0.07592f
.ends

