magic
tech sky130A
magscale 1 2
timestamp 1751017459
<< metal1 >>
rect 8731 3155 8791 3161
rect 8731 1519 8791 3095
rect 101 1327 161 1453
rect 101 789 161 1267
rect 1829 1239 1889 1453
rect 1829 789 1889 1179
rect 3557 1151 3617 1453
rect 3557 789 3617 1091
rect 5285 1063 5345 1453
rect 5285 789 5345 1003
rect 7013 975 7073 1453
rect 7013 789 7073 915
rect 8731 695 8791 1459
rect 8731 -125 8791 635
rect 8731 -191 8791 -185
<< via1 >>
rect 8731 3095 8791 3155
rect 8731 1459 8791 1519
rect 101 1267 161 1327
rect 1829 1179 1889 1239
rect 3557 1091 3617 1151
rect 5285 1003 5345 1063
rect 7013 915 7073 975
rect 8731 635 8791 695
rect 8731 -185 8791 -125
<< metal2 >>
rect 8703 3095 8731 3155
rect 8791 3095 8797 3155
rect 8703 1459 8731 1519
rect 8791 1459 8797 1519
rect 95 1267 101 1327
rect 161 1267 7079 1327
rect 95 1179 1829 1239
rect 1889 1179 7079 1239
rect 95 1091 3557 1151
rect 3617 1091 7079 1151
rect 95 1003 5285 1063
rect 5345 1003 7079 1063
rect 95 915 7013 975
rect 7073 915 7079 975
rect 8703 635 8731 695
rect 8791 635 8797 695
rect 8703 -185 8731 -125
rect 8791 -185 8797 -125
use dp_nmos_top  dp_nmos_top_0
timestamp 1750150351
transform 1 0 -18 0 1 -321
box -15 -4 8757 1244
use dp_pmos_top  dp_pmos_top_0
timestamp 1750150351
transform 1 0 -53 0 1 1304
box -10 -15 8822 2109
<< end >>
