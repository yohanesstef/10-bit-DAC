magic
tech sky130A
magscale 1 2
timestamp 1749479165
<< pwell >>
rect -150 -174 682 364
<< mvpsubdiff >>
rect -114 270 646 328
rect -114 220 -56 270
rect -114 -30 -102 220
rect -68 -30 -56 220
rect -114 -80 -56 -30
rect 588 220 646 270
rect 588 -30 600 220
rect 634 -30 646 220
rect 588 -80 646 -30
rect -114 -138 646 -80
<< mvpsubdiffcont >>
rect -102 -30 -68 220
rect 600 -30 634 220
<< locali >>
rect -102 282 634 316
rect -102 220 -68 282
rect -102 -92 -68 -30
rect 600 220 634 282
rect 600 -92 634 -30
rect -102 -126 634 -92
<< metal1 >>
rect 18 36 46 208
rect 189 -88 217 84
rect 300 45 328 217
rect 470 -103 498 69
use hnmos_2  hnmos_2_0
timestamp 1749478216
transform 1 0 -6 0 1 -5
box -4 1 548 199
<< labels >>
flabel metal1 s 18 208 18 208 4 FreeSans 480 0 0 0 vin[0]
port 0 se
flabel metal1 s 300 217 300 217 4 FreeSans 480 0 0 0 vin[1]
port 1 se
flabel metal2 s 256 138 256 138 4 FreeSans 480 0 0 0 DIN
port 2 se
flabel metal1 s 484 -87 484 -87 4 FreeSans 480 0 0 0 VH
port 3 se
flabel metal1 s 201 -60 201 -60 4 FreeSans 480 0 0 0 VL
port 4 se
flabel locali s -93 -108 -93 -108 4 FreeSans 480 0 0 0 VNB
port 5 se
<< end >>
