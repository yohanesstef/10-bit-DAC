magic
tech sky130A
magscale 1 2
timestamp 1750773250
<< mvpsubdiffcont >>
rect 4159 -3193 4205 -3159
<< mvnsubdiffcont >>
rect 4072 645 4180 679
<< viali >>
rect 4072 645 4180 679
rect 4159 -3193 4205 -3159
<< metal1 >>
rect 7127 236 7187 242
rect 7127 170 7187 176
rect 7637 -267 7643 -207
rect 7703 -267 7709 -207
rect 7180 -494 7385 -434
rect 7445 -494 7451 -434
rect 7379 -794 7385 -734
rect 7445 -794 7451 -734
rect 7637 -794 7643 -734
rect 7703 -794 7709 -734
rect 6360 -2178 6370 -2118
rect 6430 -2178 6436 -2118
rect 6360 -2559 6368 -2534
rect 6428 -2559 6436 -2534
rect 6994 -2637 7000 -2577
rect 7060 -2637 7066 -2577
rect 5981 -2932 5989 -2872
rect 6049 -2932 6057 -2872
rect 6988 -3010 6994 -2950
rect 7054 -3010 7060 -2950
rect 3924 -3597 4388 -3216
rect 6982 -3385 6988 -3325
<< via1 >>
rect 7127 176 7187 236
rect 7643 -267 7703 -207
rect 7385 -494 7445 -434
rect 7385 -794 7445 -734
rect 7643 -794 7703 -734
rect 6370 -2178 6430 -2118
rect 6368 -2559 6428 -2499
rect 7000 -2637 7060 -2577
rect 5989 -2932 6049 -2872
rect 6994 -3010 7054 -2950
rect 6988 -3385 7048 -3325
<< metal2 >>
rect 6340 176 7127 236
rect 7187 176 7193 236
rect 5041 -110 5051 -54
rect 5107 -110 5117 -54
rect 5855 -198 5865 -142
rect 5921 -198 5931 -142
rect 7637 -267 7643 -207
rect 7703 -267 7709 -207
rect 6275 -318 6430 -316
rect 6275 -374 6370 -318
rect 6426 -374 6436 -318
rect 6275 -376 6430 -374
rect 5981 -462 5991 -406
rect 6047 -462 6057 -406
rect 7385 -434 7445 -428
rect 7385 -734 7445 -494
rect 7385 -800 7445 -794
rect 7643 -734 7703 -267
rect 7643 -1264 7703 -794
rect 5178 -1324 7703 -1264
rect 5178 -1926 5238 -1324
rect 5860 -1514 5992 -1512
rect 5855 -1570 5865 -1514
rect 5921 -1570 5992 -1514
rect 5860 -1572 5992 -1570
rect 6489 -1961 6499 -1905
rect 6555 -1961 6565 -1905
rect 5041 -2044 5051 -1988
rect 5107 -2044 5117 -1988
rect 5981 -2176 5991 -2120
rect 6047 -2176 6057 -2120
rect 6360 -2178 6370 -2118
rect 6430 -2178 6436 -2118
rect 6804 -2264 6814 -2208
rect 6870 -2264 6880 -2208
rect 6930 -2352 6940 -2296
rect 6996 -2352 7006 -2296
rect 6360 -2559 6368 -2499
rect 6428 -2559 6436 -2499
rect 6489 -2579 7000 -2577
rect 6489 -2635 6499 -2579
rect 6555 -2635 7000 -2579
rect 6489 -2637 7000 -2635
rect 7060 -2637 7066 -2577
rect 5981 -2932 5989 -2872
rect 6049 -2932 6057 -2872
rect 6988 -2952 6994 -2950
rect 6930 -3008 6940 -2952
rect 6988 -3010 6994 -3008
rect 7054 -3010 7060 -2950
rect 6804 -3327 6988 -3325
rect 6804 -3383 6814 -3327
rect 6870 -3383 6988 -3327
rect 6804 -3385 6988 -3383
rect 7048 -3385 7054 -3325
<< via2 >>
rect 5051 -110 5107 -54
rect 5865 -198 5921 -142
rect 6370 -374 6426 -318
rect 5991 -462 6047 -406
rect 5865 -1570 5921 -1514
rect 6499 -1961 6555 -1905
rect 5051 -2044 5107 -1988
rect 5991 -2176 6047 -2120
rect 6370 -2176 6426 -2120
rect 6814 -2264 6870 -2208
rect 6940 -2352 6996 -2296
rect 6370 -2555 6426 -2499
rect 6499 -2635 6555 -2579
rect 5991 -2928 6047 -2872
rect 6940 -3008 6994 -2952
rect 6994 -3008 6996 -2952
rect 6814 -3383 6870 -3327
<< metal3 >>
rect 5046 -54 5112 -44
rect 5046 -110 5051 -54
rect 5107 -110 5112 -54
rect 5046 -1988 5112 -110
rect 5860 -142 5926 -132
rect 5860 -198 5865 -142
rect 5921 -198 5926 -142
rect 5860 -1514 5926 -198
rect 6365 -318 6431 -308
rect 6365 -374 6370 -318
rect 6426 -374 6431 -318
rect 5860 -1570 5865 -1514
rect 5921 -1570 5926 -1514
rect 5860 -1580 5926 -1570
rect 5986 -406 6052 -396
rect 5986 -462 5991 -406
rect 6047 -462 6052 -406
rect 5046 -2044 5051 -1988
rect 5107 -2044 5112 -1988
rect 5046 -2054 5112 -2044
rect 5986 -2120 6052 -462
rect 5986 -2176 5991 -2120
rect 6047 -2176 6052 -2120
rect 5986 -2872 6052 -2176
rect 6365 -2120 6431 -374
rect 6365 -2176 6370 -2120
rect 6426 -2176 6431 -2120
rect 6365 -2499 6431 -2176
rect 6365 -2555 6370 -2499
rect 6426 -2555 6431 -2499
rect 6365 -2565 6431 -2555
rect 6494 -1905 6560 -1895
rect 6494 -1961 6499 -1905
rect 6555 -1961 6560 -1905
rect 6494 -2579 6560 -1961
rect 6494 -2635 6499 -2579
rect 6555 -2635 6560 -2579
rect 6494 -2645 6560 -2635
rect 6809 -2208 6875 -2198
rect 6809 -2264 6814 -2208
rect 6870 -2264 6875 -2208
rect 5986 -2928 5991 -2872
rect 6047 -2928 6052 -2872
rect 5986 -2938 6052 -2928
rect 6809 -3327 6875 -2264
rect 6935 -2296 7001 -2286
rect 6935 -2352 6940 -2296
rect 6996 -2352 7001 -2296
rect 6935 -2952 7001 -2352
rect 6935 -3008 6940 -2952
rect 6996 -3008 7001 -2952
rect 6935 -3018 7001 -3008
rect 6809 -3383 6814 -3327
rect 6870 -3383 6875 -3327
rect 6809 -3388 6875 -3383
use cm2_ncell3  cm2_ncell3_0
timestamp 1750771847
transform 1 0 3595 0 1 -2894
box 1959 400 3647 1522
use cm2_ncell4  cm2_ncell4_0
timestamp 1750771847
transform 1 0 3934 0 1 -4128
box 454 531 3282 1740
use cm2_ncell  cm2_ncell_0
timestamp 1750771847
transform 1 0 3923 0 1 -2596
box -25 -646 1449 1272
use cm2_pcell3  cm2_pcell3_0
timestamp 1750201071
transform 1 0 12701 0 -1 5847
box -5785 3966 -1204 6082
use cm2_pcell4_1  cm2_pcell4_1_0
timestamp 1750204708
transform 1 0 7255 0 1 -133
box -339 -541 2041 90
use cm2_pcell4_2  cm2_pcell4_2_0
timestamp 1750205557
transform 1 0 8422 0 1 -775
box -1506 -499 -508 292
use cm2_pcell  cm2_pcell_0
timestamp 1750207421
transform 1 0 4022 0 1 568
box -154 -1842 3086 1314
<< labels >>
flabel metal1 s 7134 1669 7180 1701 0 FreeSans 480 0 0 0 ROUT
port 0 nsew
flabel metal2 s 7643 -1324 7703 -1264 0 FreeSans 480 0 0 0 VBPLV
port 1 nsew
flabel metal2 s 6368 -2559 6428 -2499 0 FreeSans 480 0 0 0 VBNLV
port 2 nsew
flabel metal2 s 6701 -1963 6761 -1903 0 FreeSans 320 0 0 0 VBPDEC
port 3 nsew
flabel metal2 s 5988 -2932 6048 -2872 0 FreeSans 320 0 0 0 VBNDEC
port 4 nsew
flabel metal1 s 3947 645 3981 679 0 FreeSans 320 0 0 0 VDDA
port 5 nsew
flabel metal1 s 3947 -1407 3981 -1373 0 FreeSans 320 0 0 0 GNDA
port 6 nsew
<< end >>
