magic
tech sky130A
magscale 1 2
timestamp 1751045299
<< nwell >>
rect 15213 13557 15995 14590
<< mvnsubdiff >>
rect 15279 14466 15929 14524
rect 15279 13681 15337 14466
rect 15871 13681 15929 14466
rect 15279 13623 15929 13681
<< locali >>
rect 15291 14478 15917 14512
rect 15291 13669 15325 14478
rect 15883 13669 15917 14478
rect 15291 13635 15917 13669
<< metal1 >>
rect 15657 14481 15709 14487
rect 15657 14412 15709 14429
rect 15499 14343 15551 14349
rect 15413 13747 15459 14329
rect 15657 14232 15709 14238
rect 15657 14167 15709 14180
rect 15499 14094 15551 14100
rect 15657 13983 15709 13989
rect 15657 13912 15709 13931
rect 15499 13845 15551 13851
rect 15749 13747 15795 14329
<< via1 >>
rect 15657 14429 15709 14481
rect 15499 14349 15551 14401
rect 15657 14180 15709 14232
rect 15499 14100 15551 14152
rect 15657 13931 15709 13983
rect 15499 13851 15551 13903
<< metal2 >>
rect 15651 14429 15657 14481
rect 15709 14429 15715 14481
rect 15493 14349 15499 14401
rect 15551 14349 15557 14401
rect 15651 14180 15657 14232
rect 15709 14180 15715 14232
rect 15493 14100 15499 14152
rect 15551 14100 15557 14152
rect 15651 13931 15657 13983
rect 15709 13931 15715 13983
rect 15493 13851 15499 13903
rect 15551 13851 15557 13903
use sky130_fd_pr__pfet_g5v0d10v5_Z832FA  sky130_fd_pr__pfet_g5v0d10v5_Z832FA_0
timestamp 1751042016
transform -1 0 15604 0 1 14074
box -253 -393 253 355
<< end >>
