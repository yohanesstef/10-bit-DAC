magic
tech sky130A
magscale 1 2
timestamp 1749567864
use hnmos_1  hnmos_1_0
timestamp 1749548291
transform 1 0 1122 0 1 -14
box -41 3 235 201
use hnmos_1  hnmos_1_1
timestamp 1749548291
transform 1 0 2530 0 1 -14
box -41 3 235 201
use hnmos_1  hnmos_1_2
timestamp 1749548291
transform 1 0 3938 0 1 -14
box -41 3 235 201
use hnmos_1  hnmos_1_3
timestamp 1749548291
transform 1 0 5346 0 1 -14
box -41 3 235 201
use hnmos_4  hnmos_4_0
timestamp 1749548291
transform 1 0 -15 0 1 -11
box -8 0 1096 198
use hnmos_4  hnmos_4_1
timestamp 1749548291
transform 1 0 1393 0 1 -11
box -8 0 1096 198
use hnmos_4  hnmos_4_2
timestamp 1749548291
transform 1 0 2801 0 1 -11
box -8 0 1096 198
use hnmos_4  hnmos_4_3
timestamp 1749548291
transform 1 0 4209 0 1 -11
box -8 0 1096 198
<< end >>
