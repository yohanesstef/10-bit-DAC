magic
tech sky130A
magscale 1 2
timestamp 1749234624
<< error_s >>
rect 2291 -2010 2349 -2004
rect 2291 -2044 2303 -2010
rect 2291 -2050 2349 -2044
rect 2291 -2222 2349 -2216
rect 2291 -2256 2303 -2222
rect 2291 -2262 2349 -2256
rect 2701 -3161 2726 -3061
rect 3237 -3135 3262 -3035
rect 3744 -3132 3769 -3032
rect 864 -8124 881 -7624
rect 918 -8173 935 -7673
rect 1385 -8219 1402 -7719
rect 1439 -8268 1456 -7768
rect 1906 -8314 1923 -7814
rect 1960 -8363 1977 -7863
rect 2427 -8409 2444 -7909
rect 2481 -8458 2498 -7958
rect 2948 -8504 2965 -8004
rect 3002 -8553 3019 -8053
rect 3469 -8599 3486 -8099
rect 3523 -8648 3540 -8148
rect 3990 -8694 4007 -8194
rect 4044 -8743 4061 -8243
<< nwell >>
rect 1544 -3334 4106 -2768
<< mvpmos >>
rect 3039 -3136 3123 -3036
rect 3334 -3135 3418 -3035
rect 3546 -3133 3630 -3033
rect 3841 -3132 3925 -3032
<< mvpdiff >>
rect 3039 -2990 3123 -2978
rect 3039 -3024 3051 -2990
rect 3111 -3024 3123 -2990
rect 3039 -3036 3123 -3024
rect 3334 -2989 3418 -2977
rect 3334 -3023 3346 -2989
rect 3406 -3023 3418 -2989
rect 3334 -3035 3418 -3023
rect 3546 -2987 3630 -2975
rect 3546 -3021 3558 -2987
rect 3618 -3021 3630 -2987
rect 3546 -3033 3630 -3021
rect 3841 -2986 3925 -2974
rect 3841 -3020 3853 -2986
rect 3913 -3020 3925 -2986
rect 3841 -3032 3925 -3020
rect 3039 -3148 3123 -3136
rect 3039 -3182 3051 -3148
rect 3111 -3182 3123 -3148
rect 3039 -3194 3123 -3182
rect 3334 -3147 3418 -3135
rect 3334 -3181 3346 -3147
rect 3406 -3181 3418 -3147
rect 3334 -3193 3418 -3181
rect 3546 -3145 3630 -3133
rect 3546 -3179 3558 -3145
rect 3618 -3179 3630 -3145
rect 3546 -3191 3630 -3179
rect 3841 -3144 3925 -3132
rect 3841 -3178 3853 -3144
rect 3913 -3178 3925 -3144
rect 3841 -3190 3925 -3178
<< mvpdiffc >>
rect 3051 -3024 3111 -2990
rect 3346 -3023 3406 -2989
rect 3558 -3021 3618 -2987
rect 3853 -3020 3913 -2986
rect 3051 -3182 3111 -3148
rect 3346 -3181 3406 -3147
rect 3558 -3179 3618 -3145
rect 3853 -3178 3913 -3144
<< poly >>
rect 3013 -3136 3039 -3036
rect 3123 -3052 3220 -3036
rect 3123 -3120 3170 -3052
rect 3204 -3120 3220 -3052
rect 3123 -3136 3220 -3120
rect 3237 -3051 3334 -3035
rect 3237 -3119 3253 -3051
rect 3287 -3119 3334 -3051
rect 3237 -3135 3334 -3119
rect 3418 -3135 3444 -3035
rect 3520 -3133 3546 -3033
rect 3630 -3049 3727 -3033
rect 3630 -3117 3677 -3049
rect 3711 -3117 3727 -3049
rect 3630 -3133 3727 -3117
rect 3744 -3048 3841 -3032
rect 3744 -3116 3760 -3048
rect 3794 -3116 3841 -3048
rect 3744 -3132 3841 -3116
rect 3925 -3132 3951 -3032
<< polycont >>
rect 3170 -3120 3204 -3052
rect 3253 -3119 3287 -3051
rect 3677 -3117 3711 -3049
rect 3760 -3116 3794 -3048
<< locali >>
rect 3035 -3024 3051 -2990
rect 3111 -3024 3127 -2990
rect 3330 -3023 3346 -2989
rect 3406 -3023 3422 -2989
rect 3542 -3021 3558 -2987
rect 3618 -3021 3634 -2987
rect 3837 -3020 3853 -2986
rect 3913 -3020 3929 -2986
rect 3170 -3052 3204 -3036
rect 3170 -3136 3204 -3120
rect 3253 -3051 3287 -3035
rect 3253 -3135 3287 -3119
rect 3677 -3049 3711 -3033
rect 3677 -3133 3711 -3117
rect 3760 -3048 3794 -3032
rect 3760 -3132 3794 -3116
rect 3035 -3182 3051 -3148
rect 3111 -3182 3127 -3148
rect 3330 -3181 3346 -3147
rect 3406 -3181 3422 -3147
rect 3542 -3179 3558 -3145
rect 3618 -3179 3634 -3145
rect 3837 -3178 3853 -3144
rect 3913 -3178 3929 -3144
<< viali >>
rect 3051 -3024 3111 -2990
rect 3346 -3023 3406 -2989
rect 3558 -3021 3618 -2987
rect 3853 -3020 3913 -2986
rect 3170 -3120 3204 -3052
rect 3253 -3119 3287 -3051
rect 3677 -3117 3711 -3049
rect 3760 -3116 3794 -3048
rect 3051 -3182 3111 -3148
rect 3346 -3181 3406 -3147
rect 3558 -3179 3618 -3145
rect 3853 -3178 3913 -3144
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 3039 -2990 3123 -2984
rect 0 -3200 200 -3000
rect 3039 -3024 3051 -2990
rect 3111 -3024 3123 -2990
rect 3039 -3030 3123 -3024
rect 3334 -2989 3418 -2983
rect 3334 -3023 3346 -2989
rect 3406 -3023 3418 -2989
rect 3334 -3029 3418 -3023
rect 3546 -2987 3630 -2981
rect 3546 -3021 3558 -2987
rect 3618 -3021 3630 -2987
rect 3546 -3027 3630 -3021
rect 3841 -2986 3925 -2980
rect 3841 -3020 3853 -2986
rect 3913 -3020 3925 -2986
rect 3841 -3026 3925 -3020
rect 3164 -3052 3210 -3040
rect 3164 -3120 3170 -3052
rect 3204 -3120 3210 -3052
rect 3164 -3132 3210 -3120
rect 3247 -3051 3293 -3039
rect 3247 -3119 3253 -3051
rect 3287 -3119 3293 -3051
rect 3247 -3131 3293 -3119
rect 3671 -3049 3717 -3037
rect 3671 -3117 3677 -3049
rect 3711 -3117 3717 -3049
rect 3671 -3129 3717 -3117
rect 3754 -3048 3800 -3036
rect 3754 -3116 3760 -3048
rect 3794 -3116 3800 -3048
rect 3754 -3128 3800 -3116
rect 3039 -3148 3123 -3142
rect 3039 -3182 3051 -3148
rect 3111 -3182 3123 -3148
rect 3039 -3188 3123 -3182
rect 3334 -3147 3418 -3141
rect 3334 -3181 3346 -3147
rect 3406 -3181 3418 -3147
rect 3334 -3187 3418 -3181
rect 3546 -3145 3630 -3139
rect 3546 -3179 3558 -3145
rect 3618 -3179 3630 -3145
rect 3546 -3185 3630 -3179
rect 3841 -3144 3925 -3138
rect 3841 -3178 3853 -3144
rect 3913 -3178 3925 -3144
rect 3841 -3184 3925 -3178
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
use rseg_3_v3  rseg_3_v3_0
timestamp 1749234624
transform 1 0 -10688 0 1 -1769
box 12478 -5378 17402 -1522
use sky130_fd_pr__pfet_01v8_M479BZ  sky130_fd_pr__pfet_01v8_M479BZ_0
timestamp 1749228705
transform 1 0 2320 0 1 -2133
box -211 -261 211 261
use sky130_fd_pr__pfet_g5v0d10v5_WJ97JY  sky130_fd_pr__pfet_g5v0d10v5_WJ97JY_0
timestamp 1749220931
transform -1 0 2306 0 1 -3077
box -174 -144 174 106
use sky130_fd_pr__pfet_g5v0d10v5_WJ97JY  sky130_fd_pr__pfet_g5v0d10v5_WJ97JY_1
timestamp 1749220931
transform 0 -1 2804 -1 0 -3111
box -174 -144 174 106
use sky130_fd_pr__pfet_g5v0d10v5_WJ97JY  sky130_fd_pr__pfet_g5v0d10v5_WJ97JY_2
timestamp 1749220931
transform 0 1 2581 -1 0 -3112
box -174 -144 174 106
use sky130_fd_pr__pfet_g5v0d10v5_WJ97JY  sky130_fd_pr__pfet_g5v0d10v5_WJ97JY_3
timestamp 1749220931
transform 0 1 3624 -1 0 -3083
box -174 -144 174 106
use sky130_fd_pr__pfet_g5v0d10v5_WJ97JY  sky130_fd_pr__pfet_g5v0d10v5_WJ97JY_4
timestamp 1749220931
transform 0 -1 3847 -1 0 -3082
box -174 -144 174 106
use sky130_fd_pr__pfet_g5v0d10v5_WJ97JY  sky130_fd_pr__pfet_g5v0d10v5_WJ97JY_5
timestamp 1749220931
transform 0 -1 3340 -1 0 -3085
box -174 -144 174 106
use sky130_fd_pr__pfet_g5v0d10v5_WJ97JY  sky130_fd_pr__pfet_g5v0d10v5_WJ97JY_6
timestamp 1749220931
transform 0 1 3117 -1 0 -3086
box -174 -144 174 106
use sky130_fd_pr__pfet_g5v0d10v5_WJ97JY  XM1
timestamp 1749220931
transform 1 0 2030 0 1 -3077
box -174 -144 174 106
use sky130_fd_pr__pfet_g5v0d10v5_5C2UEH  XM2
timestamp 1749220215
transform 1 0 639 0 1 -7851
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_5C2UEH  XM3
timestamp 1749220215
transform 1 0 1160 0 1 -7946
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_5C2UEH  XM4
timestamp 1749220215
transform 1 0 1681 0 1 -8041
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_5C2UEH  XM5
timestamp 1749220215
transform 1 0 2202 0 1 -8136
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_5C2UEH  XM6
timestamp 1749220215
transform 1 0 2723 0 1 -8231
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_5C2UEH  XM7
timestamp 1749220215
transform 1 0 3244 0 1 -8326
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_5C2UEH  XM8
timestamp 1749220215
transform 1 0 3765 0 1 -8421
box -308 -339 308 339
use sky130_fd_pr__pfet_g5v0d10v5_5C2UEH  XM9
timestamp 1749220215
transform 1 0 4286 0 1 -8516
box -308 -339 308 339
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 128 0 0 0 {vin\[0\]}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 128 0 0 0 {vin\[1\]}
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 128 0 0 0 {vin\[2\]}
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 128 0 0 0 {vin\[3\]}
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 128 0 0 0 {vin\[4\]}
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 128 0 0 0 {vin\[5\]}
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 128 0 0 0 {vin\[6\]}
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 128 0 0 0 {vin\[7\]}
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 128 0 0 0 {vin\[8\]}
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 128 0 0 0 DIN
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 128 0 0 0 {vout\[0\]}
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 128 0 0 0 {vout\[1\]}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 128 0 0 0 {vout\[2\]}
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 128 0 0 0 {vout\[3\]}
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 128 0 0 0 {}
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 128 0 0 0 {vout\[4\]}
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 128 0 0 0 {vout\[5\]}
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 128 0 0 0 {vout\[6\]}
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 128 0 0 0 {vout\[7\]}
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 128 0 0 0 {vout\[8\]}
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 128 0 0 0 VPB
port 20 nsew
<< end >>
