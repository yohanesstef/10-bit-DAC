magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1078 307 1078
<< psubdiff >>
rect -271 1008 -175 1042
rect 175 1008 271 1042
rect -271 946 -237 1008
rect 237 946 271 1008
rect -271 -1008 -237 -946
rect 237 -1008 271 -946
rect -271 -1042 -175 -1008
rect 175 -1042 271 -1008
<< psubdiffcont >>
rect -175 1008 175 1042
rect -271 -946 -237 946
rect 237 -946 271 946
rect -175 -1042 175 -1008
<< xpolycontact >>
rect -141 480 141 912
rect -141 -912 141 -480
<< xpolyres >>
rect -141 -480 141 480
<< locali >>
rect -271 1008 -175 1042
rect 175 1008 271 1042
rect -271 946 -237 1008
rect 237 946 271 1008
rect -271 -1008 -237 -946
rect 237 -1008 271 -946
rect -271 -1042 -175 -1008
rect 175 -1042 271 -1008
<< viali >>
rect -125 497 125 894
rect -125 -894 125 -497
<< metal1 >>
rect -131 894 131 906
rect -131 497 -125 894
rect 125 497 131 894
rect -131 485 131 497
rect -131 -497 131 -485
rect -131 -894 -125 -497
rect 125 -894 131 -497
rect -131 -906 131 -894
<< properties >>
string FIXED_BBOX -254 -1025 254 1025
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 4.962 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 7.305k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
