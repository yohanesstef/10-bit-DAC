magic
tech sky130A
magscale 1 2
timestamp 1749896124
use cm_pcell2_2_2  cm_pcell2_2_2_0
timestamp 1749896124
transform 1 0 6463 0 1 2673
box -31 -941 1709 943
use cm_pcell2_4_2  cm_pcell2_4_2_0
timestamp 1749896124
transform 1 0 3455 0 1 2673
box -31 -941 1621 943
use cm_pcell2_4_2  cm_pcell2_4_2_1
timestamp 1749896124
transform 1 0 4959 0 1 2673
box -31 -941 1621 943
<< end >>
