magic
tech sky130A
magscale 1 2
timestamp 1749548291
use hnmos_1  hnmos_1_0
timestamp 1749548291
transform 1 0 37 0 1 -2
box -41 3 235 201
use hnmos_1  hnmos_1_1
timestamp 1749548291
transform 1 0 313 0 1 -2
box -41 3 235 201
<< end >>
