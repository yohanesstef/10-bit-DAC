magic
tech sky130A
magscale 1 2
timestamp 1751030423
<< nwell >>
rect 4426 2776 5876 2777
rect 4244 2750 5876 2776
rect 4244 2153 4438 2750
<< metal1 >>
rect 4456 2832 4652 2852
rect 4188 2726 4652 2832
rect 4456 2688 4652 2726
rect 1964 -1656 2164 -588
rect 1964 -1844 1970 -1656
rect 2159 -1844 2164 -1656
rect 1964 -1850 2164 -1844
<< via1 >>
rect 6074 1278 6130 1334
rect 4736 1000 4792 1056
rect 1970 -1844 2159 -1656
<< metal2 >>
rect 420 1687 430 1743
rect 486 1687 496 1743
rect 1701 1334 1757 1344
rect 1701 1268 1757 1278
rect 6074 1334 6130 1344
rect 6074 1268 6130 1278
rect 1650 1112 1706 1122
rect 1650 1046 1706 1056
rect 4736 1056 4792 1066
rect 4736 990 4792 1000
rect 1964 -1656 3622 -1650
rect 1964 -1844 1970 -1656
rect 2159 -1844 3622 -1656
rect 1964 -1850 3622 -1844
rect 6599 -1889 6659 -1879
rect 6655 -1945 6659 -1889
rect 6599 -1970 6659 -1945
rect 5771 -2011 5827 -2001
rect 5771 -2077 5827 -2067
<< via2 >>
rect 430 1687 486 1743
rect 1701 1278 1757 1334
rect 6074 1278 6130 1334
rect 1650 1056 1706 1112
rect 4736 1000 4792 1056
rect 6599 -1945 6655 -1889
rect 5771 -2067 5827 -2011
<< metal3 >>
rect 425 1743 491 1753
rect 425 1687 430 1743
rect 486 1687 491 1743
rect 425 -2006 491 1687
rect 1691 1334 6140 1339
rect 1691 1278 1701 1334
rect 1757 1278 6074 1334
rect 6130 1278 6140 1334
rect 1691 1273 6140 1278
rect 1640 1112 4802 1117
rect 1640 1056 1650 1112
rect 1706 1056 4802 1112
rect 1640 1051 4736 1056
rect 4726 1000 4736 1051
rect 4792 1000 4802 1056
rect 4726 995 4802 1000
rect 1313 -1880 1379 530
rect 1313 -1884 6659 -1880
rect 1313 -1889 6665 -1884
rect 1313 -1945 6599 -1889
rect 6655 -1945 6665 -1889
rect 1313 -1946 6665 -1945
rect 6589 -1950 6665 -1946
rect 425 -2011 5837 -2006
rect 425 -2067 5771 -2011
rect 5827 -2067 5837 -2011
rect 425 -2072 5837 -2067
use top_bias_lvsf_dec  top_bias_lvsf_dec_0
timestamp 1751027542
transform 1 0 -5052 0 1 3009
box 3868 -3597 11497 1882
use top_digital_cell  top_digital_cell_0
timestamp 1751030423
transform 0 -1 5865 1 0 -22720
box 5366 -4551 25474 2301
<< end >>
