** sch_path: /home/yohanes/10-bit-DAC/xschem/top_segment_3.sch
.subckt top_segment_3 V0 V16 b[3] b[4] b[5] b[6] bb[3] bb[4] bb[5] bb[6] VH VL GND VPB
*.PININFO VH:O VPB:I b[3:6]:I VL:O bb[3:6]:I V16:I V0:I GND:I
x1 V0 V1 V2 V3 V4 V5 V6 V7 V8 bb[6] v1[0] v1[1] v1[2] v1[3] v1[4] v1[5] v1[6] v1[7] v1[8] VPB switch_pmos_1g_9o
x2 V8 V9 V10 V11 V12 V13 V14 V15 V16 b[6] v1[0] v1[1] v1[2] v1[3] v1[4] v1[5] v1[6] v1[7] v1[8] VPB switch_pmos_1g_9o
x3 v1[0] v1[1] v1[2] v1[3] v1[4] b[5] v2[0] v2[1] v2[2] v2[3] v2[4] VPB switch_pmos_1g_5o
x4 v1[4] v1[5] v1[6] v1[7] v1[8] bb[5] v2[0] v2[1] v2[2] v2[3] v2[4] VPB switch_pmos_1g_5o
x5 v2[0] v2[1] v2[2] b[4] v3[0] v3[1] v3[2] VPB switch_pmos_1g_3o
x6 v2[2] v2[3] v2[4] bb[4] v3[0] v3[1] v3[2] VPB switch_pmos_1g_3o
x7 v3[0] v3[1] b[3] VH VL VPB switch_pmos_1g_2o
x8 v3[1] v3[2] bb[3] VH VL VPB switch_pmos_1g_2o
x9 V0 V1 V2 V3 V4 V5 V6 V7 V8 V9 V10 V11 V12 V13 V14 V15 V16 GND rseg_3_v3
.ends

* expanding   symbol:  switch_pmos_1g_9o.sym # of pins=4
** sym_path: /home/yohanes/10-bit-DAC/xschem/switch_pmos_1g_9o.sym
** sch_path: /home/yohanes/10-bit-DAC/xschem/switch_pmos_1g_9o.sch
.subckt switch_pmos_1g_9o vin[0] vin[1] vin[2] vin[3] vin[4] vin[5] vin[6] vin[7] vin[8] DIN vout[0] vout[1] vout[2] vout[3]
+ vout[4] vout[5] vout[6] vout[7] vout[8] VPB
*.PININFO vin[0:8]:I vout[0:8]:O VPB:I DIN:I
.param wp=0.42 wn=0.42 l=0.5

XM1 vout[0] DIN vin[0] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM2 vout[1] DIN vin[1] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM3 vout[2] DIN vin[2] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM4 vout[3] DIN vin[3] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM5 vout[4] DIN vin[4] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM6 vout[5] DIN vin[5] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM7 vout[6] DIN vin[6] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM8 vout[7] DIN vin[7] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM9 vout[8] DIN vin[8] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
.ends


* expanding   symbol:  switch_pmos_1g_5o.sym # of pins=4
** sym_path: /home/yohanes/10-bit-DAC/xschem/switch_pmos_1g_5o.sym
** sch_path: /home/yohanes/10-bit-DAC/xschem/switch_pmos_1g_5o.sch
.subckt switch_pmos_1g_5o vin[0] vin[1] vin[2] vin[3] vin[4] DIN vout[0] vout[1] vout[2] vout[3] vout[4] VPB
*.PININFO vin[0:4]:I vout[0:4]:O VPB:I DIN:I
.param wp=0.42 wn=0.42 l=0.5

XM1 vout[0] DIN vin[0] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM2 vout[1] DIN vin[1] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM3 vout[2] DIN vin[2] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM4 vout[3] DIN vin[3] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM5 vout[4] DIN vin[4] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
.ends


* expanding   symbol:  switch_pmos_1g_3o.sym # of pins=4
** sym_path: /home/yohanes/10-bit-DAC/xschem/switch_pmos_1g_3o.sym
** sch_path: /home/yohanes/10-bit-DAC/xschem/switch_pmos_1g_3o.sch
.subckt switch_pmos_1g_3o vin[0] vin[1] vin[2] DIN vout[0] vout[1] vout[2] VPB
*.PININFO vin[0:2]:I vout[0:2]:O VPB:I DIN:I
.param wp=0.42 wn=0.42 l=0.5

XM1 vout[0] DIN vin[0] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM2 vout[1] DIN vin[1] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM3 vout[2] DIN vin[2] VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
.ends


* expanding   symbol:  switch_pmos_1g_2o.sym # of pins=5
** sym_path: /home/yohanes/10-bit-DAC/xschem/switch_pmos_1g_2o.sym
** sch_path: /home/yohanes/10-bit-DAC/xschem/switch_pmos_1g_2o.sch
.subckt switch_pmos_1g_2o vin0 vin1 DIN VH VL VPB
*.PININFO vin[0..1]:I VH:O VPB:I DIN:I VL:O
.param wp=0.42 wn=0.42 l=0.5

XM1 VL DIN vin0 VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
XM2 VH DIN vin1 VPB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 nf=1 m=1
.ends

