magic
tech sky130A
magscale 1 2
timestamp 1749525104
<< error_p >>
rect 138 567 144 573
rect 192 567 198 573
rect 2984 567 2990 573
rect 3038 567 3044 573
rect 132 561 138 567
rect 198 561 204 567
rect 2978 561 2984 567
rect 3044 561 3050 567
rect 132 507 138 513
rect 198 507 204 513
rect 2978 507 2984 513
rect 3044 507 3050 513
rect 138 501 144 507
rect 192 501 198 507
rect 2984 501 2990 507
rect 3038 501 3044 507
<< error_s >>
rect 1242 919 1248 925
rect 1296 919 1302 925
rect 1880 919 1886 925
rect 1934 919 1940 925
rect 1236 913 1242 919
rect 1302 913 1308 919
rect 1874 913 1880 919
rect 1940 913 1946 919
rect 1236 859 1242 865
rect 1302 859 1308 865
rect 1874 859 1880 865
rect 1940 859 1946 865
rect 1242 853 1248 859
rect 1296 853 1302 859
rect 1880 853 1886 859
rect 1934 853 1940 859
rect 966 831 972 837
rect 1020 831 1026 837
rect 2156 831 2162 837
rect 2210 831 2216 837
rect 960 825 966 831
rect 1026 825 1032 831
rect 2150 825 2156 831
rect 2216 825 2222 831
rect 960 771 966 777
rect 1026 771 1032 777
rect 2150 771 2156 777
rect 2216 771 2222 777
rect 966 765 972 771
rect 1020 765 1026 771
rect 2156 765 2162 771
rect 2210 765 2216 771
rect 690 743 696 749
rect 744 743 750 749
rect 2432 743 2438 749
rect 2486 743 2492 749
rect 684 737 690 743
rect 750 737 756 743
rect 2426 737 2432 743
rect 2492 737 2498 743
rect 684 683 690 689
rect 750 683 756 689
rect 2426 683 2432 689
rect 2492 683 2498 689
rect 690 677 696 683
rect 744 677 750 683
rect 2432 677 2438 683
rect 2486 677 2492 683
rect 414 655 420 661
rect 468 655 474 661
rect 2708 655 2714 661
rect 2762 655 2768 661
rect 408 649 414 655
rect 474 649 480 655
rect 2702 649 2708 655
rect 2768 649 2774 655
rect 408 595 414 601
rect 474 595 480 601
rect 2702 595 2708 601
rect 2768 595 2774 601
rect 414 589 420 595
rect 468 589 474 595
rect 2708 589 2714 595
rect 2762 589 2768 595
use hpmos_5  hpmos_5_0
timestamp 1749523501
transform 1 0 122 0 1 161
box -156 -170 1564 764
use hpmos_5  hpmos_5_1
timestamp 1749523501
transform -1 0 3060 0 1 161
box -156 -170 1564 764
<< end >>
