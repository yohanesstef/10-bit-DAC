magic
tech sky130A
magscale 1 2
timestamp 1751042016
<< mvnmos >>
rect -129 287 -29 371
rect 29 287 129 371
rect -129 47 -29 131
rect 29 47 129 131
rect -129 -193 -29 -109
rect 29 -193 129 -109
rect -129 -433 -29 -349
rect 29 -433 129 -349
<< mvndiff >>
rect -187 359 -129 371
rect -187 299 -175 359
rect -141 299 -129 359
rect -187 287 -129 299
rect -29 359 29 371
rect -29 299 -17 359
rect 17 299 29 359
rect -29 287 29 299
rect 129 359 187 371
rect 129 299 141 359
rect 175 299 187 359
rect 129 287 187 299
rect -187 119 -129 131
rect -187 59 -175 119
rect -141 59 -129 119
rect -187 47 -129 59
rect -29 119 29 131
rect -29 59 -17 119
rect 17 59 29 119
rect -29 47 29 59
rect 129 119 187 131
rect 129 59 141 119
rect 175 59 187 119
rect 129 47 187 59
rect -187 -121 -129 -109
rect -187 -181 -175 -121
rect -141 -181 -129 -121
rect -187 -193 -129 -181
rect -29 -121 29 -109
rect -29 -181 -17 -121
rect 17 -181 29 -121
rect -29 -193 29 -181
rect 129 -121 187 -109
rect 129 -181 141 -121
rect 175 -181 187 -121
rect 129 -193 187 -181
rect -187 -361 -129 -349
rect -187 -421 -175 -361
rect -141 -421 -129 -361
rect -187 -433 -129 -421
rect -29 -361 29 -349
rect -29 -421 -17 -361
rect 17 -421 29 -361
rect -29 -433 29 -421
rect 129 -361 187 -349
rect 129 -421 141 -361
rect 175 -421 187 -361
rect 129 -433 187 -421
<< mvndiffc >>
rect -175 299 -141 359
rect -17 299 17 359
rect 141 299 175 359
rect -175 59 -141 119
rect -17 59 17 119
rect 141 59 175 119
rect -175 -181 -141 -121
rect -17 -181 17 -121
rect 141 -181 175 -121
rect -175 -421 -141 -361
rect -17 -421 17 -361
rect 141 -421 175 -361
<< poly >>
rect -129 443 -29 459
rect -129 409 -113 443
rect -45 409 -29 443
rect -129 371 -29 409
rect 29 443 129 459
rect 29 409 45 443
rect 113 409 129 443
rect 29 371 129 409
rect -129 261 -29 287
rect 29 261 129 287
rect -129 203 -29 219
rect -129 169 -113 203
rect -45 169 -29 203
rect -129 131 -29 169
rect 29 203 129 219
rect 29 169 45 203
rect 113 169 129 203
rect 29 131 129 169
rect -129 21 -29 47
rect 29 21 129 47
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect -129 -219 -29 -193
rect 29 -219 129 -193
rect -129 -277 -29 -261
rect -129 -311 -113 -277
rect -45 -311 -29 -277
rect -129 -349 -29 -311
rect 29 -277 129 -261
rect 29 -311 45 -277
rect 113 -311 129 -277
rect 29 -349 129 -311
rect -129 -459 -29 -433
rect 29 -459 129 -433
<< polycont >>
rect -113 409 -45 443
rect 45 409 113 443
rect -113 169 -45 203
rect 45 169 113 203
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect -113 -311 -45 -277
rect 45 -311 113 -277
<< locali >>
rect -129 409 -113 443
rect -45 409 -29 443
rect 29 409 45 443
rect 113 409 129 443
rect -175 359 -141 375
rect -175 283 -141 299
rect -17 359 17 375
rect -17 283 17 299
rect 141 359 175 375
rect 141 283 175 299
rect -129 169 -113 203
rect -45 169 -29 203
rect 29 169 45 203
rect 113 169 129 203
rect -175 119 -141 135
rect -175 43 -141 59
rect -17 119 17 135
rect -17 43 17 59
rect 141 119 175 135
rect 141 43 175 59
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect -175 -121 -141 -105
rect -175 -197 -141 -181
rect -17 -121 17 -105
rect -17 -197 17 -181
rect 141 -121 175 -105
rect 141 -197 175 -181
rect -129 -311 -113 -277
rect -45 -311 -29 -277
rect 29 -311 45 -277
rect 113 -311 129 -277
rect -175 -361 -141 -345
rect -175 -437 -141 -421
rect -17 -361 17 -345
rect -17 -437 17 -421
rect 141 -361 175 -345
rect 141 -437 175 -421
<< viali >>
rect -105 409 -53 443
rect 53 409 105 443
rect -175 299 -141 359
rect -17 299 17 359
rect 141 299 175 359
rect -105 169 -53 203
rect 53 169 105 203
rect -175 59 -141 119
rect -17 59 17 119
rect 141 59 175 119
rect -105 -71 -53 -37
rect 53 -71 105 -37
rect -175 -181 -141 -121
rect -17 -181 17 -121
rect 141 -181 175 -121
rect -105 -311 -53 -277
rect 53 -311 105 -277
rect -175 -421 -141 -361
rect -17 -421 17 -361
rect 141 -421 175 -361
<< metal1 >>
rect -117 443 -41 449
rect -117 409 -105 443
rect -53 409 -41 443
rect -117 403 -41 409
rect 41 443 117 449
rect 41 409 53 443
rect 105 409 117 443
rect 41 403 117 409
rect -181 359 -135 371
rect -181 299 -175 359
rect -141 299 -135 359
rect -181 287 -135 299
rect -23 359 23 371
rect -23 299 -17 359
rect 17 299 23 359
rect -23 287 23 299
rect 135 359 181 371
rect 135 299 141 359
rect 175 299 181 359
rect 135 287 181 299
rect -117 203 -41 209
rect -117 169 -105 203
rect -53 169 -41 203
rect -117 163 -41 169
rect 41 203 117 209
rect 41 169 53 203
rect 105 169 117 203
rect 41 163 117 169
rect -181 119 -135 131
rect -181 59 -175 119
rect -141 59 -135 119
rect -181 47 -135 59
rect -23 119 23 131
rect -23 59 -17 119
rect 17 59 23 119
rect -23 47 23 59
rect 135 119 181 131
rect 135 59 141 119
rect 175 59 181 119
rect 135 47 181 59
rect -117 -37 -41 -31
rect -117 -71 -105 -37
rect -53 -71 -41 -37
rect -117 -77 -41 -71
rect 41 -37 117 -31
rect 41 -71 53 -37
rect 105 -71 117 -37
rect 41 -77 117 -71
rect -181 -121 -135 -109
rect -181 -181 -175 -121
rect -141 -181 -135 -121
rect -181 -193 -135 -181
rect -23 -121 23 -109
rect -23 -181 -17 -121
rect 17 -181 23 -121
rect -23 -193 23 -181
rect 135 -121 181 -109
rect 135 -181 141 -121
rect 175 -181 181 -121
rect 135 -193 181 -181
rect -117 -277 -41 -271
rect -117 -311 -105 -277
rect -53 -311 -41 -277
rect -117 -317 -41 -311
rect 41 -277 117 -271
rect 41 -311 53 -277
rect 105 -311 117 -277
rect 41 -317 117 -311
rect -181 -361 -135 -349
rect -181 -421 -175 -361
rect -141 -421 -135 -361
rect -181 -433 -135 -421
rect -23 -361 23 -349
rect -23 -421 -17 -361
rect 17 -421 23 -361
rect -23 -433 23 -421
rect 135 -361 181 -349
rect 135 -421 141 -361
rect 175 -421 181 -361
rect 135 -433 181 -421
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.420 l 0.50 m 4 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
