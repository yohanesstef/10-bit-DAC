magic
tech sky130A
magscale 1 2
timestamp 1750840520
<< magnet >>
rect 5029 -3512 5087 -3466
<< pwell >>
rect 4625 -2855 6825 -2667
rect 4625 -3696 6825 -3531
<< locali >>
rect 5058 -2891 5063 -2857
rect 5097 -2891 5104 -2857
rect 5058 -2892 5104 -2891
rect 5058 -2911 5102 -2892
rect 5061 -3472 5103 -3469
rect 5075 -3506 5103 -3472
rect 5061 -3519 5103 -3506
<< viali >>
rect 6024 -2780 6058 -2746
rect 4836 -2910 4870 -2876
rect 5063 -2891 5097 -2857
rect 5279 -2910 5313 -2876
rect 5487 -2891 5521 -2857
rect 5656 -2895 5690 -2861
rect 5753 -2910 5787 -2876
rect 5921 -2910 5955 -2876
rect 6033 -2910 6067 -2876
rect 6262 -2903 6296 -2869
rect 5573 -2990 5607 -2956
rect 5205 -3046 5239 -3012
rect 6347 -3052 6381 -3018
rect 4929 -3102 4963 -3068
rect 5750 -3429 5784 -3395
rect 4841 -3509 4875 -3475
rect 5041 -3506 5075 -3472
rect 5292 -3509 5326 -3475
rect 5477 -3518 5511 -3484
rect 5761 -3518 5795 -3484
rect 5894 -3510 5928 -3476
rect 5990 -3513 6024 -3479
rect 6125 -3509 6159 -3475
rect 6296 -3509 6330 -3475
rect 6399 -3509 6433 -3475
rect 5202 -3560 5236 -3526
rect 5635 -3575 5669 -3541
rect 6198 -3596 6232 -3562
rect 5019 -3645 5053 -3611
rect 5733 -3647 5767 -3613
<< metal1 >>
rect 6012 -2746 6070 -2740
rect 4359 -2810 4365 -2758
rect 4417 -2786 5687 -2758
rect 6012 -2780 6024 -2746
rect 6058 -2758 6070 -2746
rect 6058 -2780 6289 -2758
rect 6012 -2786 6289 -2780
rect 4417 -2810 4423 -2786
rect 4543 -2866 4549 -2814
rect 4601 -2842 5533 -2814
rect 4601 -2866 4607 -2842
rect 5051 -2857 5109 -2842
rect 4451 -2922 4457 -2870
rect 4509 -2894 4515 -2870
rect 4824 -2876 4882 -2870
rect 4824 -2894 4836 -2876
rect 4509 -2910 4836 -2894
rect 4870 -2910 4882 -2876
rect 5051 -2891 5063 -2857
rect 5097 -2891 5109 -2857
rect 5475 -2857 5533 -2842
rect 5659 -2855 5687 -2786
rect 5051 -2897 5109 -2891
rect 5267 -2876 5325 -2870
rect 4509 -2922 4882 -2910
rect 5267 -2910 5279 -2876
rect 5313 -2910 5325 -2876
rect 5475 -2891 5487 -2857
rect 5521 -2891 5533 -2857
rect 5475 -2897 5533 -2891
rect 5644 -2861 5702 -2855
rect 5644 -2895 5656 -2861
rect 5690 -2895 5702 -2861
rect 6261 -2863 6289 -2786
rect 6250 -2869 6308 -2863
rect 5644 -2901 5702 -2895
rect 5741 -2876 5799 -2870
rect 5267 -2916 5325 -2910
rect 5741 -2910 5753 -2876
rect 5787 -2910 5799 -2876
rect 5741 -2916 5799 -2910
rect 5909 -2876 5967 -2870
rect 5909 -2910 5921 -2876
rect 5955 -2910 5967 -2876
rect 5909 -2916 5967 -2910
rect 6021 -2876 6079 -2870
rect 6021 -2910 6033 -2876
rect 6067 -2910 6079 -2876
rect 6250 -2903 6262 -2869
rect 6296 -2903 6308 -2869
rect 6250 -2909 6308 -2903
rect 6021 -2916 6079 -2910
rect 4267 -2978 4273 -2926
rect 4325 -2950 4331 -2926
rect 5281 -2950 5309 -2916
rect 4325 -2978 5309 -2950
rect 5561 -2956 5619 -2950
rect 5561 -2990 5573 -2956
rect 5607 -2968 5619 -2956
rect 5771 -2968 5799 -2916
rect 5607 -2990 5799 -2968
rect 5561 -2996 5799 -2990
rect 5193 -3012 5251 -3006
rect 5193 -3046 5205 -3012
rect 5239 -3024 5251 -3012
rect 5939 -3024 5967 -2916
rect 5239 -3046 5967 -3024
rect 5193 -3052 5967 -3046
rect 4917 -3068 4975 -3062
rect 4917 -3102 4929 -3068
rect 4963 -3080 4975 -3068
rect 6051 -3080 6079 -2916
rect 4963 -3102 6079 -3080
rect 4917 -3108 6079 -3102
rect 6260 -3086 6288 -2909
rect 6335 -3018 6393 -3012
rect 6335 -3052 6347 -3018
rect 6381 -3030 6393 -3018
rect 7477 -3026 7541 -2998
rect 7477 -3030 7505 -3026
rect 6381 -3052 7505 -3030
rect 6335 -3058 7505 -3052
rect 6260 -3114 7541 -3086
rect 3899 -3148 4622 -3142
rect 4055 -3232 4622 -3148
rect 3899 -3238 4622 -3232
rect 6830 -3148 7357 -3142
rect 6830 -3232 7201 -3148
rect 6830 -3238 7357 -3232
rect 4267 -3409 4273 -3357
rect 4325 -3385 5308 -3357
rect 4325 -3409 4331 -3385
rect 4451 -3465 4457 -3413
rect 4509 -3441 5072 -3413
rect 4509 -3465 4515 -3441
rect 5029 -3466 5072 -3441
rect 4359 -3521 4365 -3469
rect 4417 -3493 4423 -3469
rect 4829 -3475 4887 -3469
rect 4829 -3493 4841 -3475
rect 4417 -3509 4841 -3493
rect 4875 -3509 4887 -3475
rect 4417 -3521 4887 -3509
rect 5029 -3472 5087 -3466
rect 5029 -3506 5041 -3472
rect 5075 -3506 5087 -3472
rect 5029 -3512 5087 -3506
rect 5280 -3469 5308 -3385
rect 5744 -3395 5790 -3383
rect 5744 -3429 5750 -3395
rect 5784 -3413 5790 -3395
rect 6136 -3385 7023 -3357
rect 5784 -3429 5916 -3413
rect 5744 -3441 5916 -3429
rect 5888 -3464 5916 -3441
rect 5280 -3475 5338 -3469
rect 5280 -3509 5292 -3475
rect 5326 -3509 5338 -3475
rect 5196 -3526 5242 -3514
rect 5280 -3515 5338 -3509
rect 5465 -3484 5523 -3478
rect 5196 -3560 5202 -3526
rect 5236 -3560 5242 -3526
rect 5196 -3567 5242 -3560
rect 5465 -3518 5477 -3484
rect 5511 -3518 5523 -3484
rect 5465 -3524 5523 -3518
rect 5755 -3484 5801 -3472
rect 5755 -3518 5761 -3484
rect 5795 -3502 5801 -3484
rect 5888 -3476 5934 -3464
rect 5795 -3518 5854 -3502
rect 5465 -3567 5493 -3524
rect 5755 -3530 5854 -3518
rect 5888 -3510 5894 -3476
rect 5928 -3510 5934 -3476
rect 5888 -3522 5934 -3510
rect 5982 -3470 6034 -3464
rect 6136 -3469 6164 -3385
rect 7017 -3409 7023 -3385
rect 7075 -3409 7081 -3357
rect 6290 -3441 6931 -3413
rect 6290 -3469 6318 -3441
rect 6925 -3465 6931 -3441
rect 6983 -3465 6989 -3413
rect 6113 -3475 6171 -3469
rect 6113 -3509 6125 -3475
rect 6159 -3509 6171 -3475
rect 6113 -3515 6171 -3509
rect 6284 -3475 6342 -3469
rect 6284 -3509 6296 -3475
rect 6330 -3509 6342 -3475
rect 6284 -3515 6342 -3509
rect 6387 -3475 6839 -3469
rect 6387 -3509 6399 -3475
rect 6433 -3497 6839 -3475
rect 6433 -3509 6445 -3497
rect 6387 -3515 6445 -3509
rect 6833 -3521 6839 -3497
rect 6891 -3521 6897 -3469
rect 5982 -3528 6034 -3522
rect 5196 -3595 5493 -3567
rect 5623 -3541 5681 -3535
rect 5623 -3575 5635 -3541
rect 5669 -3575 5681 -3541
rect 5623 -3581 5681 -3575
rect 5826 -3567 5854 -3530
rect 6184 -3562 6244 -3556
rect 6184 -3567 6198 -3562
rect 5007 -3611 5065 -3605
rect 5007 -3645 5019 -3611
rect 5053 -3623 5065 -3611
rect 5623 -3623 5651 -3581
rect 5826 -3595 6198 -3567
rect 6184 -3596 6198 -3595
rect 6232 -3596 6244 -3562
rect 6184 -3602 6244 -3596
rect 6478 -3584 6484 -3532
rect 6536 -3574 6542 -3532
rect 7489 -3574 7541 -3542
rect 6536 -3584 7541 -3574
rect 6478 -3602 7541 -3584
rect 5053 -3645 5651 -3623
rect 5007 -3651 5651 -3645
rect 5714 -3613 5779 -3606
rect 5714 -3647 5733 -3613
rect 5767 -3630 5779 -3613
rect 5767 -3647 7541 -3630
rect 5714 -3658 7541 -3647
rect 4083 -3692 4651 -3686
rect 4239 -3776 4651 -3692
rect 4083 -3782 4651 -3776
rect 6830 -3692 7541 -3686
rect 6830 -3776 7385 -3692
rect 6830 -3782 7541 -3776
<< via1 >>
rect 4365 -2810 4417 -2758
rect 4549 -2866 4601 -2814
rect 4457 -2922 4509 -2870
rect 4273 -2978 4325 -2926
rect 3899 -3232 4055 -3148
rect 7201 -3232 7357 -3148
rect 4273 -3409 4325 -3357
rect 4457 -3465 4509 -3413
rect 4365 -3521 4417 -3469
rect 7023 -3409 7075 -3357
rect 6931 -3465 6983 -3413
rect 5982 -3479 6034 -3470
rect 5982 -3513 5990 -3479
rect 5990 -3513 6024 -3479
rect 6024 -3513 6034 -3479
rect 5982 -3522 6034 -3513
rect 6839 -3521 6891 -3469
rect 6484 -3584 6536 -3532
rect 4083 -3776 4239 -3692
rect 7385 -3776 7541 -3692
<< metal2 >>
rect 3899 -3148 4055 -2598
rect 3899 -3782 4055 -3232
rect 4083 -3692 4239 -2598
rect 4083 -3782 4239 -3776
rect 4267 -2926 4331 -2694
rect 4267 -2978 4273 -2926
rect 4325 -2978 4331 -2926
rect 4267 -3357 4331 -2978
rect 4267 -3409 4273 -3357
rect 4325 -3409 4331 -3357
rect 4267 -3782 4331 -3409
rect 4359 -2758 4423 -2694
rect 4359 -2810 4365 -2758
rect 4417 -2810 4423 -2758
rect 4359 -3469 4423 -2810
rect 4359 -3521 4365 -3469
rect 4417 -3521 4423 -3469
rect 4359 -3782 4423 -3521
rect 4451 -2870 4515 -2694
rect 4451 -2922 4457 -2870
rect 4509 -2922 4515 -2870
rect 4451 -3413 4515 -2922
rect 4451 -3465 4457 -3413
rect 4509 -3465 4515 -3413
rect 4451 -3782 4515 -3465
rect 4543 -2814 4607 -2694
rect 4543 -2866 4549 -2814
rect 4601 -2866 4607 -2814
rect 4543 -3782 4607 -2866
rect 5982 -3470 6034 -3464
rect 5982 -3528 6034 -3522
rect 5994 -3532 6034 -3528
rect 6833 -3469 6897 -2694
rect 6833 -3521 6839 -3469
rect 6891 -3521 6897 -3469
rect 5994 -3560 6484 -3532
rect 6478 -3584 6484 -3560
rect 6536 -3584 6542 -3532
rect 6833 -3782 6897 -3521
rect 6925 -3413 6989 -2694
rect 6925 -3465 6931 -3413
rect 6983 -3465 6989 -3413
rect 6925 -3782 6989 -3465
rect 7017 -3357 7081 -2694
rect 7017 -3409 7023 -3357
rect 7075 -3409 7081 -3357
rect 7017 -3782 7081 -3409
rect 7109 -3782 7173 -2694
rect 7201 -3148 7357 -2598
rect 7201 -3782 7357 -3232
rect 7385 -3692 7541 -2598
rect 7385 -3782 7541 -3776
use sky130_ef_sc_hd__fill_4  sky130_ef_sc_hd__fill_4_0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6462 0 -1 -2646
box -38 -48 406 592
use sky130_ef_sc_hd__fill_4  sky130_ef_sc_hd__fill_4_1
timestamp 1704896540
transform -1 0 6830 0 1 -3734
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5358 0 -1 -2646
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1704896540
transform 1 0 6094 0 -1 -2646
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1704896540
transform 1 0 5358 0 1 -3734
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1704896540
transform 1 0 4714 0 -1 -2646
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1704896540
transform 1 0 4622 0 -1 -2646
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1704896540
transform 1 0 4622 0 1 -3734
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1704896540
transform 1 0 4714 0 1 -3734
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  x1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4806 0 -1 -2646
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x2
timestamp 1704896540
transform 1 0 5082 0 -1 -2646
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x3
timestamp 1704896540
transform 1 0 5450 0 -1 -2646
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  x4 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1749714889
transform 1 0 5726 0 -1 -2646
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  x5
timestamp 1749714889
transform 1 0 5450 0 1 -3734
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  x6
timestamp 1704896540
transform 1 0 4806 0 1 -3734
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x7
timestamp 1704896540
transform 1 0 5082 0 1 -3734
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  x8
timestamp 1749714889
transform 1 0 6094 0 1 -3734
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  x9 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1749714889
transform 1 0 6186 0 -1 -2646
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x10
timestamp 1749714889
transform 1 0 5818 0 1 -3734
box -38 -48 314 592
<< labels >>
flabel metal2 s 4267 -2704 4267 -2704 3 FreeSans 320 0 0 0 b[6]
port 0 e
flabel metal2 s 4359 -2704 4359 -2704 3 FreeSans 320 0 0 0 b[7]
port 1 e
flabel metal2 s 4451 -2704 4451 -2704 3 FreeSans 320 0 0 0 b[8]
port 2 e
flabel metal2 s 4543 -2704 4543 -2704 3 FreeSans 320 0 0 0 b[9]
port 3 e
flabel metal2 s 6833 -2707 6833 -2707 3 FreeSans 240 0 0 0 bb[6]
port 4 e
flabel metal2 s 6925 -2707 6925 -2707 3 FreeSans 240 0 0 0 bb[7]
port 5 e
flabel metal2 s 7017 -2707 7017 -2707 3 FreeSans 240 0 0 0 bb[8]
port 6 e
flabel metal2 s 3900 -2614 3900 -2614 3 FreeSans 240 0 0 0 VDD
port 11 e
flabel metal2 s 4085 -2614 4085 -2614 3 FreeSans 240 0 0 0 GND
port 12 e
flabel metal1 s 7501 -3557 7501 -3557 3 FreeSans 240 0 0 0 BSB[8]
port 9 e
flabel metal1 s 7508 -3646 7508 -3646 3 FreeSans 240 0 0 0 BS[8]
port 7 e
flabel metal1 s 7512 -3100 7512 -3100 3 FreeSans 240 0 0 0 BS[9]
port 8 e
flabel metal1 s 7513 -3011 7513 -3011 3 FreeSans 240 0 0 0 BSB[9]
port 10 e
<< end >>
