magic
tech sky130A
magscale 1 2
timestamp 1749642965
<< mvnmos >>
rect -100 -131 100 69
<< mvndiff >>
rect -158 13 -100 69
rect -158 -75 -146 13
rect -112 -75 -100 13
rect -158 -131 -100 -75
rect 100 13 158 69
rect 100 -75 112 13
rect 146 -75 158 13
rect 100 -131 158 -75
<< mvndiffc >>
rect -146 -75 -112 13
rect 112 -75 146 13
<< poly >>
rect -58 141 58 157
rect -58 124 -42 141
rect -100 107 -42 124
rect 42 124 58 141
rect 42 107 100 124
rect -100 69 100 107
rect -100 -157 100 -131
<< polycont >>
rect -42 107 42 141
<< viali >>
rect -84 107 -42 141
rect -42 107 42 141
rect 42 107 84 141
rect -146 13 -112 57
rect -146 -75 -112 13
rect -146 -119 -112 -75
rect 112 13 146 57
rect 112 -75 146 13
rect 112 -119 146 -75
<< metal1 >>
rect -96 141 96 147
rect -96 107 -84 141
rect 84 107 96 141
rect -96 101 96 107
rect -152 57 -106 69
rect -152 -119 -146 57
rect -112 -119 -106 57
rect -152 -131 -106 -119
rect 106 57 152 69
rect 106 -119 112 57
rect 146 -119 152 57
rect 106 -131 152 -119
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 1 nf 1 diffcov 50 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
