magic
tech sky130A
timestamp 1749716031
<< magnet >>
rect 29 1450 43 1464
rect -3 1418 29 1450
rect 43 1418 75 1450
rect 89 1418 121 1450
rect 135 1418 167 1450
rect 29 1404 43 1418
rect -3 1372 29 1404
rect 43 1372 75 1404
rect 89 1372 121 1404
rect 135 1372 167 1404
rect 29 1358 43 1372
rect -3 1326 29 1358
rect 43 1326 75 1358
rect 89 1326 121 1358
rect 135 1326 167 1358
rect 29 1312 43 1326
rect -3 1280 29 1312
rect 43 1280 75 1312
rect 89 1280 121 1312
rect 135 1280 167 1312
rect 29 1266 43 1280
rect -3 1234 29 1266
rect 43 1234 75 1266
rect 89 1234 121 1266
rect 135 1234 167 1266
rect 29 1220 43 1234
rect -3 1188 29 1220
rect 43 1188 75 1220
rect 89 1188 121 1220
rect 135 1188 167 1220
rect 29 1174 43 1188
rect -3 1142 29 1174
rect 43 1142 75 1174
rect 89 1142 121 1174
rect 135 1142 167 1174
rect 29 1128 43 1142
rect -3 1096 29 1128
rect 43 1096 75 1128
rect 89 1096 121 1128
rect 135 1096 167 1128
rect 29 1082 43 1096
rect -3 1050 29 1082
rect 43 1050 75 1082
rect 89 1050 121 1082
rect 135 1050 167 1082
rect 29 1036 43 1050
rect -3 1004 29 1036
rect 43 1004 75 1036
rect 89 1004 121 1036
rect 135 1004 167 1036
rect 29 990 43 1004
rect -3 958 29 990
rect 43 958 75 990
rect 89 958 121 990
rect 135 958 167 990
rect 29 944 43 958
rect -3 912 29 944
rect 43 912 75 944
rect 89 912 121 944
rect 135 912 167 944
rect 29 898 43 912
rect -3 866 29 898
rect 43 866 75 898
rect 89 866 121 898
rect 135 866 167 898
rect 29 852 43 866
rect -3 820 29 852
rect 43 820 75 852
rect 89 820 121 852
rect 135 820 167 852
rect 29 806 43 820
rect -3 774 29 806
rect 43 774 75 806
rect 89 774 121 806
rect 135 774 167 806
rect 29 760 43 774
rect -3 728 29 760
rect 43 728 75 760
rect 89 728 121 760
rect 135 728 167 760
rect 29 714 43 728
rect -3 682 29 714
rect 43 682 75 714
rect 89 682 121 714
rect 135 682 167 714
rect 29 668 43 682
rect -3 636 29 668
rect 43 636 75 668
rect 89 636 121 668
rect 135 636 167 668
rect 29 622 43 636
rect -3 590 29 622
rect 43 590 75 622
rect 89 590 121 622
rect 135 590 167 622
rect 29 576 43 590
rect -3 544 29 576
rect 43 544 75 576
rect 89 544 121 576
rect 135 544 167 576
rect 29 530 43 544
rect -3 498 29 530
rect 43 498 75 530
rect 89 498 121 530
rect 135 498 167 530
rect 29 484 43 498
rect -3 452 29 484
rect 43 452 75 484
rect 89 452 121 484
rect 135 452 167 484
rect 29 438 43 452
rect -3 406 29 438
rect 43 406 75 438
rect 89 406 121 438
rect 135 406 167 438
rect 29 392 43 406
rect -3 360 29 392
rect 43 360 75 392
rect 89 360 121 392
rect 135 360 167 392
rect 29 346 43 360
rect -3 314 29 346
rect 43 314 75 346
rect 89 314 121 346
rect 135 314 167 346
rect 29 300 43 314
rect -3 268 29 300
rect 43 268 75 300
rect 89 268 121 300
rect 135 268 167 300
rect 29 254 43 268
rect -3 222 29 254
rect 43 222 75 254
rect 89 222 121 254
rect 135 222 167 254
rect 29 208 43 222
rect -3 176 29 208
rect 43 176 75 208
rect 89 176 121 208
rect 135 176 167 208
rect 29 162 43 176
rect -3 130 29 162
rect 43 130 75 162
rect 89 130 121 162
rect 135 130 167 162
rect 29 116 43 130
rect -3 84 29 116
rect 43 84 75 116
rect 89 84 121 116
rect 135 84 167 116
rect 29 70 43 84
rect -3 38 29 70
rect 43 38 75 70
rect 89 38 121 70
rect 135 38 167 70
rect 29 24 43 38
rect -3 -8 29 24
rect 43 -8 75 24
rect 89 -8 121 24
rect 135 -8 167 24
<< end >>
