magic
tech sky130A
magscale 1 2
timestamp 1749057406
<< pwell >>
rect -307 -991 307 991
<< psubdiff >>
rect -271 921 -175 955
rect 175 921 271 955
rect -271 859 -237 921
rect 237 859 271 921
rect -271 -921 -237 -859
rect 237 -921 271 -859
rect -271 -955 -175 -921
rect 175 -955 271 -921
<< psubdiffcont >>
rect -175 921 175 955
rect -271 -859 -237 859
rect 237 -859 271 859
rect -175 -955 175 -921
<< xpolycontact >>
rect -141 393 141 825
rect -141 -825 141 -393
<< xpolyres >>
rect -141 -393 141 393
<< locali >>
rect -271 921 -175 955
rect 175 921 271 955
rect -271 859 -237 921
rect 237 859 271 921
rect -271 -921 -237 -859
rect 237 -921 271 -859
rect -271 -955 -175 -921
rect 175 -955 271 -921
<< viali >>
rect -125 410 125 807
rect -125 -807 125 -410
<< metal1 >>
rect -131 807 131 819
rect -131 410 -125 807
rect 125 410 131 807
rect -131 398 131 410
rect -131 -410 131 -398
rect -131 -807 -125 -410
rect 125 -807 131 -410
rect -131 -819 131 -807
<< properties >>
string FIXED_BBOX -254 -938 254 938
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 4.09 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 6.068k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
