magic
tech sky130A
magscale 1 2
timestamp 1749801796
<< pwell >>
rect 363 -466 1425 310
<< psubdiff >>
rect 399 -383 1389 -370
rect 399 -417 445 -383
rect 1343 -417 1389 -383
rect 399 -430 1389 -417
<< psubdiffcont >>
rect 445 -417 1343 -383
<< poly >>
rect 835 -273 865 -268
rect 769 -289 865 -273
rect 769 -323 785 -289
rect 819 -323 865 -289
rect 769 -339 865 -323
rect 923 -273 953 -268
rect 923 -289 1019 -273
rect 923 -323 969 -289
rect 1003 -323 1019 -289
rect 923 -339 1019 -323
<< polycont >>
rect 785 -323 819 -289
rect 969 -323 1003 -289
<< locali >>
rect 769 -323 785 -289
rect 819 -323 835 -289
rect 953 -323 969 -289
rect 1003 -323 1019 -289
rect 429 -417 445 -383
rect 1343 -417 1359 -383
<< viali >>
rect 785 -323 819 -289
rect 969 -323 1003 -289
rect 445 -417 1343 -383
<< metal1 >>
rect 772 -276 832 -270
rect 772 -342 832 -336
rect 864 -370 924 358
rect 956 -276 1016 -270
rect 956 -342 1016 -336
rect 399 -383 1389 -370
rect 399 -417 445 -383
rect 1343 -417 1389 -383
rect 399 -430 1389 -417
<< via1 >>
rect 772 -289 832 -276
rect 772 -323 785 -289
rect 785 -323 819 -289
rect 819 -323 832 -289
rect 772 -336 832 -323
rect 956 -289 1016 -276
rect 956 -323 969 -289
rect 969 -323 1003 -289
rect 1003 -323 1016 -289
rect 956 -336 1016 -323
<< metal2 >>
rect 772 -276 832 -270
rect 772 -342 832 -336
rect 956 -276 1016 -270
rect 956 -342 1016 -336
use sky130_fd_pr__nfet_01v8_AT5T57  sky130_fd_pr__nfet_01v8_AT5T57_0
timestamp 1749624948
transform 1 0 850 0 1 58
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_AT5T57  sky130_fd_pr__nfet_01v8_AT5T57_1
timestamp 1749624948
transform 1 0 938 0 1 58
box -73 -326 73 326
<< end >>
