magic
tech sky130A
magscale 1 2
timestamp 1751058216
<< error_p >>
rect 13380 13042 13548 13043
rect 13403 13030 13525 13036
rect 13414 13008 13514 13009
rect 13430 12992 13498 13008
rect 13176 12854 13198 12882
rect 13204 12826 13226 12910
rect 13176 12605 13198 12633
rect 13204 12577 13226 12661
rect 13176 12356 13198 12384
rect 13204 12346 13226 12412
use top_buffer_opamp  top_buffer_opamp_0
timestamp 1751058216
transform -1 0 -2156 0 1 9674
box -12462 -8798 520 13398
use top_seg_sel_interpolating  top_seg_sel_interpolating_0
timestamp 1751047404
transform 1 0 10818 0 -1 16090
box -418 2936 3076 6409
<< end >>
