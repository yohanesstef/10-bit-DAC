magic
tech sky130A
magscale 1 2
timestamp 1749835822
<< error_p >>
rect 9 2834 39 3322
rect 75 2900 105 3256
rect 1490 2900 1520 3256
rect 75 2896 391 2900
rect 451 2896 767 2900
rect 828 2896 1144 2900
rect 1204 2896 1520 2900
rect 1556 2834 1586 3322
rect 9 2830 1586 2834
rect 9 2226 1586 2230
rect 9 1873 39 2226
rect 75 2160 391 2164
rect 451 2160 767 2164
rect 828 2160 1144 2164
rect 1204 2160 1520 2164
rect 75 1873 105 2160
rect 1490 1873 1520 2160
rect 1556 1873 1586 2226
rect 9 1738 1586 1873
rect 39 1704 1556 1738
rect 9 1097 39 1585
rect 75 1163 105 1519
rect 1490 1163 1520 1519
rect 75 1159 391 1163
rect 451 1159 767 1163
rect 828 1159 1144 1163
rect 1204 1159 1520 1163
rect 1556 1097 1586 1585
rect 9 1093 1586 1097
rect 9 489 1586 493
rect 9 1 39 489
rect 75 423 391 427
rect 451 423 767 427
rect 828 423 1144 427
rect 1204 423 1520 427
rect 75 67 105 423
rect 1490 67 1520 423
rect 1556 1 1586 489
use cm_pcell1_4_4  cm_pcell1_4_4_0
timestamp 1749835822
transform 1 0 -1047 0 1 1348
box 1056 -1381 2633 2008
<< end >>
