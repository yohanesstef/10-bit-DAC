magic
tech sky130A
magscale 1 2
timestamp 1749550684
<< error_p >>
rect 37364 -7208 37370 -7202
rect 37418 -7208 37424 -7202
rect 37358 -7214 37364 -7208
rect 37424 -7214 37430 -7208
rect 37358 -7268 37364 -7262
rect 37424 -7268 37430 -7262
rect 37364 -7274 37370 -7268
rect 37418 -7274 37424 -7268
rect 37276 -7296 37282 -7290
rect 37330 -7296 37336 -7290
rect 37270 -7302 37276 -7296
rect 37336 -7302 37342 -7296
rect 37270 -7356 37276 -7350
rect 37336 -7356 37342 -7350
rect 37276 -7362 37282 -7356
rect 37330 -7362 37336 -7356
rect 37188 -7384 37194 -7378
rect 37242 -7384 37248 -7378
rect 37182 -7390 37188 -7384
rect 37248 -7390 37254 -7384
rect 37182 -7444 37188 -7438
rect 37248 -7444 37254 -7438
rect 37188 -7450 37194 -7444
rect 37242 -7450 37248 -7444
rect 37100 -7472 37106 -7466
rect 37154 -7472 37160 -7466
rect 37094 -7478 37100 -7472
rect 37160 -7478 37166 -7472
rect 37094 -7532 37100 -7526
rect 37160 -7532 37166 -7526
rect 37100 -7538 37106 -7532
rect 37154 -7538 37160 -7532
rect 33951 -7560 33957 -7554
rect 34005 -7560 34011 -7554
rect 33945 -7566 33951 -7560
rect 34011 -7566 34017 -7560
rect 33945 -7620 33951 -7614
rect 34011 -7620 34017 -7614
rect 33951 -7626 33957 -7620
rect 34005 -7626 34011 -7620
rect 33863 -7648 33869 -7642
rect 33917 -7648 33923 -7642
rect 33857 -7654 33863 -7648
rect 33923 -7654 33929 -7648
rect 33857 -7708 33863 -7702
rect 33923 -7708 33929 -7702
rect 33863 -7714 33869 -7708
rect 33917 -7714 33923 -7708
rect 33775 -7736 33781 -7730
rect 33829 -7736 33835 -7730
rect 33769 -7742 33775 -7736
rect 33835 -7742 33841 -7736
rect 33769 -7796 33775 -7790
rect 33835 -7796 33841 -7790
rect 33775 -7802 33781 -7796
rect 33829 -7802 33835 -7796
rect 33687 -7824 33693 -7818
rect 33741 -7824 33747 -7818
rect 33681 -7830 33687 -7824
rect 33747 -7830 33753 -7824
rect 33681 -7884 33687 -7878
rect 33747 -7884 33753 -7878
rect 33687 -7890 33693 -7884
rect 33741 -7890 33747 -7884
<< error_s >>
rect 40801 -5854 40807 -5848
rect 40855 -5854 40861 -5848
rect 40795 -5860 40801 -5854
rect 40861 -5860 40867 -5854
rect 40795 -5914 40801 -5908
rect 40861 -5914 40867 -5908
rect 40801 -5920 40807 -5914
rect 40855 -5920 40861 -5914
rect 40713 -5942 40719 -5936
rect 40767 -5942 40773 -5936
rect 40707 -5948 40713 -5942
rect 40773 -5948 40779 -5942
rect 40707 -6002 40713 -5996
rect 40773 -6002 40779 -5996
rect 40713 -6008 40719 -6002
rect 40767 -6008 40773 -6002
rect 40625 -6030 40631 -6024
rect 40679 -6030 40685 -6024
rect 40619 -6036 40625 -6030
rect 40685 -6036 40691 -6030
rect 40619 -6090 40625 -6084
rect 40685 -6090 40691 -6084
rect 40625 -6096 40631 -6090
rect 40679 -6096 40685 -6090
rect 40537 -6118 40543 -6112
rect 40591 -6118 40597 -6112
rect 40531 -6124 40537 -6118
rect 40597 -6124 40603 -6118
rect 40531 -6178 40537 -6172
rect 40597 -6178 40603 -6172
rect 40537 -6184 40543 -6178
rect 40591 -6184 40597 -6178
rect 40449 -6206 40455 -6200
rect 40503 -6206 40509 -6200
rect 40443 -6212 40449 -6206
rect 40509 -6212 40515 -6206
rect 40443 -6266 40449 -6260
rect 40509 -6266 40515 -6260
rect 40449 -6272 40455 -6266
rect 40503 -6272 40509 -6266
rect 40361 -6294 40367 -6288
rect 40415 -6294 40421 -6288
rect 40355 -6300 40361 -6294
rect 40421 -6300 40427 -6294
rect 40355 -6354 40361 -6348
rect 40421 -6354 40427 -6348
rect 40361 -6360 40367 -6354
rect 40415 -6360 40421 -6354
rect 40273 -6382 40279 -6376
rect 40327 -6382 40333 -6376
rect 40267 -6388 40273 -6382
rect 40333 -6388 40339 -6382
rect 40267 -6442 40273 -6436
rect 40333 -6442 40339 -6436
rect 40273 -6448 40279 -6442
rect 40327 -6448 40333 -6442
rect 40185 -6470 40191 -6464
rect 40239 -6470 40245 -6464
rect 40179 -6476 40185 -6470
rect 40245 -6476 40251 -6470
rect 40179 -6530 40185 -6524
rect 40245 -6530 40251 -6524
rect 40185 -6536 40191 -6530
rect 40239 -6536 40245 -6530
<< metal1 >>
rect 33687 -5474 34291 -5414
rect 36616 -5474 37424 -5414
rect 33687 -7824 33747 -5474
rect 33775 -5562 34291 -5502
rect 36293 -5562 37336 -5502
rect 33775 -7736 33835 -5562
rect 33863 -5650 34291 -5590
rect 36017 -5650 37248 -5590
rect 33863 -7648 33923 -5650
rect 33951 -5738 34291 -5678
rect 35741 -5738 37160 -5678
rect 33951 -7560 34011 -5738
rect 37100 -7472 37160 -5738
rect 37188 -7384 37248 -5650
rect 37276 -7296 37336 -5562
rect 37364 -7208 37424 -5474
rect 40185 -6470 40245 -5766
rect 40273 -6382 40333 -5766
rect 40361 -6294 40421 -5766
rect 40449 -6206 40509 -5766
rect 40537 -6118 40597 -5766
rect 40625 -6030 40685 -5766
rect 40713 -5942 40773 -5766
rect 40801 -5854 40861 -5766
rect 40801 -5920 40861 -5914
rect 40713 -6008 40773 -6002
rect 40625 -6096 40685 -6090
rect 40537 -6184 40597 -6178
rect 40449 -6272 40509 -6266
rect 40361 -6360 40421 -6354
rect 40273 -6448 40333 -6442
rect 40185 -6536 40245 -6530
rect 37364 -7274 37424 -7268
rect 37276 -7362 37336 -7356
rect 37188 -7450 37248 -7444
rect 37100 -7538 37160 -7532
rect 33951 -7626 34011 -7620
rect 33863 -7714 33923 -7708
rect 33775 -7802 33835 -7796
rect 33687 -7890 33747 -7884
<< via1 >>
rect 40801 -5914 40861 -5854
rect 40713 -6002 40773 -5942
rect 40625 -6090 40685 -6030
rect 40537 -6178 40597 -6118
rect 40449 -6266 40509 -6206
rect 40361 -6354 40421 -6294
rect 40273 -6442 40333 -6382
rect 40185 -6530 40245 -6470
rect 37364 -7268 37424 -7208
rect 37276 -7356 37336 -7296
rect 37188 -7444 37248 -7384
rect 37100 -7532 37160 -7472
rect 33951 -7620 34011 -7560
rect 33863 -7708 33923 -7648
rect 33775 -7796 33835 -7736
rect 33687 -7884 33747 -7824
<< metal2 >>
rect 36380 -4568 41629 -4508
rect 36104 -4656 41353 -4596
rect 35828 -4744 41077 -4684
rect 35562 -4832 40801 -4772
rect 35474 -4920 40317 -4860
rect 35208 -5008 40041 -4948
rect 34932 -5096 39765 -5036
rect 34656 -5184 39489 -5124
use nswitch_8_stage_1  nswitch_8_stage_1_0
timestamp 1749550684
transform 1 0 9756 0 1 2700
box 29523 -8466 32011 -7202
use nswitch_8_stage_2  nswitch_8_stage_2_0
timestamp 1749550684
transform 1 0 0 0 1 -88
box 34291 -5650 36817 -4414
<< end >>
