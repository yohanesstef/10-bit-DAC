magic
tech sky130A
magscale 1 2
timestamp 1750771847
<< mvpsubdiff >>
rect 1805 1933 4613 1993
rect 1805 1612 1865 1933
rect 4553 1612 4613 1933
rect 1805 1552 4613 1612
<< poly >>
rect 1876 1660 1936 1902
rect 4482 1660 4542 1902
<< locali >>
rect 4543 1980 4600 1981
rect 1818 1946 4600 1980
rect 1818 1599 1852 1946
rect 4566 1599 4600 1946
rect 1818 1565 4600 1599
rect 1818 1564 1875 1565
<< metal1 >>
rect 1795 1923 4623 2003
rect 1795 1622 1875 1923
rect 1957 1846 2310 1892
rect 1957 1814 2003 1846
rect 4415 1622 4461 1686
rect 4543 1622 4623 1923
rect 1795 1542 4623 1622
use sky130_fd_pr__nfet_g5v0d10v5_MLSP8N  sky130_fd_pr__nfet_g5v0d10v5_MLSP8N_0
timestamp 1750203240
transform 1 0 3209 0 1 1781
box -1258 -121 1258 121
<< end >>
