magic
tech sky130A
magscale 1 2
timestamp 1750863581
<< error_p >>
rect 8596 -1959 8602 -1953
rect 8654 -1959 8660 -1953
rect 12930 -1959 12936 -1953
rect 12984 -1959 12990 -1953
rect 8590 -1965 8596 -1959
rect 8660 -1965 8666 -1959
rect 12924 -1965 12930 -1959
rect 12990 -1965 12996 -1959
<< metal1 >>
rect 5748 -2019 8596 -1959
rect 8660 -2019 12930 -1959
rect 12990 -2019 23644 -1959
rect 5754 -2107 6030 -2047
rect 6094 -2107 13018 -2047
rect 13078 -2107 23644 -2047
rect 5754 -2195 8504 -2135
rect 8568 -2195 13574 -2135
rect 13634 -2195 23644 -2135
rect 5754 -2283 5938 -2223
rect 6002 -2283 13662 -2223
rect 13722 -2283 23644 -2223
rect 5754 -2371 8412 -2311
rect 8476 -2371 14218 -2311
rect 14278 -2371 23026 -2311
rect 23086 -2371 23644 -2311
rect 5754 -2459 5846 -2399
rect 5910 -2459 14306 -2399
rect 14366 -2459 23546 -2399
rect 23606 -2459 23644 -2399
rect 5754 -2547 8320 -2487
rect 8384 -2547 14862 -2487
rect 14922 -2547 20133 -2487
rect 20193 -2547 22938 -2487
rect 22998 -2547 23644 -2487
rect 5748 -2635 5754 -2575
rect 5818 -2635 14950 -2575
rect 15010 -2635 20317 -2575
rect 20377 -2635 23224 -2575
rect 23284 -2635 23644 -2575
rect 9226 -2723 15506 -2663
rect 15566 -2723 19143 -2663
rect 19203 -2723 21602 -2663
rect 21662 -2723 23644 -2663
rect 9226 -2811 15594 -2751
rect 15654 -2811 19327 -2751
rect 19387 -2811 22122 -2751
rect 22182 -2811 23644 -2751
rect 9226 -2899 16150 -2839
rect 16210 -2899 18153 -2839
rect 18213 -2899 21514 -2839
rect 21574 -2899 23644 -2839
rect 9226 -2987 16238 -2927
rect 16298 -2987 18337 -2927
rect 18397 -2987 21800 -2927
rect 21860 -2987 23644 -2927
rect 9226 -3075 16794 -3015
rect 16854 -3075 17163 -3015
rect 17223 -3075 23644 -3015
rect 9226 -3163 16882 -3103
rect 16942 -3163 17251 -3103
rect 17311 -3163 23644 -3103
rect 9226 -3251 15974 -3191
rect 16034 -3251 17438 -3191
rect 17498 -3251 23644 -3191
rect 9226 -3339 16414 -3279
rect 16474 -3339 17526 -3279
rect 17586 -3339 23644 -3279
rect 9226 -3427 15183 -3367
rect 15243 -3427 18082 -3367
rect 18142 -3427 23644 -3367
rect 9226 -3515 15367 -3455
rect 15427 -3515 18170 -3455
rect 18230 -3515 23644 -3455
rect 9226 -3603 14042 -3543
rect 14102 -3603 18726 -3543
rect 18786 -3603 23644 -3543
rect 9226 -3691 14482 -3631
rect 14542 -3691 18814 -3631
rect 18874 -3691 23644 -3631
rect 5366 -3807 24077 -3743
rect 5366 -3903 5386 -3807
rect 5542 -3903 8688 -3807
rect 8844 -3903 22539 -3807
rect 22635 -3903 23975 -3807
rect 24071 -3903 24077 -3807
rect 5564 -4447 5570 -4351
rect 5726 -4447 8872 -4351
rect 9028 -4447 20870 -4351
rect 21070 -4447 21235 -4351
rect 21331 -4447 25275 -4351
rect 25371 -4447 25377 -4351
rect 5564 -4551 25377 -4447
<< via1 >>
rect 8596 -2019 8660 -1959
rect 12930 -2019 12990 -1959
rect 6030 -2107 6094 -2047
rect 13018 -2107 13078 -2047
rect 8504 -2195 8568 -2135
rect 13574 -2195 13634 -2135
rect 5938 -2283 6002 -2223
rect 13662 -2283 13722 -2223
rect 8412 -2371 8476 -2311
rect 14218 -2371 14278 -2311
rect 23026 -2371 23086 -2311
rect 5846 -2459 5910 -2399
rect 14306 -2459 14366 -2399
rect 23546 -2459 23606 -2399
rect 8320 -2547 8384 -2487
rect 14862 -2547 14922 -2487
rect 20133 -2547 20193 -2487
rect 22938 -2547 22998 -2487
rect 5754 -2635 5818 -2575
rect 14950 -2635 15010 -2575
rect 20317 -2635 20377 -2575
rect 23224 -2635 23284 -2575
rect 15506 -2723 15566 -2663
rect 19143 -2723 19203 -2663
rect 21602 -2723 21662 -2663
rect 15594 -2811 15654 -2751
rect 19327 -2811 19387 -2751
rect 22122 -2811 22182 -2751
rect 16150 -2899 16210 -2839
rect 18153 -2899 18213 -2839
rect 21514 -2899 21574 -2839
rect 16238 -2987 16298 -2927
rect 18337 -2987 18397 -2927
rect 21800 -2987 21860 -2927
rect 16794 -3075 16854 -3015
rect 17163 -3075 17223 -3015
rect 16882 -3163 16942 -3103
rect 17251 -3163 17311 -3103
rect 15974 -3251 16034 -3191
rect 17438 -3251 17498 -3191
rect 16414 -3339 16474 -3279
rect 17526 -3339 17586 -3279
rect 15183 -3427 15243 -3367
rect 18082 -3427 18142 -3367
rect 15367 -3515 15427 -3455
rect 18170 -3515 18230 -3455
rect 14042 -3603 14102 -3543
rect 18726 -3603 18786 -3543
rect 14482 -3691 14542 -3631
rect 18814 -3691 18874 -3631
rect 5386 -3903 5542 -3807
rect 8688 -3903 8844 -3807
rect 22539 -3903 22635 -3807
rect 23975 -3903 24071 -3807
rect 5570 -4447 5726 -4351
rect 8872 -4447 9028 -4351
rect 20870 -4447 21070 -4351
rect 21235 -4447 21331 -4351
rect 25275 -4447 25371 -4351
<< metal2 >>
rect 5386 -3807 5542 -1959
rect 5386 -3909 5542 -3903
rect 5570 -4351 5726 -1959
rect 5754 -2575 5818 -1959
rect 5846 -2399 5910 -1959
rect 5938 -2223 6002 -1959
rect 6030 -2047 6094 -1959
rect 6030 -2113 6094 -2107
rect 5938 -2289 6002 -2283
rect 5846 -2465 5910 -2459
rect 8320 -2487 8384 -1959
rect 8412 -2311 8476 -1959
rect 8504 -2135 8568 -1959
rect 8596 -2025 8660 -2019
rect 8504 -2201 8568 -2195
rect 8412 -2377 8476 -2371
rect 8320 -2553 8384 -2547
rect 5754 -2641 5818 -2635
rect 8688 -3807 8844 -1959
rect 8688 -3909 8844 -3903
rect 5570 -4453 5726 -4447
rect 8872 -4351 9028 -1959
rect 12930 -3807 12990 -2019
rect 13018 -2047 13078 -2041
rect 13018 -3807 13078 -2107
rect 13574 -2135 13634 -2129
rect 13574 -3807 13634 -2195
rect 13662 -2223 13722 -2217
rect 13662 -3807 13722 -2283
rect 14042 -3543 14102 -1959
rect 14042 -3609 14102 -3603
rect 14218 -2311 14278 -2305
rect 14218 -3807 14278 -2371
rect 14306 -2399 14366 -2393
rect 14306 -3807 14366 -2459
rect 14482 -3631 14542 -1959
rect 14482 -3697 14542 -3691
rect 14862 -2487 14922 -2481
rect 14862 -3807 14922 -2547
rect 14950 -2575 15010 -2569
rect 14950 -3807 15010 -2635
rect 15183 -3367 15243 -1959
rect 15183 -3433 15243 -3427
rect 15367 -3455 15427 -1959
rect 15367 -3521 15427 -3515
rect 15506 -2663 15566 -2657
rect 15506 -3807 15566 -2723
rect 15594 -2751 15654 -2745
rect 15594 -3807 15654 -2811
rect 15974 -3191 16034 -1959
rect 15974 -3257 16034 -3251
rect 16150 -2839 16210 -2833
rect 16150 -3807 16210 -2899
rect 16238 -2927 16298 -2921
rect 16238 -3807 16298 -2987
rect 16414 -3279 16474 -1959
rect 16414 -3345 16474 -3339
rect 16794 -3015 16854 -3009
rect 16794 -3807 16854 -3075
rect 17163 -3015 17223 -1959
rect 17163 -3081 17223 -3075
rect 16882 -3103 16942 -3097
rect 16882 -3807 16942 -3163
rect 17251 -3103 17311 -1959
rect 18153 -2839 18213 -1959
rect 18153 -2905 18213 -2899
rect 18337 -2927 18397 -1959
rect 19143 -2663 19203 -1959
rect 19143 -2729 19203 -2723
rect 19327 -2751 19387 -1959
rect 20133 -2487 20193 -1959
rect 20133 -2553 20193 -2547
rect 20317 -2575 20377 -1959
rect 20317 -2641 20377 -2635
rect 19327 -2817 19387 -2811
rect 18337 -2993 18397 -2987
rect 17251 -3169 17311 -3163
rect 17438 -3191 17498 -3185
rect 17438 -3807 17498 -3251
rect 17526 -3279 17586 -3273
rect 17526 -3807 17586 -3339
rect 18082 -3367 18142 -3361
rect 18082 -3807 18142 -3427
rect 18170 -3455 18230 -3449
rect 18170 -3807 18230 -3515
rect 18726 -3543 18786 -3537
rect 18726 -3807 18786 -3603
rect 18814 -3631 18874 -3625
rect 18814 -3807 18874 -3691
rect 20870 -4351 21070 -1959
rect 13309 -4447 13369 -4387
rect 13953 -4447 14013 -4387
rect 14597 -4447 14657 -4387
rect 15241 -4447 15301 -4387
rect 15885 -4447 15945 -4387
rect 16529 -4447 16589 -4387
rect 17173 -4447 17233 -4387
rect 17817 -4447 17877 -4387
rect 18461 -4447 18521 -4387
rect 8872 -4453 9028 -4447
rect 20870 -4453 21070 -4447
rect 21235 -4351 21331 -1959
rect 21514 -2839 21574 -1959
rect 21602 -2663 21662 -1959
rect 21602 -2729 21662 -2723
rect 21514 -2905 21574 -2899
rect 21800 -2927 21860 -1959
rect 22122 -2751 22182 -1959
rect 22122 -2817 22182 -2811
rect 21800 -2993 21860 -2987
rect 22539 -3807 22635 -1959
rect 22938 -2487 22998 -1959
rect 23026 -2311 23086 -1959
rect 23026 -2377 23086 -2371
rect 22938 -2553 22998 -2547
rect 23224 -2575 23284 -1959
rect 23546 -2399 23606 -1959
rect 23546 -2465 23606 -2459
rect 23224 -2641 23284 -2635
rect 22539 -3909 22635 -3903
rect 23975 -3807 24071 -1959
rect 23975 -3909 24071 -3903
rect 21235 -4453 21331 -4447
rect 25275 -4351 25371 -1959
rect 25275 -4453 25371 -4447
use buffer_bus  buffer_bus_0
timestamp 1750863581
transform 1 0 11354 0 1 4262
box 1252 -8709 7768 -8069
<< labels >>
flabel metal2 s 18461 -4447 18521 -4387 0 FreeSans 160 180 0 0 DIN0
port 0 nsew
flabel metal2 s 17817 -4447 17877 -4387 0 FreeSans 160 180 0 0 DIN1
port 1 nsew
flabel metal2 s 17173 -4447 17233 -4387 0 FreeSans 160 180 0 0 DIN2
port 2 nsew
flabel metal2 s 16529 -4447 16589 -4387 0 FreeSans 160 180 0 0 DIN3
port 3 nsew
flabel metal2 s 15885 -4447 15945 -4387 0 FreeSans 160 180 0 0 DIN4
port 4 nsew
flabel metal2 s 15241 -4447 15301 -4387 0 FreeSans 160 180 0 0 DIN5
port 5 nsew
flabel metal2 s 14597 -4447 14657 -4387 0 FreeSans 160 180 0 0 DIN6
port 6 nsew
flabel metal2 s 13953 -4447 14013 -4387 0 FreeSans 160 180 0 0 DIN7
port 7 nsew
flabel metal2 s 13309 -4447 13369 -4387 0 FreeSans 160 180 0 0 DIN8
port 8 nsew
flabel metal2 s 18814 -3807 18874 -3747 0 FreeSans 160 0 0 0 D[0]
port 10 nsew
flabel metal2 s 18170 -3807 18230 -3747 0 FreeSans 160 0 0 0 D[1]
port 11 nsew
flabel metal2 s 17526 -3807 17586 -3747 0 FreeSans 160 0 0 0 D[2]
port 12 nsew
flabel metal2 s 16882 -3807 16942 -3747 0 FreeSans 160 0 0 0 D[3]
port 13 nsew
flabel metal2 s 16238 -3807 16298 -3747 0 FreeSans 160 0 0 0 D[4]
port 14 nsew
flabel metal2 s 15594 -3807 15654 -3747 0 FreeSans 160 0 0 0 D[5]
port 15 nsew
flabel metal2 s 14950 -3807 15010 -3747 0 FreeSans 160 0 0 0 D[6]
port 16 nsew
flabel metal2 s 14306 -3807 14366 -3747 0 FreeSans 160 0 0 0 D[7]
port 17 nsew
flabel metal2 s 13662 -3807 13722 -3747 0 FreeSans 160 0 0 0 D[8]
port 18 nsew
flabel metal2 s 13018 -3807 13078 -3747 0 FreeSans 160 0 0 0 D[9]
port 19 nsew
flabel metal2 s 18726 -3807 18786 -3747 0 FreeSans 160 180 0 0 DB[0]
port 20 nsew
flabel metal2 s 18082 -3807 18142 -3747 0 FreeSans 160 180 0 0 DB[1]
port 21 nsew
flabel metal2 s 17438 -3807 17498 -3747 0 FreeSans 160 180 0 0 DB[2]
port 22 nsew
flabel metal2 s 16794 -3807 16854 -3747 0 FreeSans 160 180 0 0 DB[3]
port 23 nsew
flabel metal2 s 16150 -3807 16210 -3747 0 FreeSans 160 180 0 0 DB[4]
port 24 nsew
flabel metal2 s 15506 -3807 15566 -3747 0 FreeSans 160 180 0 0 DB[5]
port 25 nsew
flabel metal2 s 14862 -3807 14922 -3747 0 FreeSans 160 180 0 0 DB[6]
port 26 nsew
flabel metal2 s 14218 -3807 14278 -3747 0 FreeSans 160 180 0 0 DB[7]
port 27 nsew
flabel metal2 s 13574 -3807 13634 -3747 0 FreeSans 160 180 0 0 DB[8]
port 28 nsew
flabel metal2 s 12930 -3807 12990 -3747 0 FreeSans 160 180 0 0 DB[9]
port 29 nsew
flabel metal1 s 12584 -3903 12644 -3843 0 FreeSans 160 0 0 0 VDD
port 30 nsew
flabel metal1 s 12573 -4411 12633 -4351 0 FreeSans 160 0 0 0 GND
port 31 nsew
flabel metal2 s 12665 -4447 12725 -4387 0 FreeSans 160 0 0 0 DIN9
port 9 nsew
<< end >>
