magic
tech sky130A
magscale 1 2
timestamp 1750828667
<< metal1 >>
rect 981 6 1041 941
rect 1971 52 2031 987
rect 2961 52 3021 987
use lvsf_inv  lvsf_inv_0
timestamp 1750828667
transform 1 0 -56 0 1 -17
box 11 3 1133 2956
use lvsf_inv  lvsf_inv_1
timestamp 1750828667
transform 1 0 934 0 1 -17
box 11 3 1133 2956
use lvsf_inv  lvsf_inv_2
timestamp 1750828667
transform 1 0 1924 0 1 -17
box 11 3 1133 2956
use lvsf_inv  lvsf_inv_3
timestamp 1750828667
transform 1 0 2914 0 1 -17
box 11 3 1133 2956
<< end >>
