magic
tech sky130A
magscale 1 2
timestamp 1751045931
<< error_p >>
rect -223 570 223 604
rect -253 355 253 570
rect -223 321 223 355
rect -253 106 253 321
rect -223 72 223 106
rect -253 -143 253 72
rect -223 -177 223 -143
rect -253 -392 253 -177
rect -253 -638 -223 -426
rect -187 -572 -157 -492
rect 157 -572 187 -492
rect -187 -576 187 -572
rect 223 -638 253 -426
rect -253 -642 253 -638
<< nwell >>
rect -223 358 223 604
rect -223 109 223 355
rect -223 -140 223 106
rect -223 -389 223 -143
rect -223 -638 223 -392
<< mvpmos >>
rect -129 420 -29 504
rect 29 420 129 504
rect -129 171 -29 255
rect 29 171 129 255
rect -129 -78 -29 6
rect 29 -78 129 6
rect -129 -327 -29 -243
rect 29 -327 129 -243
rect -129 -576 -29 -492
rect 29 -576 129 -492
<< mvpdiff >>
rect -187 492 -129 504
rect -187 432 -175 492
rect -141 432 -129 492
rect -187 420 -129 432
rect -29 492 29 504
rect -29 432 -17 492
rect 17 432 29 492
rect -29 420 29 432
rect 129 492 187 504
rect 129 432 141 492
rect 175 432 187 492
rect 129 420 187 432
rect -187 243 -129 255
rect -187 183 -175 243
rect -141 183 -129 243
rect -187 171 -129 183
rect -29 243 29 255
rect -29 183 -17 243
rect 17 183 29 243
rect -29 171 29 183
rect 129 243 187 255
rect 129 183 141 243
rect 175 183 187 243
rect 129 171 187 183
rect -187 -6 -129 6
rect -187 -66 -175 -6
rect -141 -66 -129 -6
rect -187 -78 -129 -66
rect -29 -6 29 6
rect -29 -66 -17 -6
rect 17 -66 29 -6
rect -29 -78 29 -66
rect 129 -6 187 6
rect 129 -66 141 -6
rect 175 -66 187 -6
rect 129 -78 187 -66
rect -187 -255 -129 -243
rect -187 -315 -175 -255
rect -141 -315 -129 -255
rect -187 -327 -129 -315
rect -29 -255 29 -243
rect -29 -315 -17 -255
rect 17 -315 29 -255
rect -29 -327 29 -315
rect 129 -255 187 -243
rect 129 -315 141 -255
rect 175 -315 187 -255
rect 129 -327 187 -315
rect -187 -504 -129 -492
rect -187 -564 -175 -504
rect -141 -564 -129 -504
rect -187 -576 -129 -564
rect -29 -504 29 -492
rect -29 -564 -17 -504
rect 17 -564 29 -504
rect -29 -576 29 -564
rect 129 -504 187 -492
rect 129 -564 141 -504
rect 175 -564 187 -504
rect 129 -576 187 -564
<< mvpdiffc >>
rect -175 432 -141 492
rect -17 432 17 492
rect 141 432 175 492
rect -175 183 -141 243
rect -17 183 17 243
rect 141 183 175 243
rect -175 -66 -141 -6
rect -17 -66 17 -6
rect 141 -66 175 -6
rect -175 -315 -141 -255
rect -17 -315 17 -255
rect 141 -315 175 -255
rect -175 -564 -141 -504
rect -17 -564 17 -504
rect 141 -564 175 -504
<< poly >>
rect -129 585 -29 601
rect -129 551 -113 585
rect -45 551 -29 585
rect -129 504 -29 551
rect 29 585 129 601
rect 29 551 45 585
rect 113 551 129 585
rect 29 504 129 551
rect -129 394 -29 420
rect 29 394 129 420
rect -129 336 -29 352
rect -129 302 -113 336
rect -45 302 -29 336
rect -129 255 -29 302
rect 29 336 129 352
rect 29 302 45 336
rect 113 302 129 336
rect 29 255 129 302
rect -129 145 -29 171
rect 29 145 129 171
rect -129 87 -29 103
rect -129 53 -113 87
rect -45 53 -29 87
rect -129 6 -29 53
rect 29 87 129 103
rect 29 53 45 87
rect 113 53 129 87
rect 29 6 129 53
rect -129 -104 -29 -78
rect 29 -104 129 -78
rect -129 -162 -29 -146
rect -129 -196 -113 -162
rect -45 -196 -29 -162
rect -129 -243 -29 -196
rect 29 -162 129 -146
rect 29 -196 45 -162
rect 113 -196 129 -162
rect 29 -243 129 -196
rect -129 -353 -29 -327
rect 29 -353 129 -327
rect -129 -411 -29 -395
rect -129 -445 -113 -411
rect -45 -445 -29 -411
rect -129 -492 -29 -445
rect 29 -411 129 -395
rect 29 -445 45 -411
rect 113 -445 129 -411
rect 29 -492 129 -445
rect -129 -602 -29 -576
rect 29 -602 129 -576
<< polycont >>
rect -113 551 -45 585
rect 45 551 113 585
rect -113 302 -45 336
rect 45 302 113 336
rect -113 53 -45 87
rect 45 53 113 87
rect -113 -196 -45 -162
rect 45 -196 113 -162
rect -113 -445 -45 -411
rect 45 -445 113 -411
<< locali >>
rect -129 551 -113 585
rect -45 551 -29 585
rect 29 551 45 585
rect 113 551 129 585
rect -175 492 -141 508
rect -175 416 -141 432
rect -17 492 17 508
rect -17 416 17 432
rect 141 492 175 508
rect 141 416 175 432
rect -129 302 -113 336
rect -45 302 -29 336
rect 29 302 45 336
rect 113 302 129 336
rect -175 243 -141 259
rect -175 167 -141 183
rect -17 243 17 259
rect -17 167 17 183
rect 141 243 175 259
rect 141 167 175 183
rect -129 53 -113 87
rect -45 53 -29 87
rect 29 53 45 87
rect 113 53 129 87
rect -175 -6 -141 10
rect -175 -82 -141 -66
rect -17 -6 17 10
rect -17 -82 17 -66
rect 141 -6 175 10
rect 141 -82 175 -66
rect -129 -196 -113 -162
rect -45 -196 -29 -162
rect 29 -196 45 -162
rect 113 -196 129 -162
rect -175 -255 -141 -239
rect -175 -331 -141 -315
rect -17 -255 17 -239
rect -17 -331 17 -315
rect 141 -255 175 -239
rect 141 -331 175 -315
rect -129 -445 -113 -411
rect -45 -445 -29 -411
rect 29 -445 45 -411
rect 113 -445 129 -411
rect -175 -504 -141 -488
rect -175 -580 -141 -564
rect -17 -504 17 -488
rect -17 -580 17 -564
rect 141 -504 175 -488
rect 141 -580 175 -564
<< viali >>
rect -105 551 -53 585
rect 53 551 105 585
rect -175 432 -141 492
rect -17 432 17 492
rect 141 432 175 492
rect -105 302 -53 336
rect 53 302 105 336
rect -175 183 -141 243
rect -17 183 17 243
rect 141 183 175 243
rect -105 53 -53 87
rect 53 53 105 87
rect -175 -66 -141 -6
rect -17 -66 17 -6
rect 141 -66 175 -6
rect -105 -196 -53 -162
rect 53 -196 105 -162
rect -175 -315 -141 -255
rect -17 -315 17 -255
rect 141 -315 175 -255
rect -105 -445 -53 -411
rect 53 -445 105 -411
rect -175 -564 -141 -504
rect -17 -564 17 -504
rect 141 -564 175 -504
<< metal1 >>
rect -117 585 -41 591
rect -117 551 -105 585
rect -53 551 -41 585
rect -117 545 -41 551
rect 41 585 117 591
rect 41 551 53 585
rect 105 551 117 585
rect 41 545 117 551
rect -181 492 -135 504
rect -181 432 -175 492
rect -141 432 -135 492
rect -181 420 -135 432
rect -23 492 23 504
rect -23 432 -17 492
rect 17 432 23 492
rect -23 420 23 432
rect 135 492 181 504
rect 135 432 141 492
rect 175 432 181 492
rect 135 420 181 432
rect -117 336 -41 342
rect -117 302 -105 336
rect -53 302 -41 336
rect -117 296 -41 302
rect 41 336 117 342
rect 41 302 53 336
rect 105 302 117 336
rect 41 296 117 302
rect -181 243 -135 255
rect -181 183 -175 243
rect -141 183 -135 243
rect -181 171 -135 183
rect -23 243 23 255
rect -23 183 -17 243
rect 17 183 23 243
rect -23 171 23 183
rect 135 243 181 255
rect 135 183 141 243
rect 175 183 181 243
rect 135 171 181 183
rect -117 87 -41 93
rect -117 53 -105 87
rect -53 53 -41 87
rect -117 47 -41 53
rect 41 87 117 93
rect 41 53 53 87
rect 105 53 117 87
rect 41 47 117 53
rect -181 -6 -135 6
rect -181 -66 -175 -6
rect -141 -66 -135 -6
rect -181 -78 -135 -66
rect -23 -6 23 6
rect -23 -66 -17 -6
rect 17 -66 23 -6
rect -23 -78 23 -66
rect 135 -6 181 6
rect 135 -66 141 -6
rect 175 -66 181 -6
rect 135 -78 181 -66
rect -117 -162 -41 -156
rect -117 -196 -105 -162
rect -53 -196 -41 -162
rect -117 -202 -41 -196
rect 41 -162 117 -156
rect 41 -196 53 -162
rect 105 -196 117 -162
rect 41 -202 117 -196
rect -181 -255 -135 -243
rect -181 -315 -175 -255
rect -141 -315 -135 -255
rect -181 -327 -135 -315
rect -23 -255 23 -243
rect -23 -315 -17 -255
rect 17 -315 23 -255
rect -23 -327 23 -315
rect 135 -255 181 -243
rect 135 -315 141 -255
rect 175 -315 181 -255
rect 135 -327 181 -315
rect -117 -411 -41 -405
rect -117 -445 -105 -411
rect -53 -445 -41 -411
rect -117 -451 -41 -445
rect 41 -411 117 -405
rect 41 -445 53 -411
rect 105 -445 117 -411
rect 41 -451 117 -445
rect -181 -504 -135 -492
rect -181 -564 -175 -504
rect -141 -564 -135 -504
rect -181 -576 -135 -564
rect -23 -504 23 -492
rect -23 -564 -17 -504
rect 17 -564 23 -504
rect -23 -576 23 -564
rect 135 -504 181 -492
rect 135 -564 141 -504
rect 175 -564 181 -504
rect 135 -576 181 -564
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.42 l 0.50 m 5 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
