magic
tech sky130A
magscale 1 2
timestamp 1749908815
<< metal1 >>
tri 36271 2000 36306 2035 se
rect 36306 2000 36393 2035
tri 36186 1915 36271 2000 se
rect 36271 1975 36393 2000
tri 36271 1915 36331 1975 nw
rect 36114 1855 36120 1915
rect 36180 1855 36211 1915
tri 36211 1855 36271 1915 nw
rect 36331 1855 36420 1915
tri 38153 1316 40154 3317 se
rect 40154 1817 40812 3317
rect 40154 1316 40274 1817
rect 38153 1315 40274 1316
tri 40274 1315 40776 1817 nw
rect 38153 -185 38774 1315
tri 38774 -185 40274 1315 nw
<< end >>
