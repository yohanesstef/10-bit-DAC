magic
tech sky130A
magscale 1 2
timestamp 1750202961
<< mvpsubdiff >>
rect 1805 1927 4153 1987
rect 1805 1612 1865 1927
rect 4093 1612 4153 1927
rect 1805 1552 4153 1612
<< poly >>
rect 1876 1660 1936 1896
rect 4022 1660 4082 1896
<< locali >>
rect 4083 1974 4140 1975
rect 1818 1940 4140 1974
rect 1818 1599 1852 1940
rect 4106 1599 4140 1940
rect 1818 1565 4140 1599
rect 1818 1564 1875 1565
<< metal1 >>
rect 1795 1917 4163 1997
rect 1795 1622 1875 1917
rect 3955 1622 4001 1686
rect 4083 1622 4163 1917
rect 1795 1542 4163 1622
use sky130_fd_pr__nfet_g5v0d10v5_TNA5KF  sky130_fd_pr__nfet_g5v0d10v5_TNA5KF_0
timestamp 1750202961
transform 1 0 2979 0 1 1778
box -1028 -118 1028 118
<< end >>
