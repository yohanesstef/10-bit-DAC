magic
tech sky130A
magscale 1 2
timestamp 1749643209
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_0
timestamp 1749643209
transform 1 0 1339 0 1 -1603
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_1
timestamp 1749643209
transform 1 0 1427 0 1 -1603
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_2
timestamp 1749643209
transform 1 0 1515 0 1 -1603
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_3
timestamp 1749643209
transform 1 0 1603 0 1 -1603
box -73 -226 73 226
<< end >>
