magic
tech sky130A
magscale 1 2
timestamp 1749563217
<< metal1 >>
rect 1540 -22764 1600 -22615
rect 1628 -22764 1688 -22615
rect 1716 -22764 1776 -22615
rect 1804 -22764 1864 -22615
rect 1892 -22764 1952 -22615
<< end >>
