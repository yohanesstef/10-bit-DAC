magic
tech sky130A
magscale 1 2
timestamp 1751017459
<< metal1 >>
rect 12 14552 9288 14609
rect 12 -16 7032 28
<< via1 >>
rect 112 14694 172 14754
rect 110 -183 170 -123
rect 7191 -401 7313 -345
<< metal2 >>
rect 102 17064 238 17066
rect 102 17008 111 17064
rect 233 17008 238 17064
rect 102 17006 238 17008
rect 4927 15281 5243 15283
rect 4927 15225 5177 15281
rect 5233 15225 5243 15281
rect 4927 15223 5243 15225
rect 104 14694 112 14754
rect 172 14694 180 14754
rect 5167 11962 5177 12018
rect 5233 11962 5243 12018
rect 104 11930 1218 11932
rect 104 11874 114 11930
rect 170 11874 1218 11930
rect 104 11872 1218 11874
rect 8058 11842 9137 11844
rect 8058 11786 9005 11842
rect 9127 11786 9137 11842
rect 8058 11784 9137 11786
rect 5167 10818 5177 10874
rect 5233 10818 5243 10874
rect 5167 10271 5177 10327
rect 5233 10271 5243 10327
rect 7306 9358 9137 9360
rect 7306 9302 9005 9358
rect 9127 9302 9137 9358
rect 7306 9300 9137 9302
rect 104 9270 1970 9272
rect 104 9214 114 9270
rect 170 9214 1970 9270
rect 104 9212 1970 9214
rect 5167 9127 5177 9183
rect 5233 9127 5243 9183
rect 4622 4599 4632 4655
rect 4688 4599 4698 4655
rect 4622 3983 4632 4039
rect 4688 3983 4698 4039
rect 4622 3083 4632 3139
rect 4688 3083 4698 3139
rect 4622 2466 4632 2522
rect 4688 2466 4698 2522
rect 102 1797 514 1800
rect 102 1741 112 1797
rect 168 1741 514 1797
rect 102 1739 514 1741
rect 102 1357 514 1360
rect 102 1301 112 1357
rect 168 1301 514 1357
rect 102 1299 514 1301
rect 102 809 514 812
rect 102 753 112 809
rect 168 753 514 809
rect 102 751 514 753
rect 102 369 514 372
rect 102 313 112 369
rect 168 313 514 369
rect 102 311 514 313
rect 102 -183 110 -123
rect 170 -183 178 -123
rect 4428 -257 4893 -255
rect 4428 -313 4632 -257
rect 4688 -313 4893 -257
rect 4428 -315 4893 -313
rect 7181 -401 7191 -345
rect 7313 -401 7323 -345
rect 4428 -553 4893 -551
rect 4428 -609 4632 -553
rect 4688 -609 4893 -553
rect 4428 -611 4893 -609
<< via2 >>
rect 111 17008 233 17064
rect 5177 15225 5233 15281
rect 114 14697 170 14753
rect 5177 11962 5233 12018
rect 114 11874 170 11930
rect 9005 11786 9127 11842
rect 5177 10818 5233 10874
rect 5177 10271 5233 10327
rect 9005 9302 9127 9358
rect 114 9214 170 9270
rect 5177 9127 5233 9183
rect 4632 4599 4688 4655
rect 4632 3983 4688 4039
rect 4632 3082 4688 3138
rect 4632 2466 4688 2522
rect 112 1741 168 1797
rect 112 1301 168 1357
rect 112 753 168 809
rect 112 313 168 369
rect 112 -180 168 -124
rect 4632 -313 4688 -257
rect 7191 -401 7313 -345
rect 4632 -609 4688 -553
<< metal3 >>
rect 106 17064 238 17204
rect 106 17008 111 17064
rect 233 17008 238 17064
rect 106 16999 238 17008
rect 5172 15281 5238 15286
rect 5172 15225 5177 15281
rect 5233 15225 5238 15281
rect 109 14753 175 14763
rect 109 14697 114 14753
rect 170 14697 175 14753
rect 109 11930 175 14697
rect 109 11874 114 11930
rect 170 11874 175 11930
rect 109 9270 175 11874
rect 109 9214 114 9270
rect 170 9214 175 9270
rect 109 9204 175 9214
rect 5172 12018 5238 15225
rect 5172 11962 5177 12018
rect 5233 11962 5238 12018
rect 5172 10874 5238 11962
rect 5172 10818 5177 10874
rect 5233 10818 5238 10874
rect 5172 10327 5238 10818
rect 5172 10271 5177 10327
rect 5233 10271 5238 10327
rect 5172 9183 5238 10271
rect 5172 9127 5177 9183
rect 5233 9127 5238 9183
rect 5172 9117 5238 9127
rect 9000 11842 9132 11852
rect 9000 11786 9005 11842
rect 9127 11786 9132 11842
rect 9000 9358 9132 11786
rect 9000 9302 9005 9358
rect 9127 9302 9132 9358
rect 9000 5006 9132 9302
rect 7186 4874 9132 5006
rect 4627 4655 4693 4665
rect 4627 4599 4632 4655
rect 4688 4599 4693 4655
rect 4627 4039 4693 4599
rect 4627 3983 4632 4039
rect 4688 3983 4693 4039
rect 4627 3138 4693 3983
rect 4627 3082 4632 3138
rect 4688 3082 4693 3138
rect 4627 2522 4693 3082
rect 4627 2466 4632 2522
rect 4688 2466 4693 2522
rect 107 1797 173 1807
rect 107 1741 112 1797
rect 168 1741 173 1797
rect 107 1357 173 1741
rect 107 1301 112 1357
rect 168 1301 173 1357
rect 107 809 173 1301
rect 107 753 112 809
rect 168 753 173 809
rect 107 369 173 753
rect 107 313 112 369
rect 168 313 173 369
rect 107 -124 173 313
rect 107 -180 112 -124
rect 168 -180 173 -124
rect 107 -190 173 -180
rect 4627 -257 4693 2466
rect 4627 -313 4632 -257
rect 4688 -313 4693 -257
rect 4627 -553 4693 -313
rect 7186 -345 7318 4874
rect 7186 -401 7191 -345
rect 7313 -401 7318 -345
rect 7186 -411 7318 -401
rect 4627 -609 4632 -553
rect 4688 -609 4693 -553
rect 4627 -619 4693 -609
use cm_ncell3  cm_ncell3_0
timestamp 1750150351
transform -1 0 9275 0 -1 -435
box -60 -455 9289 451
use cm_pcell3  cm_pcell3_0
timestamp 1750156376
transform 1 0 4623 0 -1 28738
box -4665 11508 4744 14208
use opa_input_stage  opa_input_stage_0
timestamp 1751017459
transform 1 0 -14 0 1 5133
box -30 -5131 9334 9476
<< end >>
