magic
tech sky130A
magscale 1 2
timestamp 1749664768
<< error_s >>
rect 41113 -4070 41119 -4064
rect 41167 -4070 41173 -4064
rect 41107 -4076 41113 -4070
rect 41173 -4076 41179 -4070
rect 41107 -4130 41113 -4124
rect 41173 -4130 41179 -4124
rect 41113 -4136 41119 -4130
rect 41167 -4136 41173 -4130
rect 40837 -4158 40843 -4152
rect 40891 -4158 40897 -4152
rect 40831 -4164 40837 -4158
rect 40897 -4164 40903 -4158
rect 40831 -4218 40837 -4212
rect 40897 -4218 40903 -4212
rect 40837 -4224 40843 -4218
rect 40891 -4224 40897 -4218
rect 40561 -4246 40567 -4240
rect 40615 -4246 40621 -4240
rect 40555 -4252 40561 -4246
rect 40621 -4252 40627 -4246
rect 40555 -4306 40561 -4300
rect 40621 -4306 40627 -4300
rect 40561 -4312 40567 -4306
rect 40615 -4312 40621 -4306
rect 40285 -4334 40291 -4328
rect 40339 -4334 40345 -4328
rect 40279 -4340 40285 -4334
rect 40345 -4340 40351 -4334
rect 40279 -4394 40285 -4388
rect 40345 -4394 40351 -4388
rect 40285 -4400 40291 -4394
rect 40339 -4400 40345 -4394
rect 39981 -4422 39987 -4416
rect 40035 -4422 40041 -4416
rect 39975 -4428 39981 -4422
rect 40041 -4428 40047 -4422
rect 39975 -4482 39981 -4476
rect 40041 -4482 40047 -4476
rect 39981 -4488 39987 -4482
rect 40035 -4488 40041 -4482
rect 39705 -4510 39711 -4504
rect 39759 -4510 39765 -4504
rect 39699 -4516 39705 -4510
rect 39765 -4516 39771 -4510
rect 39699 -4570 39705 -4564
rect 39765 -4570 39771 -4564
rect 39705 -4576 39711 -4570
rect 39759 -4576 39765 -4570
rect 39429 -4598 39435 -4592
rect 39483 -4598 39489 -4592
rect 39423 -4604 39429 -4598
rect 39489 -4604 39495 -4598
rect 39423 -4658 39429 -4652
rect 39489 -4658 39495 -4652
rect 39429 -4664 39435 -4658
rect 39483 -4664 39489 -4658
rect 39153 -4686 39159 -4680
rect 39207 -4686 39213 -4680
rect 39147 -4692 39153 -4686
rect 39213 -4692 39219 -4686
rect 39147 -4746 39153 -4740
rect 39213 -4746 39219 -4740
rect 39153 -4752 39159 -4746
rect 39207 -4752 39213 -4746
<< nwell >>
rect 37186 -4181 41530 -3573
<< mvnsubdiff >>
rect 37252 -3651 41464 -3639
rect 37252 -3685 37360 -3651
rect 41356 -3685 41464 -3651
rect 37252 -3697 41464 -3685
rect 37252 -3747 37310 -3697
rect 37252 -4007 37264 -3747
rect 37298 -4007 37310 -3747
rect 37252 -4057 37310 -4007
rect 41406 -3747 41464 -3697
rect 41406 -4007 41418 -3747
rect 41452 -4007 41464 -3747
rect 41406 -4057 41464 -4007
rect 37252 -4069 41464 -4057
rect 37252 -4103 37360 -4069
rect 41356 -4103 41464 -4069
rect 37252 -4115 41464 -4103
<< mvnsubdiffcont >>
rect 37360 -3685 41356 -3651
rect 37264 -4007 37298 -3747
rect 41418 -4007 41452 -3747
rect 37360 -4103 41356 -4069
<< locali >>
rect 37264 -3685 37360 -3651
rect 41356 -3685 41452 -3651
rect 37264 -3747 37298 -3685
rect 37264 -4069 37298 -4007
rect 41418 -3747 41452 -3685
rect 41418 -4069 41452 -4007
rect 37264 -4103 37360 -4069
rect 41356 -4103 41452 -4069
use pswitch_16_final  pswitch_16_final_0
timestamp 1749664768
transform 1 0 2216 0 1 526
box 34970 -5278 39314 -3861
<< end >>
