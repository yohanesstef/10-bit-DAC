magic
tech sky130A
magscale 1 2
timestamp 1749567216
<< error_p >>
rect 3213 1590 3215 1596
rect 3213 1536 3215 1542
<< error_s >>
rect 4317 1448 4323 1454
rect 4383 1448 4389 1454
rect 4323 1442 4329 1448
rect 4377 1442 4383 1448
rect 2943 1420 2949 1426
rect 2997 1420 3003 1426
rect 2937 1414 2943 1420
rect 3003 1414 3009 1420
rect 2937 1360 2943 1366
rect 3003 1360 3009 1366
rect 2943 1354 2949 1360
rect 2997 1354 3003 1360
rect 4599 1332 4605 1338
rect 4653 1332 4659 1338
rect 4593 1326 4599 1332
rect 4659 1326 4665 1332
rect 4593 1272 4599 1278
rect 4659 1272 4665 1278
rect 4599 1266 4605 1272
rect 4653 1266 4659 1272
rect 2667 1244 2673 1250
rect 2721 1244 2727 1250
rect 2661 1238 2667 1244
rect 2727 1238 2733 1244
rect 2661 1184 2667 1190
rect 2727 1184 2733 1190
rect 2667 1178 2673 1184
rect 2721 1178 2727 1184
rect 2391 1156 2397 1162
rect 2445 1156 2451 1162
rect 2385 1150 2391 1156
rect 2451 1150 2457 1156
rect 2385 1096 2391 1102
rect 2451 1096 2457 1102
rect 2391 1090 2397 1096
rect 2445 1090 2451 1096
rect 183 1068 189 1074
rect 237 1068 243 1074
rect 177 1062 183 1068
rect 243 1062 249 1068
rect 177 1008 183 1014
rect 243 1008 249 1014
rect 183 1002 189 1008
rect 237 1002 243 1008
rect 2115 980 2121 986
rect 2169 980 2175 986
rect 2109 974 2115 980
rect 2175 974 2181 980
rect 2109 920 2115 926
rect 2175 920 2181 926
rect 2115 914 2121 920
rect 2169 914 2175 920
rect 459 892 465 898
rect 513 892 519 898
rect 453 886 459 892
rect 519 886 525 892
rect 453 832 459 838
rect 519 832 525 838
rect 459 826 465 832
rect 513 826 519 832
rect 1839 804 1845 810
rect 1893 804 1899 810
rect 1833 798 1839 804
rect 1899 798 1905 804
rect 1833 744 1839 750
rect 1899 744 1905 750
rect 1839 738 1845 744
rect 1893 738 1899 744
rect 735 716 741 722
rect 789 716 795 722
rect 729 710 735 716
rect 795 710 801 716
rect 729 656 735 662
rect 795 656 801 662
rect 735 650 741 656
rect 789 650 795 656
rect 1563 628 1569 634
rect 1617 628 1623 634
rect 1557 622 1563 628
rect 1623 622 1629 628
rect 1557 568 1563 574
rect 1623 568 1629 574
rect 1563 562 1569 568
rect 1617 562 1623 568
rect 1011 540 1017 546
rect 1065 540 1071 546
rect 1005 534 1011 540
rect 1071 534 1077 540
rect 1005 480 1011 486
rect 1071 480 1077 486
rect 1011 474 1017 480
rect 1065 474 1071 480
rect 1287 452 1293 458
rect 1341 452 1347 458
rect 1281 446 1287 452
rect 1347 446 1353 452
rect 1281 392 1287 398
rect 1347 392 1353 398
rect 1287 386 1293 392
rect 1341 386 1347 392
<< pwell >>
rect -169 -173 4803 365
<< mvpsubdiff >>
rect -133 317 4767 329
rect -133 283 -25 317
rect 4659 283 4767 317
rect -133 271 4767 283
rect -133 221 -75 271
rect -133 -29 -121 221
rect -87 -29 -75 221
rect -133 -79 -75 -29
rect 4709 221 4767 271
rect 4709 -29 4721 221
rect 4755 -29 4767 221
rect 4709 -79 4767 -29
rect -133 -91 4767 -79
rect -133 -125 -25 -91
rect 4659 -125 4767 -91
rect -133 -137 4767 -125
<< mvpsubdiffcont >>
rect -25 283 4659 317
rect -121 -29 -87 221
rect 4721 -29 4755 221
rect -25 -125 4659 -91
<< locali >>
rect -121 283 -25 317
rect 4659 283 4755 317
rect -121 221 -87 283
rect -121 -91 -87 -29
rect 4721 221 4755 283
rect 4721 -91 4755 -29
rect -121 -125 -25 -91
rect 4659 -125 4755 -91
<< metal1 >>
rect 3771 1860 3831 1866
rect 3495 1772 3555 1778
rect 3219 1596 3279 1602
rect 2943 1420 3003 1426
rect 2667 1244 2727 1250
rect 2391 1156 2451 1162
rect 183 1068 243 1074
rect 183 23 243 1008
rect 2115 980 2175 986
rect 459 892 519 898
rect 459 23 519 832
rect 1839 804 1899 810
rect 735 716 795 722
rect 735 23 795 656
rect 1563 628 1623 634
rect 1011 540 1071 546
rect 1011 23 1071 480
rect 1287 452 1347 458
rect 1287 23 1347 392
rect 1563 23 1623 568
rect 1839 23 1899 744
rect 2115 23 2175 920
rect 2391 23 2451 1096
rect 2667 23 2727 1184
rect 2943 23 3003 1360
rect 3219 23 3279 1536
rect 3495 23 3555 1712
rect 3771 23 3831 1800
rect 4047 1684 4107 1690
rect 4047 23 4107 1624
rect 4323 1508 4383 1514
rect 4323 23 4383 1448
rect 4599 1332 4659 1338
rect 4599 23 4659 1272
<< via1 >>
rect 3771 1800 3831 1860
rect 3495 1712 3555 1772
rect 3219 1536 3279 1596
rect 2943 1360 3003 1420
rect 2667 1184 2727 1244
rect 2391 1096 2451 1156
rect 183 1008 243 1068
rect 2115 920 2175 980
rect 459 832 519 892
rect 1839 744 1899 804
rect 735 656 795 716
rect 1563 568 1623 628
rect 1011 480 1071 540
rect 1287 392 1347 452
rect 4047 1624 4107 1684
rect 4323 1448 4383 1508
rect 4599 1272 4659 1332
use hnmos_1  hnmos_1_1
timestamp 1749548291
transform 1 0 4428 0 1 -6
box -41 3 235 201
use hnmos_4  hnmos_4_0
timestamp 1749548291
transform 1 0 -21 0 1 -3
box -8 0 1096 198
use hnmos_4  hnmos_4_1
timestamp 1749548291
transform 1 0 1083 0 1 -3
box -8 0 1096 198
use hnmos_4  hnmos_4_2
timestamp 1749548291
transform 1 0 2187 0 1 -3
box -8 0 1096 198
use hnmos_4  hnmos_4_3
timestamp 1749548291
transform 1 0 3291 0 1 -3
box -8 0 1096 198
<< end >>
