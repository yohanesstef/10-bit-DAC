magic
tech sky130A
magscale 1 2
timestamp 1749147130
<< pwell >>
rect -307 -796 307 796
<< psubdiff >>
rect -271 726 -175 760
rect 175 726 271 760
rect -271 664 -237 726
rect 237 664 271 726
rect -271 -726 -237 -664
rect 237 -726 271 -664
rect -271 -760 -175 -726
rect 175 -760 271 -726
<< psubdiffcont >>
rect -175 726 175 760
rect -271 -664 -237 664
rect 237 -664 271 664
rect -175 -760 175 -726
<< xpolycontact >>
rect -141 198 141 630
rect -141 -630 141 -198
<< xpolyres >>
rect -141 -198 141 198
<< locali >>
rect -271 726 -175 760
rect 175 726 271 760
rect -271 664 -237 726
rect 237 664 271 726
rect -271 -726 -237 -664
rect 237 -726 271 -664
rect -271 -760 -175 -726
rect 175 -760 271 -726
<< viali >>
rect -125 215 125 612
rect -125 -612 125 -215
<< metal1 >>
rect -131 612 131 624
rect -131 215 -125 612
rect 125 215 131 612
rect -131 203 131 215
rect -131 -215 131 -203
rect -131 -612 -125 -215
rect 125 -612 131 -215
rect -131 -624 131 -612
<< properties >>
string FIXED_BBOX -254 -743 254 743
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 2.143 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 3.306k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
