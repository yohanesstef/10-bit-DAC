magic
tech sky130A
magscale 1 2
timestamp 1749488215
<< magnet >>
rect 1829 4813 1857 4841
rect 2653 4813 2681 4841
rect 2709 4813 2737 4841
rect 3533 4813 3561 4841
rect 1801 4785 1889 4813
rect 1829 4753 1889 4785
rect 1917 4753 1977 4813
rect 2005 4753 2065 4813
rect 2093 4753 2153 4813
rect 2181 4753 2241 4813
rect 2269 4753 2329 4813
rect 2357 4753 2417 4813
rect 2445 4753 2505 4813
rect 2533 4753 2593 4813
rect 2621 4785 2769 4813
rect 2621 4753 2681 4785
rect 2709 4753 2769 4785
rect 2797 4753 2857 4813
rect 2885 4753 2945 4813
rect 2973 4753 3033 4813
rect 3061 4753 3121 4813
rect 3149 4753 3209 4813
rect 3237 4753 3297 4813
rect 3325 4753 3385 4813
rect 3413 4753 3473 4813
rect 3501 4785 3589 4813
rect 3501 4753 3561 4785
rect 1829 4665 1889 4725
rect 2269 4665 2329 4725
rect 2621 4665 2681 4725
rect 2709 4665 2769 4725
rect 3149 4665 3209 4725
rect 3501 4665 3561 4725
rect 1829 4577 1889 4637
rect 2269 4577 2329 4637
rect 2621 4577 2681 4637
rect 2709 4577 2769 4637
rect 3149 4577 3209 4637
rect 3501 4577 3561 4637
rect 1829 4489 1889 4549
rect 2269 4489 2329 4549
rect 2621 4489 2681 4549
rect 2709 4489 2769 4549
rect 3149 4489 3209 4549
rect 3501 4489 3561 4549
rect 1829 4401 1889 4461
rect 2269 4401 2329 4461
rect 2621 4401 2681 4461
rect 2709 4401 2769 4461
rect 3149 4401 3209 4461
rect 3501 4401 3561 4461
rect 1829 4313 1889 4373
rect 2269 4313 2329 4373
rect 2621 4313 2681 4373
rect 2709 4313 2769 4373
rect 3149 4313 3209 4373
rect 3501 4313 3561 4373
rect 1829 4225 1889 4285
rect 2269 4225 2329 4285
rect 2621 4225 2681 4285
rect 2709 4225 2769 4285
rect 3149 4225 3209 4285
rect 3501 4225 3561 4285
rect 1829 4137 1889 4197
rect 2269 4137 2329 4197
rect 2621 4137 2681 4197
rect 2709 4137 2769 4197
rect 3149 4137 3209 4197
rect 3501 4137 3561 4197
rect 1829 4049 1889 4109
rect 2269 4049 2329 4109
rect 2621 4049 2681 4109
rect 2709 4049 2769 4109
rect 3149 4049 3209 4109
rect 3501 4049 3561 4109
rect 1829 3989 1889 4021
rect 1801 3961 1889 3989
rect 1917 3961 1977 4021
rect 2005 3961 2065 4021
rect 2093 3961 2153 4021
rect 2181 3961 2241 4021
rect 2269 3961 2329 4021
rect 2357 3961 2417 4021
rect 2445 3961 2505 4021
rect 2533 3961 2593 4021
rect 2621 3989 2681 4021
rect 2709 3989 2769 4021
rect 2621 3961 2769 3989
rect 2797 3961 2857 4021
rect 2885 3961 2945 4021
rect 2973 3961 3033 4021
rect 3061 3961 3121 4021
rect 3149 3961 3209 4021
rect 3237 3961 3297 4021
rect 3325 3961 3385 4021
rect 3413 3961 3473 4021
rect 3501 3989 3561 4021
rect 3501 3961 3589 3989
rect 1829 3933 1857 3961
rect 2653 3933 2681 3961
rect 2709 3933 2737 3961
rect 3533 3933 3561 3961
rect 1801 3905 1889 3933
rect 1829 3873 1889 3905
rect 1917 3873 1977 3933
rect 2005 3873 2065 3933
rect 2093 3873 2153 3933
rect 2181 3873 2241 3933
rect 2269 3873 2329 3933
rect 2357 3873 2417 3933
rect 2445 3873 2505 3933
rect 2533 3873 2593 3933
rect 2621 3905 2769 3933
rect 2621 3873 2681 3905
rect 2709 3873 2769 3905
rect 2797 3873 2857 3933
rect 2885 3873 2945 3933
rect 2973 3873 3033 3933
rect 3061 3873 3121 3933
rect 3149 3873 3209 3933
rect 3237 3873 3297 3933
rect 3325 3873 3385 3933
rect 3413 3873 3473 3933
rect 3501 3905 3589 3933
rect 3501 3873 3561 3905
rect 1829 3785 1889 3845
rect 2269 3785 2329 3845
rect 2621 3785 2681 3845
rect 2709 3785 2769 3845
rect 3149 3785 3209 3845
rect 3501 3785 3561 3845
rect 1829 3697 1889 3757
rect 2269 3697 2329 3757
rect 2621 3697 2681 3757
rect 2709 3697 2769 3757
rect 3149 3697 3209 3757
rect 3501 3697 3561 3757
rect 1829 3609 1889 3669
rect 2269 3609 2329 3669
rect 2621 3609 2681 3669
rect 2709 3609 2769 3669
rect 3149 3609 3209 3669
rect 3501 3609 3561 3669
rect 1829 3521 1889 3581
rect 2269 3521 2329 3581
rect 2621 3521 2681 3581
rect 2709 3521 2769 3581
rect 3149 3521 3209 3581
rect 3501 3521 3561 3581
rect 1829 3433 1889 3493
rect 2269 3433 2329 3493
rect 2621 3433 2681 3493
rect 2709 3433 2769 3493
rect 3149 3433 3209 3493
rect 3501 3433 3561 3493
rect 1829 3345 1889 3405
rect 2269 3345 2329 3405
rect 2621 3345 2681 3405
rect 2709 3345 2769 3405
rect 3149 3345 3209 3405
rect 3501 3345 3561 3405
rect 1829 3257 1889 3317
rect 2269 3257 2329 3317
rect 2621 3257 2681 3317
rect 2709 3257 2769 3317
rect 3149 3257 3209 3317
rect 3501 3257 3561 3317
rect 1829 3169 1889 3229
rect 2269 3169 2329 3229
rect 2621 3169 2681 3229
rect 2709 3169 2769 3229
rect 3149 3169 3209 3229
rect 3501 3169 3561 3229
rect 1829 3109 1889 3141
rect 1801 3081 1889 3109
rect 1917 3081 1977 3141
rect 2005 3081 2065 3141
rect 2093 3081 2153 3141
rect 2181 3081 2241 3141
rect 2269 3081 2329 3141
rect 2357 3081 2417 3141
rect 2445 3081 2505 3141
rect 2533 3081 2593 3141
rect 2621 3109 2681 3141
rect 2709 3109 2769 3141
rect 2621 3081 2769 3109
rect 2797 3081 2857 3141
rect 2885 3081 2945 3141
rect 2973 3081 3033 3141
rect 3061 3081 3121 3141
rect 3149 3081 3209 3141
rect 3237 3081 3297 3141
rect 3325 3081 3385 3141
rect 3413 3081 3473 3141
rect 3501 3109 3561 3141
rect 3501 3081 3589 3109
rect 1829 3053 1857 3081
rect 2653 3053 2681 3081
rect 2709 3053 2737 3081
rect 3533 3053 3561 3081
<< end >>
