magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -781 307 781
<< psubdiff >>
rect -271 711 -175 745
rect 175 711 271 745
rect -271 649 -237 711
rect 237 649 271 711
rect -271 -711 -237 -649
rect 237 -711 271 -649
rect -271 -745 -175 -711
rect 175 -745 271 -711
<< psubdiffcont >>
rect -175 711 175 745
rect -271 -649 -237 649
rect 237 -649 271 649
rect -175 -745 175 -711
<< xpolycontact >>
rect -141 183 141 615
rect -141 -615 141 -183
<< xpolyres >>
rect -141 -183 141 183
<< locali >>
rect -271 711 -175 745
rect 175 711 271 745
rect -271 649 -237 711
rect 237 649 271 711
rect -271 -711 -237 -649
rect 237 -711 271 -649
rect -271 -745 -175 -711
rect 175 -745 271 -711
<< viali >>
rect -125 200 125 597
rect -125 -597 125 -200
<< metal1 >>
rect -131 597 131 609
rect -131 200 -125 597
rect 125 200 131 597
rect -131 188 131 200
rect -131 -200 131 -188
rect -131 -597 -125 -200
rect 125 -597 131 -200
rect -131 -609 131 -597
<< properties >>
string FIXED_BBOX -254 -728 254 728
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.989 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 3.088k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
