magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1129 307 1129
<< psubdiff >>
rect -271 1059 -175 1093
rect 175 1059 271 1093
rect -271 997 -237 1059
rect 237 997 271 1059
rect -271 -1059 -237 -997
rect 237 -1059 271 -997
rect -271 -1093 -175 -1059
rect 175 -1093 271 -1059
<< psubdiffcont >>
rect -175 1059 175 1093
rect -271 -997 -237 997
rect 237 -997 271 997
rect -175 -1093 175 -1059
<< xpolycontact >>
rect -141 531 141 963
rect -141 -963 141 -531
<< xpolyres >>
rect -141 -531 141 531
<< locali >>
rect -271 1059 -175 1093
rect 175 1059 271 1093
rect -271 997 -237 1059
rect 237 997 271 1059
rect -271 -1059 -237 -997
rect 237 -1059 271 -997
rect -271 -1093 -175 -1059
rect 175 -1093 271 -1059
<< viali >>
rect -125 548 125 945
rect -125 -945 125 -548
<< metal1 >>
rect -131 945 131 957
rect -131 548 -125 945
rect 125 548 131 945
rect -131 536 131 548
rect -131 -548 131 -536
rect -131 -945 -125 -548
rect 125 -945 131 -548
rect -131 -957 131 -945
<< properties >>
string FIXED_BBOX -254 -1076 254 1076
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 5.474 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 8.031k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
