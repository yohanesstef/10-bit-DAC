magic
tech sky130A
magscale 1 2
timestamp 1749147130
<< pwell >>
rect -307 -760 307 760
<< psubdiff >>
rect -271 690 -175 724
rect 175 690 271 724
rect -271 628 -237 690
rect 237 628 271 690
rect -271 -690 -237 -628
rect 237 -690 271 -628
rect -271 -724 -175 -690
rect 175 -724 271 -690
<< psubdiffcont >>
rect -175 690 175 724
rect -271 -628 -237 628
rect 237 -628 271 628
rect -175 -724 175 -690
<< xpolycontact >>
rect -141 162 141 594
rect -141 -594 141 -162
<< xpolyres >>
rect -141 -162 141 162
<< locali >>
rect -271 690 -175 724
rect 175 690 271 724
rect -271 628 -237 690
rect 237 628 271 690
rect -271 -690 -237 -628
rect 237 -690 271 -628
rect -271 -724 -175 -690
rect 175 -724 271 -690
<< viali >>
rect -125 179 125 576
rect -125 -576 125 -179
<< metal1 >>
rect -131 576 131 588
rect -131 179 -125 576
rect 125 179 131 576
rect -131 167 131 179
rect -131 -179 131 -167
rect -131 -576 -125 -179
rect 125 -576 131 -179
rect -131 -588 131 -576
<< properties >>
string FIXED_BBOX -254 -707 254 707
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.784 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 2.797k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
