magic
tech sky130A
magscale 1 2
timestamp 1750052349
<< mvnsubdiffcont >>
rect 12732 1529 12766 3161
rect 21906 1529 21940 3161
rect 12732 1495 21940 1529
rect 12732 -137 12766 1495
rect 21906 -137 21940 1495
<< metal2 >>
rect 17362 2694 17536 2696
rect 17362 2638 17371 2694
rect 17427 2638 17536 2694
rect 17362 2636 17536 2638
rect 17142 2606 17310 2608
rect 17142 2550 17245 2606
rect 17301 2550 17310 2606
rect 17142 2548 17310 2550
rect 17488 2342 18105 2344
rect 17488 2286 17497 2342
rect 17553 2286 18105 2342
rect 17488 2284 18105 2286
rect 16937 738 17562 740
rect 16937 682 17497 738
rect 17553 682 17562 738
rect 16937 680 17562 682
rect 17236 474 17533 476
rect 17236 418 17245 474
rect 17301 418 17533 474
rect 17236 416 17533 418
rect 17121 386 17436 388
rect 17121 330 17371 386
rect 17427 330 17436 386
rect 17121 328 17436 330
<< via2 >>
rect 17119 3078 17175 3134
rect 16993 2990 17049 3046
rect 16741 2814 16797 2870
rect 17371 2638 17427 2694
rect 17245 2550 17301 2606
rect 17497 2286 17553 2342
rect 16867 2198 16923 2254
rect 17749 1670 17805 1726
rect 17623 1582 17679 1638
rect 17623 1386 17679 1442
rect 17749 1298 17805 1354
rect 16867 770 16923 826
rect 17497 682 17553 738
rect 17245 418 17301 474
rect 17371 330 17427 386
rect 16741 154 16797 210
rect 16993 -22 17049 34
rect 17119 -110 17175 -54
<< metal3 >>
rect 16736 2870 16802 3174
rect 16736 2814 16741 2870
rect 16797 2814 16802 2870
rect 16736 210 16802 2814
rect 16862 2254 16928 3174
rect 16862 2198 16867 2254
rect 16923 2198 16928 2254
rect 16862 826 16928 2198
rect 16862 770 16867 826
rect 16923 770 16928 826
rect 16862 765 16928 770
rect 16988 3046 17054 3174
rect 16988 2990 16993 3046
rect 17049 2990 17054 3046
rect 16736 154 16741 210
rect 16797 154 16802 210
rect 16736 149 16802 154
rect 16988 34 17054 2990
rect 16988 -22 16993 34
rect 17049 -22 17054 34
rect 16988 -29 17054 -22
rect 17114 3134 17180 3174
rect 17114 3078 17119 3134
rect 17175 3078 17180 3134
rect 17114 -54 17180 3078
rect 17240 2606 17306 3174
rect 17240 2550 17245 2606
rect 17301 2550 17306 2606
rect 17240 474 17306 2550
rect 17240 418 17245 474
rect 17301 418 17306 474
rect 17240 413 17306 418
rect 17366 2694 17432 3174
rect 17366 2638 17371 2694
rect 17427 2638 17432 2694
rect 17366 386 17432 2638
rect 17492 2342 17558 3174
rect 17492 2286 17497 2342
rect 17553 2286 17558 2342
rect 17492 738 17558 2286
rect 17618 1638 17684 3174
rect 17618 1582 17623 1638
rect 17679 1582 17684 1638
rect 17618 1442 17684 1582
rect 17618 1386 17623 1442
rect 17679 1386 17684 1442
rect 17618 1381 17684 1386
rect 17744 1726 17810 3174
rect 17744 1670 17749 1726
rect 17805 1670 17810 1726
rect 17744 1354 17810 1670
rect 17744 1298 17749 1354
rect 17805 1298 17810 1354
rect 17744 1293 17810 1298
rect 17492 682 17497 738
rect 17553 682 17558 738
rect 17492 677 17558 682
rect 17366 330 17371 386
rect 17427 330 17432 386
rect 17366 325 17432 330
rect 17114 -110 17119 -54
rect 17175 -110 17180 -54
rect 17114 -122 17180 -110
use cm_pcell2_half  cm_pcell2_half_0
timestamp 1749897485
transform 1 0 12450 0 1 3120
box 204 -1704 9568 180
use cm_pcell2_half  cm_pcell2_half_1
timestamp 1749897485
transform -1 0 22222 0 -1 -96
box 204 -1704 9568 180
<< end >>
