magic
tech sky130A
magscale 1 2
timestamp 1750167460
use top_buffer_opamp  top_buffer_opamp_0
timestamp 1750156376
transform -1 0 -2156 0 1 9674
box -12462 -8798 520 13398
use top_digital_cell  top_digital_cell_0
timestamp 1750151992
transform 0 -1 43880 1 0 1486
box -31 -831 19579 4114
use top_segment_1  top_segment_1_0
timestamp 1749633251
transform 1 0 25398 0 1 1220
box -385 -49 14453 8429
use top_segment_2  top_segment_2_0
timestamp 1749580325
transform -1 0 32595 0 -1 22873
box -870 14 15704 7051
use top_segment_3  top_segment_3_0
timestamp 1749552768
transform -1 0 22205 0 -1 23118
box 5007 266 11251 6636
use top_segment_4  top_segment_4_1
timestamp 1749664768
transform 1 0 -18626 0 1 13460
box 29493 -12226 43322 -3773
<< end >>
