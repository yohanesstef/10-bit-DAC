magic
tech sky130A
magscale 1 2
timestamp 1750150226
<< metal3 >>
rect 2268 9190 6412 9206
rect 2268 9126 2285 9190
rect 2349 9126 3297 9190
rect 3361 9126 4309 9190
rect 4373 9126 5322 9190
rect 5386 9126 6333 9190
rect 6397 9126 6412 9190
rect 2268 9110 6412 9126
rect -3804 8470 340 8486
rect -3804 8406 -3787 8470
rect -3723 8406 -2775 8470
rect -2711 8406 -1763 8470
rect -1699 8406 -751 8470
rect -687 8406 261 8470
rect 325 8406 340 8470
rect -3804 8390 340 8406
rect 820 7670 3664 7766
<< via3 >>
rect 2285 9126 2349 9190
rect 3297 9126 3361 9190
rect 4309 9126 4373 9190
rect 5322 9126 5386 9190
rect 6333 9126 6397 9190
rect -3787 8406 -3723 8470
rect -2775 8406 -2711 8470
rect -1763 8406 -1699 8470
rect -751 8406 -687 8470
rect 261 8406 325 8470
use opa_cap_cell  opa_cap_cell_0
timestamp 1750148716
transform 1 0 -571 0 1 10026
box 1635 -3628 8479 452
use opa_cap_cell  opa_cap_cell_1
timestamp 1750148716
transform 1 0 -6643 0 1 10026
box 1635 -3628 8479 452
<< end >>
