magic
tech sky130A
magscale 1 2
timestamp 1749736748
<< magnet >>
rect 2595 -4415 2647 -4363
<< pwell >>
rect 579 -4820 2781 -4413
rect 579 -5683 2781 -5501
<< locali >>
rect 2370 -4394 2378 -4367
rect 2616 -4367 2650 -4360
rect 2344 -4401 2378 -4394
rect 2639 -4394 2650 -4367
rect 690 -4847 724 -4832
rect 690 -4866 706 -4847
rect 1097 -4865 1289 -4831
rect 695 -5459 729 -5439
rect 695 -5473 720 -5459
rect 1185 -5473 1187 -5439
rect 1221 -5473 1240 -5439
rect 1185 -5489 1240 -5473
<< viali >>
rect 1060 -4293 1094 -4259
rect 1341 -4317 1375 -4283
rect 698 -4394 732 -4360
rect 866 -4393 900 -4359
rect 978 -4394 1012 -4360
rect 1132 -4394 1166 -4360
rect 1244 -4394 1278 -4360
rect 1412 -4394 1446 -4360
rect 1580 -4394 1614 -4360
rect 1902 -4394 1936 -4360
rect 2071 -4394 2105 -4360
rect 2183 -4394 2217 -4360
rect 2336 -4394 2370 -4360
rect 2448 -4394 2482 -4360
rect 2605 -4401 2639 -4367
rect 1984 -4450 2018 -4416
rect 867 -4506 901 -4472
rect 2336 -4506 2370 -4472
rect 2532 -4503 2566 -4469
rect 904 -4732 938 -4698
rect 1343 -4732 1377 -4698
rect 1435 -4732 1469 -4698
rect 1810 -4794 1844 -4760
rect 706 -4881 740 -4847
rect 809 -4881 843 -4847
rect 1063 -4865 1097 -4831
rect 1615 -4849 1649 -4815
rect 1716 -4865 1750 -4831
rect 1901 -4877 1935 -4843
rect 2033 -4866 2067 -4832
rect 2496 -4865 2530 -4831
rect 1516 -4951 1550 -4917
rect 973 -5007 1007 -4973
rect 720 -5493 754 -5459
rect 866 -5473 900 -5439
rect 978 -5473 1012 -5439
rect 1187 -5473 1221 -5439
rect 1340 -5473 1374 -5439
rect 1427 -5474 1461 -5440
rect 1617 -5473 1651 -5439
rect 1790 -5473 1824 -5439
rect 1902 -5473 1936 -5439
rect 1988 -5483 2022 -5449
rect 2101 -5493 2135 -5459
rect 2202 -5494 2236 -5460
rect 2354 -5494 2388 -5460
rect 2504 -5485 2538 -5451
rect 1156 -5559 1190 -5525
rect 878 -5606 912 -5572
rect 1902 -5573 1936 -5539
rect 2342 -5594 2376 -5560
<< metal1 >>
rect -147 -4030 714 -4024
rect 9 -4114 714 -4030
rect -147 -4120 714 -4114
rect 2692 -4030 3311 -4024
rect 2692 -4114 3155 -4030
rect 2692 -4120 3311 -4114
rect 221 -4159 1163 -4153
rect 221 -4211 227 -4159
rect 279 -4181 1163 -4159
rect 279 -4211 285 -4181
rect 221 -4217 285 -4211
rect 313 -4215 1009 -4209
rect 313 -4267 319 -4215
rect 371 -4237 1009 -4215
rect 371 -4267 377 -4237
rect 313 -4273 377 -4267
rect 405 -4271 897 -4265
rect 405 -4323 411 -4271
rect 463 -4293 897 -4271
rect 463 -4323 469 -4293
rect 405 -4329 469 -4323
rect 869 -4353 897 -4293
rect 686 -4360 744 -4354
rect 686 -4363 698 -4360
rect 497 -4369 698 -4363
rect 497 -4421 503 -4369
rect 555 -4391 698 -4369
rect 555 -4421 561 -4391
rect 686 -4394 698 -4391
rect 732 -4394 744 -4360
rect 686 -4400 744 -4394
rect 854 -4359 912 -4353
rect 981 -4354 1009 -4237
rect 1051 -4250 1103 -4244
rect 1051 -4308 1103 -4302
rect 1135 -4354 1163 -4181
rect 2073 -4159 2943 -4153
rect 2073 -4181 2885 -4159
rect 1341 -4277 1611 -4265
rect 1329 -4283 1611 -4277
rect 1329 -4317 1341 -4283
rect 1375 -4293 1611 -4283
rect 1375 -4317 1387 -4293
rect 1329 -4323 1387 -4317
rect 1224 -4351 1284 -4345
rect 854 -4393 866 -4359
rect 900 -4393 912 -4359
rect 854 -4399 912 -4393
rect 966 -4360 1024 -4354
rect 966 -4394 978 -4360
rect 1012 -4394 1024 -4360
rect 966 -4400 1024 -4394
rect 1120 -4360 1178 -4354
rect 1120 -4394 1132 -4360
rect 1166 -4394 1178 -4360
rect 1120 -4400 1178 -4394
rect 1276 -4360 1284 -4351
rect 1583 -4354 1611 -4293
rect 1886 -4347 1892 -4295
rect 1944 -4347 1950 -4295
rect 1886 -4353 1950 -4347
rect 2073 -4348 2101 -4181
rect 2185 -4237 2759 -4209
rect 2879 -4211 2885 -4181
rect 2937 -4211 2943 -4159
rect 2879 -4217 2943 -4211
rect 2185 -4348 2213 -4237
rect 2339 -4293 2703 -4265
rect 2339 -4348 2367 -4293
rect 1278 -4394 1284 -4360
rect 1276 -4403 1284 -4394
rect 1400 -4360 1458 -4354
rect 1400 -4394 1412 -4360
rect 1446 -4394 1458 -4360
rect 1400 -4400 1458 -4394
rect 1568 -4360 1626 -4354
rect 1568 -4394 1580 -4360
rect 1614 -4394 1626 -4360
rect 1568 -4400 1626 -4394
rect 1896 -4360 1942 -4353
rect 1896 -4394 1902 -4360
rect 1936 -4394 1942 -4360
rect 1224 -4409 1284 -4403
rect 497 -4427 561 -4421
rect 855 -4472 913 -4466
rect 855 -4506 867 -4472
rect 901 -4475 913 -4472
rect 1415 -4475 1443 -4400
rect 1896 -4406 1942 -4394
rect 2065 -4360 2111 -4348
rect 2065 -4394 2071 -4360
rect 2105 -4394 2111 -4360
rect 1975 -4407 2027 -4401
rect 2065 -4406 2111 -4394
rect 2177 -4360 2223 -4348
rect 2177 -4394 2183 -4360
rect 2217 -4394 2223 -4360
rect 2177 -4406 2223 -4394
rect 2330 -4360 2376 -4348
rect 2330 -4394 2336 -4360
rect 2370 -4394 2376 -4360
rect 2330 -4406 2376 -4394
rect 2442 -4360 2488 -4348
rect 2442 -4394 2448 -4360
rect 2482 -4394 2488 -4360
rect 2442 -4406 2488 -4394
rect 2593 -4363 2647 -4355
rect 1972 -4456 1975 -4410
rect 2027 -4456 2030 -4410
rect 1975 -4465 2027 -4459
rect 901 -4503 1443 -4475
rect 2324 -4472 2382 -4466
rect 901 -4506 913 -4503
rect 855 -4512 913 -4506
rect 2324 -4506 2336 -4472
rect 2370 -4475 2382 -4472
rect 2451 -4475 2479 -4406
rect 2593 -4415 2595 -4363
rect 2593 -4421 2647 -4415
rect 2675 -4401 2703 -4293
rect 2731 -4345 2759 -4237
rect 2971 -4315 3035 -4309
rect 2971 -4345 2977 -4315
rect 2731 -4367 2977 -4345
rect 3029 -4367 3035 -4315
rect 2731 -4373 3035 -4367
rect 3063 -4371 3127 -4365
rect 3063 -4401 3069 -4371
rect 2675 -4423 3069 -4401
rect 3121 -4423 3127 -4371
rect 2675 -4429 3127 -4423
rect 2370 -4503 2479 -4475
rect 2523 -4460 2575 -4454
rect 2370 -4506 2382 -4503
rect 2324 -4512 2382 -4506
rect 2523 -4518 2575 -4512
rect 37 -4574 714 -4568
rect 193 -4658 714 -4574
rect 37 -4664 714 -4658
rect 2691 -4574 3495 -4568
rect 2691 -4658 3339 -4574
rect 2691 -4664 3495 -4658
rect 892 -4698 950 -4692
rect 892 -4701 904 -4698
rect 405 -4707 904 -4701
rect 405 -4759 411 -4707
rect 463 -4729 904 -4707
rect 463 -4759 469 -4729
rect 892 -4732 904 -4729
rect 938 -4701 950 -4698
rect 1331 -4698 1389 -4692
rect 1331 -4701 1343 -4698
rect 938 -4729 1343 -4701
rect 938 -4732 950 -4729
rect 892 -4738 950 -4732
rect 1331 -4732 1343 -4729
rect 1377 -4732 1389 -4698
rect 1331 -4738 1389 -4732
rect 1423 -4698 1481 -4692
rect 1423 -4732 1435 -4698
rect 1469 -4732 1481 -4698
rect 1423 -4738 1481 -4732
rect 1633 -4720 2907 -4692
rect 405 -4765 469 -4759
rect 1423 -4766 1451 -4738
rect 221 -4792 285 -4786
rect 221 -4844 227 -4792
rect 279 -4822 285 -4792
rect 614 -4794 1451 -4766
rect 614 -4822 642 -4794
rect 1633 -4809 1661 -4720
rect 2879 -4744 2907 -4720
rect 1800 -4760 2045 -4748
rect 1800 -4794 1810 -4760
rect 1844 -4776 2045 -4760
rect 1844 -4794 1858 -4776
rect 1800 -4806 1858 -4794
rect 1603 -4815 1661 -4809
rect 279 -4844 642 -4822
rect 221 -4850 642 -4844
rect 694 -4847 752 -4836
rect 694 -4878 706 -4847
rect 313 -4881 706 -4878
rect 740 -4881 752 -4847
rect 313 -4884 752 -4881
rect 313 -4936 319 -4884
rect 371 -4886 752 -4884
rect 797 -4847 855 -4841
rect 797 -4881 809 -4847
rect 843 -4881 855 -4847
rect 1044 -4874 1051 -4822
rect 1103 -4874 1109 -4822
rect 1603 -4849 1615 -4815
rect 1649 -4849 1661 -4815
rect 1603 -4855 1661 -4849
rect 1704 -4831 1765 -4825
rect 1704 -4865 1716 -4831
rect 1750 -4865 1765 -4831
rect 2017 -4826 2045 -4776
rect 2879 -4750 2943 -4744
rect 2879 -4802 2885 -4750
rect 2937 -4802 2943 -4750
rect 2879 -4808 2943 -4802
rect 2017 -4832 2079 -4826
rect 1704 -4871 1765 -4865
rect 371 -4906 747 -4886
rect 797 -4887 855 -4881
rect 371 -4936 377 -4906
rect 313 -4942 377 -4936
rect 813 -5056 841 -4887
rect 1504 -4917 1562 -4911
rect 1504 -4951 1516 -4917
rect 1550 -4933 1562 -4917
rect 1737 -4933 1765 -4871
rect 1889 -4843 1947 -4837
rect 1889 -4877 1901 -4843
rect 1935 -4877 1947 -4843
rect 2017 -4866 2033 -4832
rect 2067 -4866 2079 -4832
rect 2017 -4872 2079 -4866
rect 2481 -4871 2487 -4819
rect 2539 -4871 2545 -4819
rect 1889 -4883 1947 -4877
rect 1550 -4951 1765 -4933
rect 1504 -4961 1765 -4951
rect 961 -4973 1019 -4967
rect 961 -5007 973 -4973
rect 1007 -4989 1019 -4973
rect 1905 -4989 1933 -4883
rect 1007 -5007 1933 -4989
rect 961 -5017 1933 -5007
rect 2787 -5026 2851 -5020
rect 2787 -5056 2793 -5026
rect 813 -5078 2793 -5056
rect 2845 -5078 2851 -5026
rect 813 -5084 2851 -5078
rect -147 -5118 714 -5112
rect 9 -5202 714 -5118
rect -147 -5208 714 -5202
rect 2692 -5118 3311 -5112
rect 2692 -5202 3155 -5118
rect 2692 -5208 3311 -5202
rect 221 -5266 285 -5260
rect 221 -5318 227 -5266
rect 279 -5283 285 -5266
rect 279 -5311 1443 -5283
rect 1603 -5292 1609 -5240
rect 1661 -5292 1667 -5240
rect 2879 -5253 2943 -5247
rect 2879 -5283 2885 -5253
rect 279 -5318 285 -5311
rect 221 -5324 285 -5318
rect 313 -5345 1009 -5339
rect 313 -5397 319 -5345
rect 371 -5367 1009 -5345
rect 371 -5397 377 -5367
rect 313 -5403 377 -5397
rect 405 -5422 469 -5416
rect 405 -5474 411 -5422
rect 463 -5451 469 -5422
rect 609 -5421 673 -5415
rect 609 -5451 615 -5421
rect 463 -5473 615 -5451
rect 667 -5473 673 -5421
rect 851 -5447 857 -5395
rect 909 -5447 915 -5395
rect 981 -5433 1009 -5367
rect 1175 -5395 1233 -5389
rect 1175 -5419 1178 -5395
rect 966 -5439 1024 -5433
rect 463 -5474 673 -5473
rect 405 -5479 673 -5474
rect 711 -5459 761 -5447
rect 405 -5480 469 -5479
rect 711 -5493 720 -5459
rect 754 -5493 761 -5459
rect 854 -5473 866 -5447
rect 900 -5473 912 -5447
rect 854 -5479 912 -5473
rect 966 -5473 978 -5439
rect 1012 -5473 1024 -5439
rect 1172 -5447 1178 -5419
rect 1230 -5419 1233 -5395
rect 1230 -5447 1236 -5419
rect 1172 -5448 1187 -5447
rect 966 -5479 1024 -5473
rect 1175 -5473 1187 -5448
rect 1221 -5448 1236 -5447
rect 1322 -5439 1386 -5432
rect 1221 -5473 1233 -5448
rect 1175 -5479 1233 -5473
rect 1322 -5451 1340 -5439
rect 1374 -5451 1386 -5439
rect 711 -5507 761 -5493
rect 1322 -5503 1328 -5451
rect 1380 -5503 1386 -5451
rect 1415 -5434 1443 -5311
rect 1639 -5433 1667 -5292
rect 1793 -5305 2885 -5283
rect 2937 -5305 2943 -5253
rect 1793 -5311 2943 -5305
rect 1793 -5433 1821 -5311
rect 1905 -5345 2851 -5339
rect 1905 -5367 2793 -5345
rect 1905 -5433 1933 -5367
rect 2787 -5397 2793 -5367
rect 2845 -5397 2851 -5345
rect 2787 -5403 2851 -5397
rect 2675 -5425 2739 -5419
rect 1415 -5440 1473 -5434
rect 1415 -5474 1427 -5440
rect 1461 -5474 1473 -5440
rect 1415 -5480 1473 -5474
rect 1605 -5439 1667 -5433
rect 1605 -5473 1617 -5439
rect 1651 -5473 1667 -5439
rect 1605 -5479 1667 -5473
rect 1778 -5439 1836 -5433
rect 1778 -5473 1790 -5439
rect 1824 -5473 1836 -5439
rect 1778 -5479 1836 -5473
rect 1890 -5439 1948 -5433
rect 1890 -5473 1902 -5439
rect 1936 -5473 1948 -5439
rect 1890 -5479 1948 -5473
rect 1976 -5449 2034 -5443
rect 1976 -5483 1988 -5449
rect 2022 -5483 2034 -5449
rect 2492 -5451 2550 -5445
rect 1976 -5489 2034 -5483
rect 1976 -5507 2004 -5489
rect 2086 -5503 2092 -5451
rect 2144 -5503 2150 -5451
rect 2186 -5503 2192 -5451
rect 2244 -5503 2250 -5451
rect 2338 -5503 2344 -5451
rect 2396 -5503 2402 -5451
rect 2492 -5463 2504 -5451
rect 2430 -5485 2504 -5463
rect 2538 -5485 2550 -5451
rect 2675 -5477 2681 -5425
rect 2733 -5455 2739 -5425
rect 2971 -5426 3035 -5420
rect 2971 -5455 2977 -5426
rect 2733 -5477 2977 -5455
rect 2675 -5478 2977 -5477
rect 3029 -5478 3035 -5426
rect 2675 -5483 3035 -5478
rect 2971 -5484 3035 -5483
rect 2430 -5491 2550 -5485
rect 498 -5508 761 -5507
rect 497 -5514 761 -5508
rect 497 -5566 503 -5514
rect 555 -5535 761 -5514
rect 555 -5566 561 -5535
rect 1142 -5559 1148 -5507
rect 1200 -5559 1206 -5507
rect 1905 -5533 2004 -5507
rect 497 -5572 561 -5566
rect 863 -5615 869 -5563
rect 921 -5615 928 -5563
rect 1142 -5565 1206 -5559
rect 1890 -5535 2004 -5533
rect 1890 -5539 1948 -5535
rect 1890 -5573 1902 -5539
rect 1936 -5573 1948 -5539
rect 1890 -5579 1948 -5573
rect 2330 -5560 2388 -5554
rect 2330 -5594 2342 -5560
rect 2376 -5563 2388 -5560
rect 2430 -5563 2458 -5491
rect 2376 -5591 2458 -5563
rect 2675 -5518 3127 -5512
rect 2675 -5570 2681 -5518
rect 2733 -5540 3069 -5518
rect 2733 -5570 2739 -5540
rect 2675 -5576 2739 -5570
rect 3063 -5570 3069 -5540
rect 3121 -5570 3127 -5518
rect 3063 -5576 3127 -5570
rect 2376 -5594 2388 -5591
rect 2330 -5600 2388 -5594
rect 37 -5662 714 -5656
rect 193 -5746 714 -5662
rect 37 -5752 714 -5746
rect 2663 -5662 3495 -5656
rect 2663 -5746 3339 -5662
rect 2663 -5752 3495 -5746
<< via1 >>
rect -147 -4114 9 -4030
rect 3155 -4114 3311 -4030
rect 227 -4211 279 -4159
rect 319 -4267 371 -4215
rect 411 -4323 463 -4271
rect 503 -4421 555 -4369
rect 1051 -4259 1103 -4250
rect 1051 -4293 1060 -4259
rect 1060 -4293 1094 -4259
rect 1094 -4293 1103 -4259
rect 1051 -4302 1103 -4293
rect 1224 -4360 1276 -4351
rect 1892 -4347 1944 -4295
rect 2885 -4211 2937 -4159
rect 1224 -4394 1244 -4360
rect 1244 -4394 1276 -4360
rect 1224 -4403 1276 -4394
rect 1975 -4416 2027 -4407
rect 1975 -4450 1984 -4416
rect 1984 -4450 2018 -4416
rect 2018 -4450 2027 -4416
rect 1975 -4459 2027 -4450
rect 2595 -4367 2647 -4363
rect 2595 -4401 2605 -4367
rect 2605 -4401 2639 -4367
rect 2639 -4401 2647 -4367
rect 2595 -4415 2647 -4401
rect 2977 -4367 3029 -4315
rect 3069 -4423 3121 -4371
rect 2523 -4469 2575 -4460
rect 2523 -4503 2532 -4469
rect 2532 -4503 2566 -4469
rect 2566 -4503 2575 -4469
rect 2523 -4512 2575 -4503
rect 37 -4658 193 -4574
rect 3339 -4658 3495 -4574
rect 411 -4759 463 -4707
rect 227 -4844 279 -4792
rect 319 -4936 371 -4884
rect 1051 -4831 1103 -4822
rect 1051 -4865 1063 -4831
rect 1063 -4865 1097 -4831
rect 1097 -4865 1103 -4831
rect 1051 -4874 1103 -4865
rect 2885 -4802 2937 -4750
rect 2487 -4831 2539 -4819
rect 2487 -4865 2496 -4831
rect 2496 -4865 2530 -4831
rect 2530 -4865 2539 -4831
rect 2487 -4871 2539 -4865
rect 2793 -5078 2845 -5026
rect -147 -5202 9 -5118
rect 3155 -5202 3311 -5118
rect 227 -5318 279 -5266
rect 1609 -5292 1661 -5240
rect 319 -5397 371 -5345
rect 411 -5474 463 -5422
rect 615 -5473 667 -5421
rect 857 -5439 909 -5395
rect 857 -5447 866 -5439
rect 866 -5447 900 -5439
rect 900 -5447 909 -5439
rect 1178 -5439 1230 -5395
rect 1178 -5447 1187 -5439
rect 1187 -5447 1221 -5439
rect 1221 -5447 1230 -5439
rect 1328 -5473 1340 -5451
rect 1340 -5473 1374 -5451
rect 1374 -5473 1380 -5451
rect 1328 -5503 1380 -5473
rect 2885 -5305 2937 -5253
rect 2793 -5397 2845 -5345
rect 2092 -5459 2144 -5451
rect 2092 -5493 2101 -5459
rect 2101 -5493 2135 -5459
rect 2135 -5493 2144 -5459
rect 2092 -5503 2144 -5493
rect 2192 -5460 2244 -5451
rect 2192 -5494 2202 -5460
rect 2202 -5494 2236 -5460
rect 2236 -5494 2244 -5460
rect 2192 -5503 2244 -5494
rect 2344 -5460 2396 -5451
rect 2344 -5494 2354 -5460
rect 2354 -5494 2388 -5460
rect 2388 -5494 2396 -5460
rect 2344 -5503 2396 -5494
rect 2681 -5477 2733 -5425
rect 2977 -5478 3029 -5426
rect 503 -5566 555 -5514
rect 1148 -5525 1200 -5507
rect 1148 -5559 1156 -5525
rect 1156 -5559 1190 -5525
rect 1190 -5559 1200 -5525
rect 869 -5572 921 -5563
rect 869 -5606 878 -5572
rect 878 -5606 912 -5572
rect 912 -5606 921 -5572
rect 869 -5615 921 -5606
rect 2681 -5570 2733 -5518
rect 3069 -5570 3121 -5518
rect 37 -5746 193 -5662
rect 3339 -5746 3495 -5662
<< metal2 >>
rect -147 -4030 9 -4024
rect -147 -5118 9 -4114
rect -147 -5752 9 -5202
rect 37 -4574 193 -4024
rect 37 -5662 193 -4658
rect 37 -5752 193 -5746
rect 221 -4159 285 -4024
rect 221 -4211 227 -4159
rect 279 -4211 285 -4159
rect 221 -4792 285 -4211
rect 221 -4844 227 -4792
rect 279 -4844 285 -4792
rect 221 -5266 285 -4844
rect 221 -5318 227 -5266
rect 279 -5318 285 -5266
rect 221 -5752 285 -5318
rect 313 -4215 377 -4024
rect 313 -4267 319 -4215
rect 371 -4267 377 -4215
rect 313 -4884 377 -4267
rect 313 -4936 319 -4884
rect 371 -4936 377 -4884
rect 313 -5345 377 -4936
rect 313 -5397 319 -5345
rect 371 -5397 377 -5345
rect 313 -5752 377 -5397
rect 405 -4271 469 -4024
rect 405 -4323 411 -4271
rect 463 -4323 469 -4271
rect 405 -4707 469 -4323
rect 405 -4759 411 -4707
rect 463 -4759 469 -4707
rect 405 -5422 469 -4759
rect 405 -5474 411 -5422
rect 463 -5474 469 -5422
rect 405 -5752 469 -5474
rect 497 -4369 561 -4024
rect 1051 -4250 1103 -4244
rect 1051 -4308 1103 -4302
rect 497 -4421 503 -4369
rect 555 -4421 561 -4369
rect 1075 -4363 1103 -4308
rect 1224 -4351 1276 -4345
rect 1886 -4347 1892 -4295
rect 1944 -4307 1950 -4295
rect 2787 -4307 2851 -4024
rect 1944 -4335 2851 -4307
rect 1944 -4347 1950 -4335
rect 1075 -4391 1224 -4363
rect 1224 -4409 1276 -4403
rect 2005 -4391 2595 -4363
rect 2005 -4407 2033 -4391
rect 497 -4947 561 -4421
rect 1969 -4459 1975 -4407
rect 2027 -4459 2033 -4407
rect 2589 -4415 2595 -4391
rect 2647 -4415 2653 -4363
rect 2523 -4460 2575 -4454
rect 2507 -4512 2523 -4475
rect 2507 -4518 2575 -4512
rect 2507 -4819 2535 -4518
rect 1044 -4835 1051 -4822
rect 757 -4863 1051 -4835
rect 757 -4947 785 -4863
rect 1044 -4874 1051 -4863
rect 1103 -4874 1109 -4822
rect 2481 -4871 2487 -4819
rect 2539 -4871 2545 -4819
rect 497 -4975 785 -4947
rect 497 -5514 561 -4975
rect 2787 -5026 2851 -4335
rect 2787 -5078 2793 -5026
rect 2845 -5078 2851 -5026
rect 645 -5240 1667 -5227
rect 645 -5255 1609 -5240
rect 645 -5415 673 -5255
rect 1603 -5292 1609 -5255
rect 1661 -5292 1667 -5240
rect 1737 -5255 2703 -5227
rect 1737 -5339 1765 -5255
rect 1093 -5367 1765 -5339
rect 1093 -5395 1121 -5367
rect 609 -5421 673 -5415
rect 609 -5473 615 -5421
rect 667 -5473 673 -5421
rect 851 -5447 857 -5395
rect 909 -5423 1121 -5395
rect 909 -5447 915 -5423
rect 1172 -5447 1178 -5395
rect 1230 -5423 2647 -5395
rect 1230 -5447 1236 -5423
rect 609 -5479 673 -5473
rect 1322 -5503 1328 -5451
rect 1380 -5479 2092 -5451
rect 1380 -5503 1386 -5479
rect 2086 -5503 2092 -5479
rect 2144 -5503 2150 -5451
rect 2186 -5503 2192 -5451
rect 2244 -5503 2250 -5451
rect 2338 -5475 2344 -5451
rect 2283 -5503 2344 -5475
rect 2396 -5503 2402 -5451
rect 497 -5566 503 -5514
rect 555 -5566 561 -5514
rect 1142 -5559 1148 -5507
rect 1200 -5531 1206 -5507
rect 2186 -5531 2214 -5503
rect 1200 -5559 2214 -5531
rect 497 -5752 561 -5566
rect 863 -5615 869 -5563
rect 921 -5587 928 -5563
rect 2283 -5587 2311 -5503
rect 2619 -5512 2647 -5423
rect 2675 -5419 2703 -5255
rect 2787 -5345 2851 -5078
rect 2787 -5397 2793 -5345
rect 2845 -5397 2851 -5345
rect 2675 -5425 2739 -5419
rect 2675 -5477 2681 -5425
rect 2733 -5477 2739 -5425
rect 2675 -5483 2739 -5477
rect 2619 -5518 2739 -5512
rect 2619 -5540 2681 -5518
rect 2675 -5570 2681 -5540
rect 2733 -5570 2739 -5518
rect 2675 -5576 2739 -5570
rect 921 -5615 2311 -5587
rect 2787 -5752 2851 -5397
rect 2879 -4159 2943 -4024
rect 2879 -4211 2885 -4159
rect 2937 -4211 2943 -4159
rect 2879 -4750 2943 -4211
rect 2879 -4802 2885 -4750
rect 2937 -4802 2943 -4750
rect 2879 -5253 2943 -4802
rect 2879 -5305 2885 -5253
rect 2937 -5305 2943 -5253
rect 2879 -5752 2943 -5305
rect 2971 -4315 3035 -4024
rect 2971 -4367 2977 -4315
rect 3029 -4367 3035 -4315
rect 2971 -5426 3035 -4367
rect 2971 -5478 2977 -5426
rect 3029 -5478 3035 -5426
rect 2971 -5752 3035 -5478
rect 3063 -4371 3127 -4024
rect 3063 -4423 3069 -4371
rect 3121 -4423 3127 -4371
rect 3063 -5518 3127 -4423
rect 3063 -5570 3069 -5518
rect 3121 -5570 3127 -5518
rect 3063 -5752 3127 -5570
rect 3155 -4030 3311 -4024
rect 3155 -5118 3311 -4114
rect 3155 -5752 3311 -5202
rect 3339 -4574 3495 -4024
rect 3339 -5662 3495 -4658
rect 3339 -5752 3495 -5746
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1749714889
transform 1 0 1956 0 -1 -4616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1749714889
transform 1 0 2416 0 -1 -4616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1749714889
transform 1 0 1496 0 1 -4616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1749714889
transform 1 0 2416 0 1 -5704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1864 0 1 -4616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1704896540
transform 1 0 2232 0 -1 -4616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1704896540
transform 1 0 2324 0 -1 -4616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1704896540
transform 1 0 2692 0 1 -5704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1704896540
transform 1 0 576 0 1 -5704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1704896540
transform 1 0 576 0 1 -4616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1704896540
transform 1 0 576 0 -1 -4616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1704896540
transform 1 0 2692 0 -1 -4616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1704896540
transform 1 0 2692 0 1 -4616
box -38 -48 130 592
use seg_selector_1_logic  x1
timestamp 1749667264
transform 1 0 1234 0 1 -2656
box 592 -2008 1496 -1368
use seg_selector_2_logic  x2
timestamp 1749736748
transform 1 0 131 0 1 -2259
box 499 -3493 2323 -2853
use seg_selector_3_logic  x3
timestamp 1749714889
transform 1 0 -62 0 -1 -6976
box 692 -2408 2056 -1768
use seg_selector_4_logic  x4
timestamp 1749664768
transform 1 0 380 0 1 -2402
box 250 -2262 1154 -1622
<< labels >>
flabel metal2 s 221 -4024 221 -4024 4 FreeSans 240 0 0 0 b[6]
port 0 se
flabel metal2 s 313 -4024 313 -4024 4 FreeSans 240 0 0 0 b[7]
port 1 se
flabel metal2 s 405 -4024 405 -4024 4 FreeSans 240 0 0 0 b[8]
port 2 se
flabel metal2 s 497 -4024 497 -4024 4 FreeSans 240 0 0 0 b[9]
port 3 se
flabel metal2 s 2787 -4024 2787 -4024 4 FreeSans 240 0 0 0 bb[6]
port 4 se
flabel metal2 s 2879 -4024 2879 -4024 4 FreeSans 240 0 0 0 bb[7]
port 5 se
flabel metal2 s 2971 -4024 2971 -4024 4 FreeSans 240 0 0 0 bb[8]
port 6 se
flabel metal2 s 3063 -4024 3063 -4024 4 FreeSans 240 0 0 0 bb[9]
port 7 se
flabel metal2 s 2514 -4807 2514 -4807 4 FreeSans 240 0 0 0 S[1]
port 8 se
flabel metal1 s 2433 -5465 2433 -5465 4 FreeSans 240 0 0 0 S[2]
port 9 se
flabel metal1 s 1953 -4752 1953 -4752 4 FreeSans 240 0 0 0 S[3]
port 10 se
flabel metal1 s 1482 -4271 1482 -4271 4 FreeSans 240 0 0 0 S[4]
port 11 se
flabel locali s 2584 -4875 2584 -4875 4 FreeSans 240 0 0 0 SB[1]
port 12 se
flabel locali s 2582 -5449 2582 -5449 4 FreeSans 240 0 0 0 SB[2]
port 13 se
flabel locali s 2123 -4822 2123 -4822 4 FreeSans 240 0 0 0 SB[3]
port 14 se
flabel locali s 1664 -4350 1664 -4350 4 FreeSans 240 0 0 0 SB[4]
port 15 se
flabel metal2 s -145 -4027 -145 -4027 4 FreeSans 480 0 0 0 VDD
port 16 se
flabel metal2 s 39 -4026 39 -4026 4 FreeSans 480 0 0 0 GND
port 17 se
<< end >>
