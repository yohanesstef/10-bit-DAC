magic
tech sky130A
magscale 1 2
timestamp 1750052349
<< mvnsubdiffcont >>
rect -90 602 8998 636
rect -150 -488 -116 576
rect 9024 -488 9058 576
rect -150 -522 9058 -488
rect -150 -1586 -116 -522
rect 9024 -1586 9058 -522
rect -90 -1646 8998 -1612
<< metal1 >>
rect 4361 -221 4421 -215
rect 4361 -287 4421 -281
rect 4487 -221 4547 -215
rect 4487 -287 4547 -281
rect 4284 -978 4380 -918
rect 4536 -978 4624 -918
rect 4284 -1081 4344 -978
rect 4284 -1147 4344 -1141
rect 4564 -1169 4624 -978
rect 4564 -1235 4624 -1229
<< via1 >>
rect 4361 -281 4421 -221
rect 4487 -281 4547 -221
rect 4284 -1141 4344 -1081
rect 4564 -1229 4624 -1169
<< metal2 >>
rect 3849 493 3859 549
rect 3915 493 3925 549
rect 1034 393 7122 395
rect 1034 337 4237 393
rect 4293 337 7122 393
rect 1034 335 7122 337
rect 1786 305 7874 307
rect 1786 249 4111 305
rect 4167 249 7874 305
rect 1786 247 7874 249
rect 2162 41 7498 43
rect 2162 -15 3985 41
rect 4041 -15 7498 41
rect 2162 -17 7498 -15
rect 717 -47 8191 -45
rect 717 -103 4867 -47
rect 4923 -103 8191 -47
rect 717 -105 8191 -103
rect 3666 -135 5994 -133
rect 3666 -191 4741 -135
rect 4797 -191 5994 -135
rect 3666 -193 5994 -191
rect 4354 -281 4361 -221
rect 4421 -281 4428 -221
rect 4480 -281 4487 -221
rect 4547 -281 4554 -221
rect 4606 -223 5242 -221
rect 4606 -279 4615 -223
rect 4671 -279 5242 -223
rect 4606 -281 5242 -279
rect 3849 -435 3859 -379
rect 3915 -435 3925 -379
rect 3849 -631 3859 -575
rect 3915 -631 3925 -575
rect 3666 -731 4680 -729
rect 3666 -787 4615 -731
rect 4671 -787 4680 -731
rect 3666 -789 4680 -787
rect 2914 -819 5242 -817
rect 2914 -875 4741 -819
rect 4797 -875 5242 -819
rect 2914 -877 5242 -875
rect 717 -907 8191 -905
rect 717 -963 4867 -907
rect 4923 -963 8191 -907
rect 717 -965 8191 -963
rect 1410 -995 6746 -993
rect 1410 -1051 3985 -995
rect 4041 -1051 6746 -995
rect 1410 -1053 6746 -1051
rect 4278 -1141 4284 -1081
rect 4344 -1083 4554 -1081
rect 4344 -1139 4489 -1083
rect 4545 -1139 4554 -1083
rect 4344 -1141 4554 -1139
rect 4354 -1171 4564 -1169
rect 4354 -1227 4363 -1171
rect 4419 -1227 4564 -1171
rect 4354 -1229 4564 -1227
rect 4624 -1229 4630 -1169
rect 1034 -1259 7122 -1257
rect 1034 -1315 4111 -1259
rect 4167 -1315 7122 -1259
rect 1034 -1317 7122 -1315
rect 1786 -1347 7874 -1345
rect 1786 -1403 4237 -1347
rect 4293 -1403 7874 -1347
rect 1786 -1405 7874 -1403
rect 3849 -1559 3859 -1503
rect 3915 -1559 3925 -1503
<< via2 >>
rect 3859 493 3915 549
rect 4237 337 4293 393
rect 4111 249 4167 305
rect 3985 -15 4041 41
rect 4867 -103 4923 -47
rect 4741 -191 4797 -135
rect 4363 -279 4419 -223
rect 4489 -279 4545 -223
rect 4615 -279 4671 -223
rect 3859 -435 3915 -379
rect 3859 -631 3915 -575
rect 4615 -787 4671 -731
rect 4741 -875 4797 -819
rect 4867 -963 4923 -907
rect 3985 -1051 4041 -995
rect 4489 -1139 4545 -1083
rect 4363 -1227 4419 -1171
rect 4111 -1315 4167 -1259
rect 4237 -1403 4293 -1347
rect 3859 -1559 3915 -1503
<< metal3 >>
rect 3854 549 3920 559
rect 3854 493 3859 549
rect 3915 493 3920 549
rect 3854 -379 3920 493
rect 4232 393 4298 403
rect 4232 337 4237 393
rect 4293 337 4298 393
rect 4106 305 4172 315
rect 4106 249 4111 305
rect 4167 249 4172 305
rect 3854 -435 3859 -379
rect 3915 -435 3920 -379
rect 3854 -575 3920 -435
rect 3854 -631 3859 -575
rect 3915 -631 3920 -575
rect 3854 -1503 3920 -631
rect 3854 -1559 3859 -1503
rect 3915 -1559 3920 -1503
rect 3854 -1659 3920 -1559
rect 3980 41 4046 51
rect 3980 -15 3985 41
rect 4041 -15 4046 41
rect 3980 -995 4046 -15
rect 3980 -1051 3985 -995
rect 4041 -1051 4046 -995
rect 3980 -1659 4046 -1051
rect 4106 -1259 4172 249
rect 4106 -1315 4111 -1259
rect 4167 -1315 4172 -1259
rect 4106 -1659 4172 -1315
rect 4232 -1347 4298 337
rect 4862 -47 4928 -37
rect 4862 -103 4867 -47
rect 4923 -103 4928 -47
rect 4736 -135 4802 -125
rect 4736 -191 4741 -135
rect 4797 -191 4802 -135
rect 4232 -1403 4237 -1347
rect 4293 -1403 4298 -1347
rect 4232 -1659 4298 -1403
rect 4358 -223 4424 -213
rect 4358 -279 4363 -223
rect 4419 -279 4424 -223
rect 4358 -1171 4424 -279
rect 4358 -1227 4363 -1171
rect 4419 -1227 4424 -1171
rect 4358 -1659 4424 -1227
rect 4484 -223 4550 -213
rect 4484 -279 4489 -223
rect 4545 -279 4550 -223
rect 4484 -1083 4550 -279
rect 4484 -1139 4489 -1083
rect 4545 -1139 4550 -1083
rect 4484 -1659 4550 -1139
rect 4610 -223 4676 -211
rect 4610 -279 4615 -223
rect 4671 -279 4676 -223
rect 4610 -731 4676 -279
rect 4610 -787 4615 -731
rect 4671 -787 4676 -731
rect 4610 -1659 4676 -787
rect 4736 -819 4802 -191
rect 4736 -875 4741 -819
rect 4797 -875 4802 -819
rect 4736 -1659 4802 -875
rect 4862 -907 4928 -103
rect 4862 -963 4867 -907
rect 4923 -963 4928 -907
rect 4862 -1659 4928 -963
use cm_pcell1_left  cm_pcell1_left_0
timestamp 1749890363
transform 1 0 -116 0 1 -588
box -112 -14 4652 1304
use cm_pcell1_left  cm_pcell1_left_1
timestamp 1749890363
transform -1 0 9024 0 -1 -422
box -112 -14 4652 1304
use cm_pcell1_right  cm_pcell1_right_0
timestamp 1749890363
transform 1 0 -498 0 1 -2147
box 4870 1545 9634 2863
use cm_pcell1_right  cm_pcell1_right_1
timestamp 1749890363
transform -1 0 9406 0 -1 1137
box 4870 1545 9634 2863
<< labels >>
flabel metal3 s 3854 -1659 3854 -1659 2 FreeSans 320 0 0 0 G1
port 0 ne
flabel metal3 s 4232 -1659 4232 -1659 2 FreeSans 320 0 0 0 io0
port 1 ne
flabel metal3 s 4106 -1659 4106 -1659 2 FreeSans 320 0 0 0 io1
port 2 ne
flabel metal3 s 3980 -1659 3980 -1659 2 FreeSans 320 0 0 0 io2
port 3 ne
flabel metal3 s 4358 -1659 4358 -1659 2 FreeSans 320 0 0 0 ho0
port 4 ne
flabel metal3 s 4484 -1659 4484 -1659 2 FreeSans 320 0 0 0 ho1
port 5 ne
flabel metal3 s 4610 -1659 4610 -1659 2 FreeSans 320 0 0 0 ho2
port 6 ne
flabel metal3 s 4736 -1659 4736 -1659 2 FreeSans 320 0 0 0 ho3
port 7 ne
flabel metal3 s 4862 -1659 4862 -1659 2 FreeSans 320 0 0 0 ho4
port 8 ne
flabel metal1 s 3589 -1669 3589 -1669 2 FreeSans 480 0 0 0 VDDA
port 9 ne
<< end >>
