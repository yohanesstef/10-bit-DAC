magic
tech sky130A
magscale 1 2
timestamp 1750066786
<< error_p >>
rect -353 -398 -323 330
rect -287 -332 -257 264
rect 257 -332 287 264
rect -287 -336 287 -332
rect 323 -398 353 330
rect -353 -402 353 -398
<< nwell >>
rect -323 -398 323 364
<< mvpmos >>
rect -229 -336 -29 264
rect 29 -336 229 264
<< mvpdiff >>
rect -287 252 -229 264
rect -287 -324 -275 252
rect -241 -324 -229 252
rect -287 -336 -229 -324
rect -29 252 29 264
rect -29 -324 -17 252
rect 17 -324 29 252
rect -29 -336 29 -324
rect 229 252 287 264
rect 229 -324 241 252
rect 275 -324 287 252
rect 229 -336 287 -324
<< mvpdiffc >>
rect -275 -324 -241 252
rect -17 -324 17 252
rect 241 -324 275 252
<< poly >>
rect -229 345 -29 361
rect -229 311 -213 345
rect -45 311 -29 345
rect -229 264 -29 311
rect 29 345 229 361
rect 29 311 45 345
rect 213 311 229 345
rect 29 264 229 311
rect -229 -362 -29 -336
rect 29 -362 229 -336
<< polycont >>
rect -213 311 -45 345
rect 45 311 213 345
<< locali >>
rect -229 311 -213 345
rect -45 311 -29 345
rect 29 311 45 345
rect 213 311 229 345
rect -275 252 -241 268
rect -275 -340 -241 -324
rect -17 252 17 268
rect -17 -340 17 -324
rect 241 252 275 268
rect 241 -340 275 -324
<< viali >>
rect -192 311 -66 345
rect 66 311 192 345
rect -275 -324 -241 252
rect -17 -324 17 252
rect 241 -324 275 252
<< metal1 >>
rect -204 345 -54 351
rect -204 311 -192 345
rect -66 311 -54 345
rect -204 305 -54 311
rect 54 345 204 351
rect 54 311 66 345
rect 192 311 204 345
rect 54 305 204 311
rect -281 252 -235 264
rect -281 -324 -275 252
rect -241 -324 -235 252
rect -281 -336 -235 -324
rect -23 252 23 264
rect -23 -324 -17 252
rect 17 -324 23 252
rect -23 -336 23 -324
rect 235 252 281 264
rect 235 -324 241 252
rect 275 -324 281 252
rect 235 -336 281 -324
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
