magic
tech sky130A
magscale 1 2
timestamp 1751047404
<< error_s >>
rect 2358 3706 2380 3734
rect 2386 3678 2408 3744
rect 2358 3457 2380 3485
rect 2386 3429 2408 3513
rect 2358 3208 2380 3236
rect 2386 3180 2408 3264
rect 2612 3082 2680 3098
rect 2596 3081 2696 3082
rect 2585 3054 2707 3060
rect 2562 3047 2730 3048
<< nwell >>
rect 2160 3208 2180 3236
<< metal1 >>
rect -252 4206 -200 4216
rect -252 4148 -200 4154
rect 174 4206 226 4216
rect 174 4148 226 4154
rect 1520 4206 1572 4216
rect 1520 4148 1572 4154
rect 1946 4206 1998 4216
rect 1946 4148 1998 4154
rect -252 3966 -200 3976
rect -252 3908 -200 3914
rect 174 3966 226 3976
rect 1520 3966 1572 3976
rect 382 3928 608 3956
rect 174 3908 226 3914
rect 1520 3908 1572 3914
rect 1946 3966 1998 3976
rect 1946 3908 1998 3914
rect -252 3726 -200 3736
rect -252 3668 -200 3674
rect 174 3726 226 3736
rect 1520 3726 1572 3736
rect 382 3688 608 3716
rect 174 3668 226 3674
rect 1520 3668 1572 3674
rect 1946 3726 1998 3736
rect 2154 3706 2380 3734
rect 1946 3668 1998 3674
rect -252 3486 -200 3496
rect -252 3428 -200 3434
rect 174 3486 226 3496
rect 1520 3486 1572 3496
rect 382 3448 608 3476
rect 174 3428 226 3434
rect 1520 3428 1572 3434
rect 1946 3486 1998 3496
rect 2154 3457 2380 3485
rect 1946 3428 1998 3434
rect -252 3246 -200 3256
rect -252 3188 -200 3194
rect 174 3246 226 3256
rect 1520 3246 1572 3256
rect 382 3208 608 3236
rect 174 3188 226 3194
rect 1520 3188 1572 3194
rect 1946 3246 1998 3256
rect 2160 3208 2380 3236
rect 1946 3188 1998 3194
<< via1 >>
rect -252 4154 -200 4206
rect 174 4154 226 4206
rect 1520 4154 1572 4206
rect 1946 4154 1998 4206
rect -252 3914 -200 3966
rect 174 3914 226 3966
rect 1520 3914 1572 3966
rect 1946 3914 1998 3966
rect -252 3674 -200 3726
rect 174 3674 226 3726
rect 1520 3674 1572 3726
rect 1946 3674 1998 3726
rect -252 3434 -200 3486
rect 174 3434 226 3486
rect 1520 3434 1572 3486
rect 1946 3434 1998 3486
rect -252 3194 -200 3246
rect 174 3194 226 3246
rect 1520 3194 1572 3246
rect 1946 3194 1998 3246
<< metal2 >>
rect -252 4210 -196 4220
rect -252 4144 -196 4154
rect 174 4210 230 4220
rect 174 4144 230 4154
rect 1520 4210 1576 4220
rect 1520 4144 1576 4154
rect 1946 4210 2002 4220
rect 1946 4144 2002 4154
rect -252 3970 -196 3980
rect -252 3904 -196 3914
rect 174 3970 230 3980
rect 174 3904 230 3914
rect 1520 3970 1576 3980
rect 1520 3904 1576 3914
rect 1946 3970 2002 3980
rect 1946 3904 2002 3914
rect -252 3730 -196 3740
rect -252 3664 -196 3674
rect 174 3730 230 3740
rect 174 3664 230 3674
rect 1520 3730 1576 3740
rect 1520 3664 1576 3674
rect 1946 3730 2002 3740
rect 1946 3664 2002 3674
rect -252 3490 -196 3500
rect -252 3424 -196 3434
rect 174 3490 230 3500
rect 174 3424 230 3434
rect 1520 3490 1576 3500
rect 1520 3424 1576 3434
rect 1946 3490 2002 3500
rect 1946 3424 2002 3434
rect -252 3250 -196 3260
rect -252 3184 -196 3194
rect 174 3250 230 3260
rect 174 3184 230 3194
rect 1520 3250 1576 3260
rect 1520 3184 1576 3194
rect 1946 3250 2002 3260
rect 1946 3184 2002 3194
<< via2 >>
rect -252 4206 -196 4210
rect -252 4154 -200 4206
rect -200 4154 -196 4206
rect 174 4206 230 4210
rect 174 4154 226 4206
rect 226 4154 230 4206
rect 1520 4206 1576 4210
rect 1520 4154 1572 4206
rect 1572 4154 1576 4206
rect 1946 4206 2002 4210
rect 1946 4154 1998 4206
rect 1998 4154 2002 4206
rect -252 3966 -196 3970
rect -252 3914 -200 3966
rect -200 3914 -196 3966
rect 174 3966 230 3970
rect 174 3914 226 3966
rect 226 3914 230 3966
rect 1520 3966 1576 3970
rect 1520 3914 1572 3966
rect 1572 3914 1576 3966
rect 1946 3966 2002 3970
rect 1946 3914 1998 3966
rect 1998 3914 2002 3966
rect -252 3726 -196 3730
rect -252 3674 -200 3726
rect -200 3674 -196 3726
rect 174 3726 230 3730
rect 174 3674 226 3726
rect 226 3674 230 3726
rect 1520 3726 1576 3730
rect 1520 3674 1572 3726
rect 1572 3674 1576 3726
rect 1946 3726 2002 3730
rect 1946 3674 1998 3726
rect 1998 3674 2002 3726
rect -252 3486 -196 3490
rect -252 3434 -200 3486
rect -200 3434 -196 3486
rect 174 3486 230 3490
rect 174 3434 226 3486
rect 226 3434 230 3486
rect 1520 3486 1576 3490
rect 1520 3434 1572 3486
rect 1572 3434 1576 3486
rect 1946 3486 2002 3490
rect 1946 3434 1998 3486
rect 1998 3434 2002 3486
rect -252 3246 -196 3250
rect -252 3194 -200 3246
rect -200 3194 -196 3246
rect 174 3246 230 3250
rect 174 3194 226 3246
rect 226 3194 230 3246
rect 1520 3246 1576 3250
rect 1520 3194 1572 3246
rect 1572 3194 1576 3246
rect 1946 3246 2002 3250
rect 1946 3194 1998 3246
rect 1998 3194 2002 3246
<< metal3 >>
rect -262 4210 2012 4215
rect -262 4154 -252 4210
rect -196 4154 174 4210
rect 230 4154 1520 4210
rect 1576 4154 1946 4210
rect 2002 4154 2012 4210
rect -262 4149 2012 4154
rect -262 3970 2012 3975
rect -262 3914 -252 3970
rect -196 3914 174 3970
rect 230 3914 1520 3970
rect 1576 3914 1946 3970
rect 2002 3914 2012 3970
rect -262 3909 2012 3914
rect -262 3730 2012 3735
rect -262 3674 -252 3730
rect -196 3674 174 3730
rect 230 3674 1520 3730
rect 1576 3674 1946 3730
rect 2002 3674 2012 3730
rect -262 3669 2012 3674
rect -262 3490 2012 3495
rect -262 3434 -252 3490
rect -196 3434 174 3490
rect 230 3434 1520 3490
rect 1576 3434 1946 3490
rect 2002 3434 2012 3490
rect -262 3429 2012 3434
rect -262 3250 2012 3255
rect -262 3194 -252 3250
rect -196 3194 174 3250
rect 230 3194 1520 3250
rect 1576 3194 1946 3250
rect 2002 3194 2012 3250
rect -262 3189 2012 3194
use interpolation_s2  interpolation_s2_0
timestamp 1751042016
transform 1 0 585 0 1 3118
box -151 -134 689 1279
use interpolation_s3  interpolation_s3_0
timestamp 1751042016
transform 1 0 2357 0 1 3100
box -181 -164 719 1105
use interpolation_switch  interpolation_switch_0
timestamp 1751047215
transform 1 0 559 0 1 5062
box -188 -172 1374 1062
use seg_sel_1  seg_sel_1_0
timestamp 1750845293
transform 1 0 -351 0 1 3052
box -67 -68 489 1430
use seg_sel_2  seg_sel_2_0
timestamp 1750845353
transform 1 0 87 0 1 3058
box -79 -74 477 1424
use seg_sel_3  seg_sel_3_0
timestamp 1750845438
transform 1 0 1846 0 1 3045
box -96 -109 520 1495
use seg_sel_4  seg_sel_4_0
timestamp 1750845534
transform 1 0 1420 0 1 3041
box -96 -105 520 1499
use seg_sel_nmos  seg_sel_nmos_0
timestamp 1751047180
transform 1 0 701 0 1 5081
box -930 -169 -200 1309
use seg_sel_pmos  seg_sel_pmos_0
timestamp 1751047404
transform 1 0 -4488 0 1 4596
box 6231 294 7013 1813
<< end >>
