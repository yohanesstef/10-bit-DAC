magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1217 307 1217
<< psubdiff >>
rect -271 1147 -175 1181
rect 175 1147 271 1181
rect -271 1085 -237 1147
rect 237 1085 271 1147
rect -271 -1147 -237 -1085
rect 237 -1147 271 -1085
rect -271 -1181 -175 -1147
rect 175 -1181 271 -1147
<< psubdiffcont >>
rect -175 1147 175 1181
rect -271 -1085 -237 1085
rect 237 -1085 271 1085
rect -175 -1181 175 -1147
<< xpolycontact >>
rect -141 619 141 1051
rect -141 -1051 141 -619
<< xpolyres >>
rect -141 -619 141 619
<< locali >>
rect -271 1147 -175 1181
rect 175 1147 271 1181
rect -271 1085 -237 1147
rect 237 1085 271 1147
rect -271 -1147 -237 -1085
rect 237 -1147 271 -1085
rect -271 -1181 -175 -1147
rect 175 -1181 271 -1147
<< viali >>
rect -125 636 125 1033
rect -125 -1033 125 -636
<< metal1 >>
rect -131 1033 131 1045
rect -131 636 -125 1033
rect 125 636 131 1033
rect -131 624 131 636
rect -131 -636 131 -624
rect -131 -1033 -125 -636
rect 125 -1033 131 -636
rect -131 -1045 131 -1033
<< properties >>
string FIXED_BBOX -254 -1164 254 1164
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 6.346 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 9.268k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
