magic
tech sky130A
magscale 1 2
timestamp 1749147327
<< xpolycontact >>
rect -141 239 141 671
rect -141 -671 141 -239
<< xpolyres >>
rect -141 -239 141 239
<< viali >>
rect -125 256 125 653
rect -125 -653 125 -256
<< metal1 >>
rect -131 653 131 665
rect -131 256 -125 653
rect 125 256 131 653
rect -131 244 131 256
rect -131 -256 131 -244
rect -131 -653 -125 -256
rect 125 -653 131 -256
rect -131 -665 131 -653
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 2.553 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 3.888k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
