magic
tech sky130A
magscale 1 2
timestamp 1749548291
<< error_s >>
rect 1074 684 1080 690
rect 1128 684 1134 690
rect 1068 678 1074 684
rect 1134 678 1140 684
rect 1068 624 1074 630
rect 1134 624 1140 630
rect 1074 618 1080 624
rect 1128 618 1134 624
rect 798 596 804 602
rect 852 596 858 602
rect 792 590 798 596
rect 858 590 864 596
rect 792 536 798 542
rect 858 536 864 542
rect 798 530 804 536
rect 852 530 858 536
rect 522 508 528 514
rect 576 508 582 514
rect 516 502 522 508
rect 582 502 588 508
rect 516 448 522 454
rect 582 448 588 454
rect 522 442 528 448
rect 576 442 582 448
rect 246 420 252 426
rect 300 420 306 426
rect 240 414 246 420
rect 306 414 312 420
rect 240 360 246 366
rect 306 360 312 366
rect 246 354 252 360
rect 300 354 306 360
rect 891 -45 897 -39
rect 945 -45 951 -39
rect 885 -51 891 -45
rect 951 -51 957 -45
rect 885 -105 891 -99
rect 951 -105 957 -99
rect 891 -111 897 -105
rect 945 -111 951 -105
rect 615 -133 621 -127
rect 669 -133 675 -127
rect 609 -139 615 -133
rect 675 -139 681 -133
rect 609 -193 615 -187
rect 675 -193 681 -187
rect 615 -199 621 -193
rect 669 -199 675 -193
rect 339 -221 345 -215
rect 393 -221 399 -215
rect 333 -227 339 -221
rect 399 -227 405 -221
rect 333 -281 339 -275
rect 399 -281 405 -275
rect 339 -287 345 -281
rect 393 -287 399 -281
rect 63 -309 69 -303
rect 117 -309 123 -303
rect 57 -315 63 -309
rect 123 -315 129 -309
rect 57 -369 63 -363
rect 123 -369 129 -363
rect 63 -375 69 -369
rect 117 -375 123 -369
<< metal1 >>
rect 1074 684 1134 690
rect 798 596 858 602
rect 522 508 582 514
rect 246 420 306 426
rect 246 70 306 360
rect 522 70 582 448
rect 63 -309 123 70
rect 339 -221 399 70
rect 615 -133 675 71
rect 798 70 858 536
rect 1074 70 1134 624
rect 891 -45 951 70
rect 891 -111 951 -105
rect 615 -199 675 -193
rect 339 -287 399 -281
rect 63 -375 123 -369
<< via1 >>
rect 1074 624 1134 684
rect 798 536 858 596
rect 522 448 582 508
rect 246 360 306 420
rect 891 -105 951 -45
rect 615 -193 675 -133
rect 339 -281 399 -221
rect 63 -369 123 -309
use hnmos_4  hnmos_4_0
timestamp 1749548291
transform 1 0 42 0 1 44
box -8 0 1096 198
<< end >>
