magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -714 307 714
<< psubdiff >>
rect -271 644 -175 678
rect 175 644 271 678
rect -271 582 -237 644
rect 237 582 271 644
rect -271 -644 -237 -582
rect 237 -644 271 -582
rect -271 -678 -175 -644
rect 175 -678 271 -644
<< psubdiffcont >>
rect -175 644 175 678
rect -271 -582 -237 582
rect 237 -582 271 582
rect -175 -678 175 -644
<< xpolycontact >>
rect -141 116 141 548
rect -141 -548 141 -116
<< xpolyres >>
rect -141 -116 141 116
<< locali >>
rect -271 644 -175 678
rect 175 644 271 678
rect -271 582 -237 644
rect 237 582 271 644
rect -271 -644 -237 -582
rect 237 -644 271 -582
rect -271 -678 -175 -644
rect 175 -678 271 -644
<< viali >>
rect -125 133 125 530
rect -125 -530 125 -133
<< metal1 >>
rect -131 530 131 542
rect -131 133 -125 530
rect 125 133 131 530
rect -131 121 131 133
rect -131 -133 131 -121
rect -131 -530 -125 -133
rect 125 -530 131 -133
rect -131 -542 131 -530
<< properties >>
string FIXED_BBOX -254 -661 254 661
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.323 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 2.143k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
