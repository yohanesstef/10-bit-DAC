magic
tech sky130A
magscale 1 2
timestamp 1750017183
<< mvpsubdiff >>
rect -374 1313 1184 1373
rect -374 578 -314 1313
rect 1124 578 1184 1313
<< poly >>
rect -16 670 44 1104
rect 766 670 826 1104
<< locali >>
rect -361 1326 1171 1360
rect -361 578 -327 1326
rect 1137 578 1171 1326
<< metal1 >>
rect -280 1103 -220 1109
rect -280 578 -220 1043
rect -192 578 -132 1285
rect 148 1043 154 1103
rect 280 1043 286 1103
rect 323 1016 369 1121
rect 441 1016 487 1121
rect 524 1043 530 1103
rect 656 1043 662 1103
rect 942 578 1002 1285
<< via1 >>
rect -280 1043 -220 1103
rect 154 1043 280 1103
rect 530 1043 656 1103
<< metal2 >>
rect -286 1043 -280 1103
rect -220 1043 154 1103
rect 280 1043 530 1103
rect 656 1043 662 1103
use sky130_fd_pr__nfet_g5v0d10v5_YZ2SRG  sky130_fd_pr__nfet_g5v0d10v5_YZ2SRG_0
timestamp 1750017183
transform 1 0 217 0 1 887
box -158 -217 158 217
use sky130_fd_pr__nfet_g5v0d10v5_YZ2SRG  sky130_fd_pr__nfet_g5v0d10v5_YZ2SRG_1
timestamp 1750017183
transform 1 0 593 0 1 887
box -158 -217 158 217
<< end >>
