magic
tech sky130A
magscale 1 2
timestamp 1749485587
<< metal1 >>
rect 18462 -23125 18522 -21181
rect 18550 -22476 18610 -21181
rect 18638 -21828 18698 -21181
rect 18726 -21505 18865 -21180
rect 18638 -22153 18865 -21828
rect 18550 -22801 18865 -22476
rect 18462 -23449 18865 -23125
<< end >>
