magic
tech sky130A
magscale 1 2
timestamp 1750150351
<< nwell >>
rect 3009 -235 4699 2767
<< mvnsubdiffcont >>
rect 3148 2654 4560 2688
rect 3088 -96 3122 2628
rect 4586 -96 4620 2628
rect 3148 -156 4560 -122
<< metal1 >>
rect 4303 2607 4363 2613
rect 3759 2547 3765 2607
rect 3825 2547 3831 2607
rect 3345 2519 3405 2525
rect 3169 95 3229 2437
rect 3257 1236 3317 1242
rect 3257 13 3317 1176
rect 3345 73 3405 2459
rect 3772 2454 3818 2547
rect 3877 2459 3883 2519
rect 3943 2459 3949 2519
rect 3890 2454 3936 2459
rect 3514 1356 3560 1384
rect 4148 1356 4194 1384
rect 3514 1296 3725 1356
rect 3999 1296 4194 1356
rect 3514 1176 3520 1236
rect 3580 1176 3710 1236
rect 3941 1176 4128 1236
rect 4188 1176 4194 1236
rect 3514 1148 3560 1176
rect 4148 1136 4194 1176
rect 3772 73 3818 79
rect 3345 13 3818 73
rect 3890 73 3936 78
rect 4303 73 4363 2547
rect 3890 13 4363 73
rect 4391 1236 4451 1242
rect 4391 13 4451 1176
<< via1 >>
rect 3765 2547 3825 2607
rect 4303 2547 4363 2607
rect 3345 2459 3405 2519
rect 3257 1176 3317 1236
rect 3883 2459 3943 2519
rect 3520 1176 3580 1236
rect 4128 1176 4188 1236
rect 4391 1176 4451 1236
<< metal2 >>
rect 3759 2547 3765 2607
rect 3825 2547 4303 2607
rect 4363 2547 4369 2607
rect 3339 2459 3345 2519
rect 3405 2459 3883 2519
rect 3943 2459 3949 2519
rect 3251 1176 3257 1236
rect 3317 1176 3520 1236
rect 3580 1176 3586 1236
rect 4122 1176 4128 1236
rect 4188 1176 4391 1236
rect 4451 1176 4457 1236
use cross_pair  cross_pair_0
timestamp 1750150351
transform 1 0 -32404 0 1 -679
box 36114 1855 36403 2035
use monticelli_pmos_2  monticelli_pmos_2_0
timestamp 1750003173
transform 1 0 3449 0 1 1328
box -440 -128 1250 1439
use monticelli_pmos_2  monticelli_pmos_2_1
timestamp 1750003173
transform 1 0 3449 0 -1 1204
box -440 -128 1250 1439
<< end >>
