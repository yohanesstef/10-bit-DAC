magic
tech sky130A
magscale 1 2
timestamp 1743275510
<< pwell >>
rect -201 -663 201 663
<< psubdiff >>
rect -165 593 -69 627
rect 69 593 165 627
rect -165 531 -131 593
rect 131 531 165 593
rect -165 -593 -131 -531
rect 131 -593 165 -531
rect -165 -627 -69 -593
rect 69 -627 165 -593
<< psubdiffcont >>
rect -69 593 69 627
rect -165 -531 -131 531
rect 131 -531 165 531
rect -69 -627 69 -593
<< xpolycontact >>
rect -35 65 35 497
rect -35 -497 35 -65
<< xpolyres >>
rect -35 -65 35 65
<< locali >>
rect -165 593 -69 627
rect 69 593 165 627
rect -165 531 -131 593
rect 131 531 165 593
rect -165 -593 -131 -531
rect 131 -593 165 -531
rect -165 -627 -69 -593
rect 69 -627 165 -593
<< viali >>
rect -19 82 19 479
rect -19 -479 19 -82
<< metal1 >>
rect -25 479 25 491
rect -25 82 -19 479
rect 19 82 25 479
rect -25 70 25 82
rect -25 -82 25 -70
rect -25 -479 -19 -82
rect 19 -479 25 -82
rect -25 -491 25 -479
<< properties >>
string FIXED_BBOX -148 -610 148 610
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.812 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 5.715k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
