magic
tech sky130A
magscale 1 2
timestamp 1750058993
<< mvnmos >>
rect -100 -91 100 29
<< mvndiff >>
rect -158 17 -100 29
rect -158 -79 -146 17
rect -112 -79 -100 17
rect -158 -91 -100 -79
rect 100 17 158 29
rect 100 -79 112 17
rect 146 -79 158 17
rect 100 -91 158 -79
<< mvndiffc >>
rect -146 -79 -112 17
rect 112 -79 146 17
<< poly >>
rect -100 101 100 117
rect -100 67 -84 101
rect 84 67 100 101
rect -100 29 100 67
rect -100 -117 100 -91
<< polycont >>
rect -84 67 84 101
<< locali >>
rect -100 67 -84 101
rect 84 67 100 101
rect -146 17 -112 33
rect -146 -95 -112 -79
rect 112 17 146 33
rect 112 -95 146 -79
<< viali >>
rect -63 67 63 101
rect -146 -79 -112 17
rect 112 -79 146 17
<< metal1 >>
rect -75 101 75 107
rect -75 67 -63 101
rect 63 67 75 101
rect -75 61 75 67
rect -152 17 -106 29
rect -152 -79 -146 17
rect -112 -79 -106 17
rect -152 -91 -106 -79
rect 106 17 152 29
rect 106 -79 112 17
rect 146 -79 152 17
rect 106 -91 152 -79
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.6 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
