magic
tech sky130A
magscale 1 2
timestamp 1749915489
<< error_s >>
rect -555 957 1365 1023
rect -555 79 -489 957
rect -429 831 1239 897
rect -429 79 -363 831
rect -555 13 -363 79
rect -206 17 -176 745
rect -140 83 -110 679
rect 920 83 950 679
rect -140 79 950 83
rect 986 17 1016 745
rect -206 13 1016 17
rect 1173 79 1239 831
rect 1299 79 1365 957
rect 1173 13 1365 79
<< mvnsubdiff >>
rect -489 897 1299 957
rect -489 79 -429 897
rect 1239 79 1299 897
<< poly >>
rect -215 53 -155 776
rect 965 53 1025 776
<< locali >>
rect -476 910 1286 944
rect -476 79 -442 910
rect 1252 79 1286 910
<< metal1 >>
rect -391 79 -331 859
rect -303 79 -243 859
rect -51 793 -45 853
rect 81 793 87 853
rect -51 765 87 793
rect 723 793 729 853
rect 855 793 861 853
rect 207 705 213 765
rect 339 705 345 765
rect 465 705 471 765
rect 597 705 603 765
rect 723 760 861 793
rect 117 227 177 233
rect 117 161 177 167
rect 633 227 693 233
rect 633 161 693 167
<< via1 >>
rect -45 793 81 853
rect 729 793 855 853
rect 213 705 339 765
rect 471 705 597 765
rect 117 167 177 227
rect 633 167 693 227
<< metal2 >>
rect -397 793 -45 853
rect 81 793 729 853
rect 855 793 892 853
rect -397 705 213 765
rect 339 705 471 765
rect 597 705 892 765
rect 111 167 117 227
rect 177 167 633 227
rect 693 167 699 227
use sky130_fd_pr__pfet_g5v0d10v5_V8EYZH  sky130_fd_pr__pfet_g5v0d10v5_V8EYZH_0
timestamp 1749911905
transform 1 0 405 0 1 415
box -611 -402 611 364
<< end >>
