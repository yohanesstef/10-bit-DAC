magic
tech sky130A
magscale 1 2
timestamp 1750201071
<< nwell >>
rect -5785 3966 -1204 6082
<< mvnsubdiff >>
rect -5719 6003 -1270 6016
rect -5719 5969 -5646 6003
rect -1343 5969 -1270 6003
rect -5719 5956 -1270 5969
rect -5719 5943 -5659 5956
rect -5719 4105 -5706 5943
rect -5672 4105 -5659 5943
rect -1330 5943 -1270 5956
rect -5719 4092 -5659 4105
rect -1330 4105 -1317 5943
rect -1283 4105 -1270 5943
rect -1330 4092 -1270 4105
rect -5719 4079 -1270 4092
rect -5719 4045 -5646 4079
rect -1343 4045 -1270 4079
rect -5719 4032 -1270 4045
<< mvnsubdiffcont >>
rect -5646 5969 -1343 6003
rect -5706 4105 -5672 5943
rect -1317 4105 -1283 5943
rect -5646 4045 -1343 4079
<< poly >>
rect -5648 5020 -5588 5028
rect -5515 5020 -1515 5028
rect -1442 5020 -1382 5028
<< viali >>
rect -5706 5969 -5646 6003
rect -5646 5969 -1343 6003
rect -1343 5969 -1283 6003
rect -5706 5943 -5672 5969
rect -5706 4105 -5672 5943
rect -5706 4079 -5672 4105
rect -1317 5943 -1283 5969
rect -1317 4105 -1283 5943
rect -1317 4079 -1283 4105
rect -5706 4045 -5646 4079
rect -5646 4045 -1343 4079
rect -1343 4045 -1283 4079
<< metal1 >>
rect -5729 6003 -1260 6026
rect -5729 4045 -5706 6003
rect -5672 5946 -1317 5969
rect -5672 4102 -5649 5946
rect -5567 5054 -5521 5542
rect -1509 5414 -1463 5542
rect -1509 4994 -1463 5054
rect -5567 4593 -5521 4634
rect -5567 4547 -5015 4593
rect -5567 4506 -5521 4547
rect -1510 4506 -1464 4634
rect -1340 4102 -1317 5946
rect -5672 4079 -1317 4102
rect -1283 4045 -1260 6003
rect -5729 4022 -1260 4045
use cm2_pcell3_cell  cm2_pcell3_cell_0
timestamp 1750201071
transform 1 0 -3823 0 -1 13345
box -1825 7377 2441 7903
use cm2_pcell3_cell  cm2_pcell3_cell_1
timestamp 1750201071
transform 1 0 -3823 0 1 -2389
box -1825 7377 2441 7903
use cm2_pcell3_cell  cm2_pcell3_cell_2
timestamp 1750201071
transform 1 0 -3823 0 -1 12437
box -1825 7377 2441 7903
use cm2_pcell3_cell  cm2_pcell3_cell_3
timestamp 1750201071
transform 1 0 -3823 0 1 -3297
box -1825 7377 2441 7903
<< end >>
