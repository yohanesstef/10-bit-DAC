magic
tech sky130A
magscale 1 2
timestamp 1749538868
<< metal1 >>
rect 16306 -23125 16366 -21181
rect 16394 -22477 16454 -21181
rect 16482 -21829 16542 -21181
rect 16570 -21443 16575 -21181
rect 16575 -21505 16991 -21443
rect 17575 -21505 17635 -21181
rect 17552 -21767 17635 -21505
rect 17131 -21829 17552 -21767
rect 16482 -22091 16570 -21829
rect 16482 -22110 16991 -22091
rect 16570 -22153 16991 -22110
rect 17663 -22153 17723 -21181
rect 17552 -22415 17723 -22153
rect 17136 -22477 17552 -22415
rect 16394 -22739 16565 -22477
rect 16570 -22801 16986 -22739
rect 17751 -22801 17811 -21181
rect 17552 -23063 17811 -22801
rect 17136 -23125 17552 -23063
rect 16306 -23387 16565 -23125
rect 16565 -23449 16981 -23387
use sky130_fd_pr__res_xhigh_po_1p41_6E4SWG  sky130_fd_pr__res_xhigh_po_1p41_6E4SWG_0
timestamp 1748944356
transform 0 -1 17061 1 0 -22608
box -141 -502 141 502
use sky130_fd_pr__res_xhigh_po_1p41_9JVM35  sky130_fd_pr__res_xhigh_po_1p41_9JVM35_0
timestamp 1748944356
transform 0 -1 17061 1 0 -23580
box -141 -507 141 507
use sky130_fd_pr__res_xhigh_po_1p41_9JVP35  sky130_fd_pr__res_xhigh_po_1p41_9JVP35_0
timestamp 1749123188
transform 0 -1 17061 1 0 -23904
box -141 -507 141 507
use sky130_fd_pr__res_xhigh_po_1p41_B5ZH9J  sky130_fd_pr__res_xhigh_po_1p41_B5ZH9J_0
timestamp 1749202939
transform 0 -1 17061 1 0 -20988
box -141 -492 141 492
use sky130_fd_pr__res_xhigh_po_1p41_6E4SWG  XR42
timestamp 1748944356
transform 0 -1 17061 1 0 -23256
box -141 -502 141 502
use sky130_fd_pr__res_xhigh_po_1p41_53UW4Z  XR43
timestamp 1748944356
transform 0 -1 17061 1 0 -22932
box -141 -497 141 497
use sky130_fd_pr__res_xhigh_po_1p41_53UW4Z  XR45
timestamp 1748944356
transform 0 -1 17061 1 0 -22284
box -141 -497 141 497
use sky130_fd_pr__res_xhigh_po_1p41_53UW4Z  XR46
timestamp 1748944356
transform 0 -1 17061 1 0 -21960
box -141 -497 141 497
use sky130_fd_pr__res_xhigh_po_1p41_53UW4Z  XR47
timestamp 1748944356
transform 0 -1 17061 1 0 -21636
box -141 -497 141 497
use sky130_fd_pr__res_xhigh_po_1p41_B5ZK9J  XR48
timestamp 1748944356
transform 0 -1 17061 1 0 -21312
box -141 -492 141 492
<< end >>
