magic
tech sky130A
magscale 1 2
timestamp 1751042016
<< error_s >>
rect 255 -18 323 -2
rect 239 -19 339 -18
rect 228 -46 350 -40
rect 205 -53 373 -52
<< nwell >>
rect -181 -164 719 1105
<< mvnsubdiff >>
rect -115 981 653 1039
rect -115 -40 -57 981
rect 595 -40 653 981
rect -115 -98 653 -40
<< locali >>
rect -103 993 641 1027
rect -103 -52 -69 993
rect 607 -52 641 993
rect -103 -86 641 -52
<< metal1 >>
rect 29 146 57 644
use sky130_fd_pr__pfet_g5v0d10v5_ZG42FA  sky130_fd_pr__pfet_g5v0d10v5_ZG42FA_0
timestamp 1750847642
transform 1 0 289 0 -1 317
box -174 -393 174 355
use sky130_fd_pr__pfet_g5v0d10v5_ZG42FA  sky130_fd_pr__pfet_g5v0d10v5_ZG42FA_1
timestamp 1750847642
transform 1 0 131 0 1 389
box -174 -393 174 355
<< end >>
