magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -658 307 658
<< psubdiff >>
rect -271 588 -175 622
rect 175 588 271 622
rect -271 526 -237 588
rect 237 526 271 588
rect -271 -588 -237 -526
rect 237 -588 271 -526
rect -271 -622 -175 -588
rect 175 -622 271 -588
<< psubdiffcont >>
rect -175 588 175 622
rect -271 -526 -237 526
rect 237 -526 271 526
rect -175 -622 175 -588
<< xpolycontact >>
rect -141 60 141 492
rect -141 -492 141 -60
<< xpolyres >>
rect -141 -60 141 60
<< locali >>
rect -271 588 -175 622
rect 175 588 271 622
rect -271 526 -237 588
rect 237 526 271 588
rect -271 -588 -237 -526
rect 237 -588 271 -526
rect -271 -622 -175 -588
rect 175 -622 271 -588
<< viali >>
rect -125 77 125 474
rect -125 -474 125 -77
<< metal1 >>
rect -131 474 131 486
rect -131 77 -125 474
rect 125 77 131 474
rect -131 65 131 77
rect -131 -77 131 -65
rect -131 -474 -125 -77
rect 125 -474 131 -77
rect -131 -486 131 -474
<< properties >>
string FIXED_BBOX -254 -605 254 605
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 0.759 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 1.343k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
