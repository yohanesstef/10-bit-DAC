magic
tech sky130A
magscale 1 2
timestamp 1749528210
<< error_s >>
rect 4591 2016 4597 2022
rect 4645 2016 4651 2022
rect 4585 2010 4591 2016
rect 4651 2010 4657 2016
rect 4585 1956 4591 1962
rect 4651 1956 4657 1962
rect 4591 1950 4597 1956
rect 4645 1950 4651 1956
rect 4315 1928 4321 1934
rect 4369 1928 4375 1934
rect 4309 1922 4315 1928
rect 4375 1922 4381 1928
rect 4309 1868 4315 1874
rect 4375 1868 4381 1874
rect 4315 1862 4321 1868
rect 4369 1862 4375 1868
rect 4039 1840 4045 1846
rect 4093 1840 4099 1846
rect 4033 1834 4039 1840
rect 4099 1834 4105 1840
rect 4033 1780 4039 1786
rect 4099 1780 4105 1786
rect 4039 1774 4045 1780
rect 4093 1774 4099 1780
rect 3763 1752 3769 1758
rect 3817 1752 3823 1758
rect 3757 1746 3763 1752
rect 3823 1746 3829 1752
rect 3757 1692 3763 1698
rect 3823 1692 3829 1698
rect 3763 1686 3769 1692
rect 3817 1686 3823 1692
rect 3487 1664 3493 1670
rect 3541 1664 3547 1670
rect 3481 1658 3487 1664
rect 3547 1658 3553 1664
rect 3481 1604 3487 1610
rect 3547 1604 3553 1610
rect 3487 1598 3493 1604
rect 3541 1598 3547 1604
rect 3211 1576 3217 1582
rect 3265 1576 3271 1582
rect 3205 1570 3211 1576
rect 3271 1570 3277 1576
rect 3205 1516 3211 1522
rect 3271 1516 3277 1522
rect 3211 1510 3217 1516
rect 3265 1510 3271 1516
rect 2935 1488 2941 1494
rect 2989 1488 2995 1494
rect 2929 1482 2935 1488
rect 2995 1482 3001 1488
rect 2929 1428 2935 1434
rect 2995 1428 3001 1434
rect 2935 1422 2941 1428
rect 2989 1422 2995 1428
rect 2659 1400 2665 1406
rect 2713 1400 2719 1406
rect 2653 1394 2659 1400
rect 2719 1394 2725 1400
rect 2653 1340 2659 1346
rect 2719 1340 2725 1346
rect 2659 1334 2665 1340
rect 2713 1334 2719 1340
rect 2437 1312 2443 1318
rect 2443 1306 2449 1312
rect 2443 1252 2449 1258
rect 2437 1246 2443 1252
<< nwell >>
rect 2208 736 5032 1344
<< mvnsubdiff >>
rect 2274 1266 4966 1278
rect 2274 1232 2382 1266
rect 4858 1232 4966 1266
rect 2274 1220 4966 1232
rect 2274 1170 2332 1220
rect 2274 910 2286 1170
rect 2320 910 2332 1170
rect 2274 860 2332 910
rect 4908 1170 4966 1220
rect 4908 910 4920 1170
rect 4954 910 4966 1170
rect 4908 860 4966 910
rect 2274 848 4966 860
rect 2274 814 2382 848
rect 4858 814 4966 848
rect 2274 802 4966 814
<< mvnsubdiffcont >>
rect 2382 1232 4858 1266
rect 2286 910 2320 1170
rect 4920 910 4954 1170
rect 2382 814 4858 848
<< locali >>
rect 2286 1232 2382 1266
rect 4858 1232 4954 1266
rect 2286 1170 2320 1232
rect 2286 848 2320 910
rect 4920 1170 4954 1232
rect 4920 848 4954 910
rect 2286 814 2382 848
rect 4858 814 4954 848
<< metal1 >>
rect 4591 2016 4651 2022
rect 4315 1928 4375 1934
rect 4039 1840 4099 1846
rect 3763 1752 3823 1758
rect 3487 1664 3547 1670
rect 3211 1576 3271 1582
rect 2935 1488 2995 1494
rect 2659 1400 2719 1406
rect 2383 1312 2443 1318
rect 2383 1161 2443 1252
rect 2659 1161 2719 1340
rect 2935 1161 2995 1428
rect 3211 1161 3271 1516
rect 3487 1161 3547 1604
rect 3763 1161 3823 1692
rect 4039 1161 4099 1780
rect 4315 1161 4375 1868
rect 4591 1161 4651 1956
rect 2383 1059 2442 1161
rect 2659 1059 2718 1161
rect 2935 1059 2994 1161
rect 3211 1059 3270 1161
rect 3487 1059 3546 1161
rect 3763 1059 3822 1161
rect 4039 1059 4098 1161
rect 4315 1059 4374 1161
rect 4591 1059 4650 1161
rect 2383 962 2443 1059
rect 2452 962 2453 1022
rect 2659 962 2719 1059
rect 2935 962 2995 1059
rect 3211 962 3271 1059
rect 3487 962 3547 1059
rect 3763 962 3823 1059
rect 4039 962 4099 1059
rect 4315 962 4375 1059
rect 4591 962 4651 1059
<< via1 >>
rect 4591 1956 4651 2016
rect 4315 1868 4375 1928
rect 4039 1780 4099 1840
rect 3763 1692 3823 1752
rect 3487 1604 3547 1664
rect 3211 1516 3271 1576
rect 2935 1428 2995 1488
rect 2659 1340 2719 1400
rect 2383 1252 2443 1312
<< metal2 >>
rect 2377 1252 2383 1312
use hpmos_1  hpmos_1_1
timestamp 1749230053
transform 1 0 2694 0 1 4117
box 1856 -3221 2204 -2971
use hpmos_4  hpmos_4_0
timestamp 1749384553
transform 1 0 1964 0 1 865
box 378 31 1554 281
use hpmos_4  hpmos_4_1
timestamp 1749384553
transform 1 0 3068 0 1 865
box 378 31 1554 281
<< end >>
