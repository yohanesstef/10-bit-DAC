magic
tech sky130A
magscale 1 2
timestamp 1750060026
<< mvnmos >>
rect -2000 -91 2000 29
<< mvndiff >>
rect -2058 17 -2000 29
rect -2058 -79 -2046 17
rect -2012 -79 -2000 17
rect -2058 -91 -2000 -79
rect 2000 17 2058 29
rect 2000 -79 2012 17
rect 2046 -79 2058 17
rect 2000 -91 2058 -79
<< mvndiffc >>
rect -2046 -79 -2012 17
rect 2012 -79 2046 17
<< poly >>
rect -2000 101 2000 117
rect -2000 67 -1984 101
rect 1984 67 2000 101
rect -2000 29 2000 67
rect -2000 -117 2000 -91
<< polycont >>
rect -1984 67 1984 101
<< locali >>
rect -2000 67 -1984 101
rect 1984 67 2000 101
rect -2046 17 -2012 33
rect -2046 -95 -2012 -79
rect 2012 17 2046 33
rect 2012 -95 2046 -79
<< viali >>
rect -1488 67 1488 101
rect -2046 -79 -2012 17
rect 2012 -79 2046 17
<< metal1 >>
rect -1500 101 1500 107
rect -1500 67 -1488 101
rect 1488 67 1500 101
rect -1500 61 1500 67
rect -2052 17 -2006 29
rect -2052 -79 -2046 17
rect -2012 -79 -2006 17
rect -2052 -91 -2006 -79
rect 2006 17 2052 29
rect 2006 -79 2012 17
rect 2046 -79 2052 17
rect 2006 -91 2052 -79
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.6 l 20 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
