magic
tech sky130A
magscale 1 2
timestamp 1749895928
<< error_s >>
rect -1475 2365 -1448 2375
rect -1501 2305 -1448 2365
rect -1475 2295 -1448 2305
rect -1447 2365 -1420 2375
rect 1534 2365 1561 2375
rect -1447 2305 -1394 2365
rect 1508 2305 1561 2365
rect -1447 2295 -1420 2305
rect 1534 2295 1561 2305
rect 1562 2365 1589 2375
rect 1562 2305 1615 2365
rect 1562 2295 1589 2305
rect -1475 2207 -1448 2267
rect -1447 2207 -1420 2267
rect 1534 2207 1561 2267
rect 1562 2207 1589 2267
rect -1475 1279 -1448 1339
rect -1447 1279 -1420 1339
rect 1534 1279 1561 1339
rect 1562 1279 1589 1339
rect -1475 1241 -1448 1251
rect -1501 1181 -1448 1241
rect -1475 1171 -1448 1181
rect -1447 1241 -1420 1251
rect 1534 1241 1561 1251
rect -1447 1181 -1394 1241
rect 1508 1181 1561 1241
rect -1447 1171 -1420 1181
rect 1534 1171 1561 1181
rect 1562 1241 1589 1251
rect 1562 1181 1615 1241
rect 1562 1171 1589 1181
rect -1475 1083 -1448 1143
rect -1447 1083 -1420 1143
rect 1534 1083 1561 1143
rect 1562 1083 1589 1143
rect -1475 155 -1448 215
rect -1447 155 -1420 215
rect 1534 155 1561 215
rect 1562 155 1589 215
rect -1475 117 -1448 127
rect -1501 57 -1448 117
rect -1475 47 -1448 57
rect -1447 117 -1420 127
rect 1534 117 1561 127
rect -1447 57 -1394 117
rect 1508 57 1561 117
rect -1447 47 -1420 57
rect 1534 47 1561 57
rect 1562 117 1589 127
rect 1562 57 1615 117
rect 1562 47 1589 57
use cm_pcell1_4_4  cm_pcell1_4_4_0
timestamp 1749895928
transform 1 0 -1035 0 1 591
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_1
timestamp 1749895928
transform 1 0 470 0 1 591
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_2
timestamp 1749895928
transform -1 0 -356 0 1 591
box 1026 -600 2672 1840
use cm_pcell1_4_4  cm_pcell1_4_4_3
timestamp 1749895928
transform -1 0 1149 0 1 591
box 1026 -600 2672 1840
<< end >>
