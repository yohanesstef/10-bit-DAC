magic
tech sky130A
magscale 1 2
timestamp 1743275510
<< pwell >>
rect -201 -654 201 654
<< psubdiff >>
rect -165 584 -69 618
rect 69 584 165 618
rect -165 522 -131 584
rect 131 522 165 584
rect -165 -584 -131 -522
rect 131 -584 165 -522
rect -165 -618 -69 -584
rect 69 -618 165 -584
<< psubdiffcont >>
rect -69 584 69 618
rect -165 -522 -131 522
rect 131 -522 165 522
rect -69 -618 69 -584
<< xpolycontact >>
rect -35 56 35 488
rect -35 -488 35 -56
<< xpolyres >>
rect -35 -56 35 56
<< locali >>
rect -165 584 -69 618
rect 69 584 165 618
rect -165 522 -131 584
rect 131 522 165 584
rect -165 -584 -131 -522
rect 131 -584 165 -522
rect -165 -618 -69 -584
rect 69 -618 165 -584
<< viali >>
rect -19 73 19 470
rect -19 -470 19 -73
<< metal1 >>
rect -25 470 25 482
rect -25 73 -19 470
rect 19 73 25 470
rect -25 61 25 73
rect -25 -73 25 -61
rect -25 -470 -19 -73
rect 19 -470 25 -73
rect -25 -482 25 -470
<< properties >>
string FIXED_BBOX -148 -601 148 601
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.718 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 5.178k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
