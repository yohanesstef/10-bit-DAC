magic
tech sky130A
magscale 1 2
timestamp 1749382758
<< metal1 >>
rect 1839 3483 1899 3489
rect 1751 3395 1811 3401
rect 1663 3219 1723 3225
rect 1575 3131 1635 3137
rect 1575 2955 1635 3071
rect 1663 2955 1723 3159
rect 1751 2955 1811 3335
rect 1839 2955 1899 3423
rect 2015 3131 2075 3659
rect 2103 3219 2163 3659
rect 2191 3307 2251 3659
rect 2279 3395 2339 3659
rect 2279 3329 2339 3335
rect 2191 3241 2251 3247
rect 2103 3153 2163 3159
rect 2367 3219 2427 3659
rect 2455 3483 2515 3659
rect 2455 3417 2515 3423
rect 2543 3395 2603 3659
rect 2543 3329 2603 3335
rect 2367 3153 2427 3159
rect 2015 3065 2075 3071
rect 2631 3043 2691 3659
rect 2279 2983 2691 3043
rect 2279 2955 2339 2983
<< via1 >>
rect 1839 3423 1899 3483
rect 1751 3335 1811 3395
rect 1663 3159 1723 3219
rect 1575 3071 1635 3131
rect 2279 3335 2339 3395
rect 2191 3247 2251 3307
rect 2103 3159 2163 3219
rect 2455 3423 2515 3483
rect 2543 3335 2603 3395
rect 2367 3159 2427 3219
rect 2015 3071 2075 3131
<< metal2 >>
rect 1833 3423 1839 3483
rect 1899 3423 2455 3483
rect 2515 3423 2521 3483
rect 1745 3335 1751 3395
rect 1811 3335 2279 3395
rect 2339 3335 2345 3395
rect 2537 3335 2543 3395
rect 2603 3335 2796 3395
rect 2185 3247 2191 3307
rect 2251 3247 2796 3307
rect 1657 3159 1663 3219
rect 1723 3159 2103 3219
rect 2163 3159 2169 3219
rect 2361 3159 2367 3219
rect 2427 3159 2796 3219
rect 1569 3071 1575 3131
rect 1635 3071 2015 3131
rect 2075 3071 2081 3131
<< end >>
