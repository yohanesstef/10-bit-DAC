magic
tech sky130A
magscale 1 2
timestamp 1750064013
<< error_p >>
rect -353 -578 -323 510
rect -287 -512 -257 444
rect 257 -512 287 444
rect -287 -516 287 -512
rect 323 -578 353 510
rect -353 -582 353 -578
<< nwell >>
rect -323 -578 323 544
<< mvpmos >>
rect -229 -516 -29 444
rect 29 -516 229 444
<< mvpdiff >>
rect -287 432 -229 444
rect -287 -504 -275 432
rect -241 -504 -229 432
rect -287 -516 -229 -504
rect -29 432 29 444
rect -29 -504 -17 432
rect 17 -504 29 432
rect -29 -516 29 -504
rect 229 432 287 444
rect 229 -504 241 432
rect 275 -504 287 432
rect 229 -516 287 -504
<< mvpdiffc >>
rect -275 -504 -241 432
rect -17 -504 17 432
rect 241 -504 275 432
<< poly >>
rect -229 525 -29 541
rect -229 491 -213 525
rect -45 491 -29 525
rect -229 444 -29 491
rect 29 525 229 541
rect 29 491 45 525
rect 213 491 229 525
rect 29 444 229 491
rect -229 -542 -29 -516
rect 29 -542 229 -516
<< polycont >>
rect -213 491 -45 525
rect 45 491 213 525
<< locali >>
rect -229 491 -213 525
rect -45 491 -29 525
rect 29 491 45 525
rect 213 491 229 525
rect -275 432 -241 448
rect -275 -520 -241 -504
rect -17 432 17 448
rect -17 -520 17 -504
rect 241 432 275 448
rect 241 -520 275 -504
<< viali >>
rect -192 491 -66 525
rect 66 491 192 525
rect -275 -504 -241 432
rect -17 -504 17 432
rect 241 -504 275 432
<< metal1 >>
rect -204 525 -54 531
rect -204 491 -192 525
rect -66 491 -54 525
rect -204 485 -54 491
rect 54 525 204 531
rect 54 491 66 525
rect 192 491 204 525
rect 54 485 204 491
rect -281 432 -235 444
rect -281 -504 -275 432
rect -241 -504 -235 432
rect -281 -516 -235 -504
rect -23 432 23 444
rect -23 -504 -17 432
rect 17 -504 23 432
rect -23 -516 23 -504
rect 235 432 281 444
rect 235 -504 241 432
rect 275 -504 281 432
rect 235 -516 281 -504
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.8 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
