magic
tech sky130A
magscale 1 2
timestamp 1750195772
<< error_s >>
rect 102 517 686 523
rect 48 463 740 469
<< pwell >>
rect 1985 1416 3621 1496
rect 1985 506 2065 1416
rect 3541 506 3621 1416
rect 1985 426 3621 506
<< mvpsubdiff >>
rect 1995 1426 3611 1486
rect 1995 496 2055 1426
rect 3551 496 3611 1426
rect 1995 436 3611 496
<< poly >>
rect 2181 982 2241 1216
rect 3365 982 3425 1216
rect 2181 706 2241 940
rect 3365 706 3425 940
<< locali >>
rect 2008 1439 3598 1473
rect 2008 483 2042 1439
rect 3564 483 3598 1439
rect 2008 449 3598 483
<< metal1 >>
rect 1985 1416 3621 1496
rect 1985 506 2065 1416
rect 3453 1382 3513 1388
rect 2391 1322 2397 1382
rect 2457 1322 2463 1382
rect 2093 1294 2153 1300
rect 2093 776 2153 1234
rect 2397 1206 2457 1322
rect 2358 1146 2364 1206
rect 2490 1146 2496 1206
rect 3110 1146 3116 1206
rect 3242 1146 3248 1206
rect 2093 710 2153 716
rect 2181 1008 2275 1128
rect 2526 1079 2586 1085
rect 3073 1019 3247 1079
rect 2526 1013 2586 1019
rect 2181 688 2241 1008
rect 2651 997 2697 1008
rect 2909 997 2955 1008
rect 2644 991 2704 997
rect 2644 925 2704 931
rect 2902 991 2962 997
rect 3101 980 3107 991
rect 2902 925 2962 931
rect 3027 940 3107 980
rect 2651 914 2697 925
rect 2909 914 2955 925
rect 3027 914 3073 940
rect 3101 931 3107 940
rect 3167 931 3173 991
rect 3201 909 3247 1019
rect 3331 1008 3425 1128
rect 2526 903 2586 909
rect 2526 837 2586 843
rect 3195 903 3255 909
rect 3195 837 3255 843
rect 2181 622 2241 628
rect 2275 606 2321 794
rect 2358 716 2364 776
rect 2490 716 2496 776
rect 3110 716 3116 776
rect 3242 716 3248 776
rect 3285 694 3331 795
rect 3277 688 3337 694
rect 3277 622 3337 628
rect 2268 600 2328 606
rect 2268 534 2328 540
rect 3365 600 3425 1008
rect 3453 776 3513 1322
rect 3453 710 3513 716
rect 3365 534 3425 540
rect 3541 506 3621 1416
rect 1985 426 3621 506
<< via1 >>
rect 2397 1322 2457 1382
rect 3453 1322 3513 1382
rect 2093 1234 2153 1294
rect 2364 1146 2490 1206
rect 3116 1146 3242 1206
rect 2093 716 2153 776
rect 2526 1019 2586 1079
rect 2644 931 2704 991
rect 2902 931 2962 991
rect 3107 931 3167 991
rect 2526 843 2586 903
rect 3195 843 3255 903
rect 2181 628 2241 688
rect 2364 716 2490 776
rect 3116 716 3242 776
rect 3277 628 3337 688
rect 2268 540 2328 600
rect 3453 716 3513 776
rect 3365 540 3425 600
<< metal2 >>
rect 2391 1322 2397 1382
rect 2457 1322 3453 1382
rect 3513 1322 3519 1382
rect 2087 1234 2093 1294
rect 2153 1234 3248 1294
rect 3110 1206 3248 1234
rect 2358 1146 2364 1206
rect 2490 1146 2496 1206
rect 3110 1146 3116 1206
rect 3242 1146 3248 1206
rect 2520 1019 2526 1079
rect 2586 1019 3167 1079
rect 3107 991 3167 1019
rect 2638 931 2644 991
rect 2704 931 2710 991
rect 2896 931 2902 991
rect 2962 931 2968 991
rect 3101 931 3107 991
rect 3167 931 3173 991
rect 2520 843 2526 903
rect 2586 843 3195 903
rect 3255 843 3261 903
rect 2087 716 2093 776
rect 2153 716 2364 776
rect 2490 716 2496 776
rect 3110 716 3116 776
rect 3242 716 3453 776
rect 3513 716 3519 776
rect 2175 628 2181 688
rect 2241 628 3277 688
rect 3337 628 3344 688
rect 2262 540 2268 600
rect 2328 540 3365 600
rect 3425 540 3431 600
use sky130_fd_pr__nfet_g5v0d10v5_EZHYDL  sky130_fd_pr__nfet_g5v0d10v5_EZHYDL_0
timestamp 1750195294
transform 1 0 370 0 1 218
box -457 -287 457 287
use sky130_fd_pr__nfet_g5v0d10v5_QKV39N  sky130_fd_pr__nfet_g5v0d10v5_QKV39N_0 ~/10-bit-DAC/mag
timestamp 1750058993
transform 1 0 2427 0 1 1099
box -158 -117 158 117
use sky130_fd_pr__nfet_g5v0d10v5_QKV39N  sky130_fd_pr__nfet_g5v0d10v5_QKV39N_1
timestamp 1750058993
transform 1 0 2803 0 1 1099
box -158 -117 158 117
use sky130_fd_pr__nfet_g5v0d10v5_QKV39N  sky130_fd_pr__nfet_g5v0d10v5_QKV39N_2
timestamp 1750058993
transform 1 0 3179 0 1 1099
box -158 -117 158 117
use sky130_fd_pr__nfet_g5v0d10v5_QKV39N  sky130_fd_pr__nfet_g5v0d10v5_QKV39N_3
timestamp 1750058993
transform 1 0 2427 0 -1 823
box -158 -117 158 117
use sky130_fd_pr__nfet_g5v0d10v5_QKV39N  sky130_fd_pr__nfet_g5v0d10v5_QKV39N_4
timestamp 1750058993
transform 1 0 2803 0 -1 823
box -158 -117 158 117
use sky130_fd_pr__nfet_g5v0d10v5_QKV39N  sky130_fd_pr__nfet_g5v0d10v5_QKV39N_5
timestamp 1750058993
transform 1 0 3179 0 -1 823
box -158 -117 158 117
use sky130_fd_pr__nfet_g5v0d10v5_ZUMGVX  sky130_fd_pr__nfet_g5v0d10v5_ZUMGVX_0
timestamp 1750195294
transform 1 0 394 0 1 1238
box -328 -757 328 757
<< end >>
