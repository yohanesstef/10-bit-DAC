magic
tech sky130A
magscale 1 2
timestamp 1749714889
<< magnet >>
rect -7 1616 7 1630
rect 511 1616 525 1630
rect 539 1616 553 1630
rect 1057 1616 1071 1630
rect 1085 1616 1099 1630
rect 1603 1616 1617 1630
rect 1631 1616 1645 1630
rect 2149 1616 2163 1630
rect -21 1602 21 1616
rect -7 1588 21 1602
rect 49 1588 77 1616
rect 105 1588 133 1616
rect 161 1588 189 1616
rect 217 1588 245 1616
rect 273 1588 301 1616
rect 329 1588 357 1616
rect 385 1588 413 1616
rect 441 1588 469 1616
rect 497 1602 567 1616
rect 497 1588 525 1602
rect 539 1588 567 1602
rect 595 1588 623 1616
rect 651 1588 679 1616
rect 707 1588 735 1616
rect 763 1588 791 1616
rect 819 1588 847 1616
rect 875 1588 903 1616
rect 931 1588 959 1616
rect 987 1588 1015 1616
rect 1043 1602 1113 1616
rect 1043 1588 1071 1602
rect 1085 1588 1113 1602
rect 1141 1588 1169 1616
rect 1197 1588 1225 1616
rect 1253 1588 1281 1616
rect 1309 1588 1337 1616
rect 1365 1588 1393 1616
rect 1421 1588 1449 1616
rect 1477 1588 1505 1616
rect 1533 1588 1561 1616
rect 1589 1602 1659 1616
rect 1589 1588 1617 1602
rect 1631 1588 1659 1602
rect 1687 1588 1715 1616
rect 1743 1588 1771 1616
rect 1799 1588 1827 1616
rect 1855 1588 1883 1616
rect 1911 1588 1939 1616
rect 1967 1588 1995 1616
rect 2023 1588 2051 1616
rect 2079 1588 2107 1616
rect 2135 1602 2177 1616
rect 2135 1588 2163 1602
rect -7 1532 21 1560
rect 49 1532 77 1560
rect 105 1532 133 1560
rect 161 1532 189 1560
rect 217 1532 245 1560
rect 273 1532 301 1560
rect 329 1532 357 1560
rect 385 1532 413 1560
rect 441 1532 469 1560
rect 497 1532 525 1560
rect 539 1532 567 1560
rect 595 1532 623 1560
rect 651 1532 679 1560
rect 707 1532 735 1560
rect 763 1532 791 1560
rect 819 1532 847 1560
rect 875 1532 903 1560
rect 931 1532 959 1560
rect 987 1532 1015 1560
rect 1043 1532 1071 1560
rect 1085 1532 1113 1560
rect 1141 1532 1169 1560
rect 1197 1532 1225 1560
rect 1253 1532 1281 1560
rect 1309 1532 1337 1560
rect 1365 1532 1393 1560
rect 1421 1532 1449 1560
rect 1477 1532 1505 1560
rect 1533 1532 1561 1560
rect 1589 1532 1617 1560
rect 1631 1532 1659 1560
rect 1687 1532 1715 1560
rect 1743 1532 1771 1560
rect 1799 1532 1827 1560
rect 1855 1532 1883 1560
rect 1911 1532 1939 1560
rect 1967 1532 1995 1560
rect 2023 1532 2051 1560
rect 2079 1532 2107 1560
rect 2135 1532 2163 1560
rect -7 1476 21 1504
rect 49 1476 77 1504
rect 105 1476 133 1504
rect 161 1476 189 1504
rect 217 1476 245 1504
rect 273 1476 301 1504
rect 329 1476 357 1504
rect 385 1476 413 1504
rect 441 1476 469 1504
rect 497 1476 525 1504
rect 539 1476 567 1504
rect 595 1476 623 1504
rect 651 1476 679 1504
rect 707 1476 735 1504
rect 763 1476 791 1504
rect 819 1476 847 1504
rect 875 1476 903 1504
rect 931 1476 959 1504
rect 987 1476 1015 1504
rect 1043 1476 1071 1504
rect 1085 1476 1113 1504
rect 1141 1476 1169 1504
rect 1197 1476 1225 1504
rect 1253 1476 1281 1504
rect 1309 1476 1337 1504
rect 1365 1476 1393 1504
rect 1421 1476 1449 1504
rect 1477 1476 1505 1504
rect 1533 1476 1561 1504
rect 1589 1476 1617 1504
rect 1631 1476 1659 1504
rect 1687 1476 1715 1504
rect 1743 1476 1771 1504
rect 1799 1476 1827 1504
rect 1855 1476 1883 1504
rect 1911 1476 1939 1504
rect 1967 1476 1995 1504
rect 2023 1476 2051 1504
rect 2079 1476 2107 1504
rect 2135 1476 2163 1504
rect -7 1420 21 1448
rect 49 1420 77 1448
rect 105 1420 133 1448
rect 161 1420 189 1448
rect 217 1420 245 1448
rect 273 1420 301 1448
rect 329 1420 357 1448
rect 385 1420 413 1448
rect 441 1420 469 1448
rect 497 1420 525 1448
rect 539 1420 567 1448
rect 595 1420 623 1448
rect 651 1420 679 1448
rect 707 1420 735 1448
rect 763 1420 791 1448
rect 819 1420 847 1448
rect 875 1420 903 1448
rect 931 1420 959 1448
rect 987 1420 1015 1448
rect 1043 1420 1071 1448
rect 1085 1420 1113 1448
rect 1141 1420 1169 1448
rect 1197 1420 1225 1448
rect 1253 1420 1281 1448
rect 1309 1420 1337 1448
rect 1365 1420 1393 1448
rect 1421 1420 1449 1448
rect 1477 1420 1505 1448
rect 1533 1420 1561 1448
rect 1589 1420 1617 1448
rect 1631 1420 1659 1448
rect 1687 1420 1715 1448
rect 1743 1420 1771 1448
rect 1799 1420 1827 1448
rect 1855 1420 1883 1448
rect 1911 1420 1939 1448
rect 1967 1420 1995 1448
rect 2023 1420 2051 1448
rect 2079 1420 2107 1448
rect 2135 1420 2163 1448
rect -7 1364 21 1392
rect 49 1364 77 1392
rect 105 1364 133 1392
rect 161 1364 189 1392
rect 217 1364 245 1392
rect 273 1364 301 1392
rect 329 1364 357 1392
rect 385 1364 413 1392
rect 441 1364 469 1392
rect 497 1364 525 1392
rect 539 1364 567 1392
rect 595 1364 623 1392
rect 651 1364 679 1392
rect 707 1364 735 1392
rect 763 1364 791 1392
rect 819 1364 847 1392
rect 875 1364 903 1392
rect 931 1364 959 1392
rect 987 1364 1015 1392
rect 1043 1364 1071 1392
rect 1085 1364 1113 1392
rect 1141 1364 1169 1392
rect 1197 1364 1225 1392
rect 1253 1364 1281 1392
rect 1309 1364 1337 1392
rect 1365 1364 1393 1392
rect 1421 1364 1449 1392
rect 1477 1364 1505 1392
rect 1533 1364 1561 1392
rect 1589 1364 1617 1392
rect 1631 1364 1659 1392
rect 1687 1364 1715 1392
rect 1743 1364 1771 1392
rect 1799 1364 1827 1392
rect 1855 1364 1883 1392
rect 1911 1364 1939 1392
rect 1967 1364 1995 1392
rect 2023 1364 2051 1392
rect 2079 1364 2107 1392
rect 2135 1364 2163 1392
rect -7 1308 21 1336
rect 49 1308 77 1336
rect 105 1308 133 1336
rect 161 1308 189 1336
rect 217 1308 245 1336
rect 273 1308 301 1336
rect 329 1308 357 1336
rect 385 1308 413 1336
rect 441 1308 469 1336
rect 497 1308 525 1336
rect 539 1308 567 1336
rect 595 1308 623 1336
rect 651 1308 679 1336
rect 707 1308 735 1336
rect 763 1308 791 1336
rect 819 1308 847 1336
rect 875 1308 903 1336
rect 931 1308 959 1336
rect 987 1308 1015 1336
rect 1043 1308 1071 1336
rect 1085 1308 1113 1336
rect 1141 1308 1169 1336
rect 1197 1308 1225 1336
rect 1253 1308 1281 1336
rect 1309 1308 1337 1336
rect 1365 1308 1393 1336
rect 1421 1308 1449 1336
rect 1477 1308 1505 1336
rect 1533 1308 1561 1336
rect 1589 1308 1617 1336
rect 1631 1308 1659 1336
rect 1687 1308 1715 1336
rect 1743 1308 1771 1336
rect 1799 1308 1827 1336
rect 1855 1308 1883 1336
rect 1911 1308 1939 1336
rect 1967 1308 1995 1336
rect 2023 1308 2051 1336
rect 2079 1308 2107 1336
rect 2135 1308 2163 1336
rect -7 1252 21 1280
rect 49 1252 77 1280
rect 105 1252 133 1280
rect 161 1252 189 1280
rect 217 1252 245 1280
rect 273 1252 301 1280
rect 329 1252 357 1280
rect 385 1252 413 1280
rect 441 1252 469 1280
rect 497 1252 525 1280
rect 539 1252 567 1280
rect 595 1252 623 1280
rect 651 1252 679 1280
rect 707 1252 735 1280
rect 763 1252 791 1280
rect 819 1252 847 1280
rect 875 1252 903 1280
rect 931 1252 959 1280
rect 987 1252 1015 1280
rect 1043 1252 1071 1280
rect 1085 1252 1113 1280
rect 1141 1252 1169 1280
rect 1197 1252 1225 1280
rect 1253 1252 1281 1280
rect 1309 1252 1337 1280
rect 1365 1252 1393 1280
rect 1421 1252 1449 1280
rect 1477 1252 1505 1280
rect 1533 1252 1561 1280
rect 1589 1252 1617 1280
rect 1631 1252 1659 1280
rect 1687 1252 1715 1280
rect 1743 1252 1771 1280
rect 1799 1252 1827 1280
rect 1855 1252 1883 1280
rect 1911 1252 1939 1280
rect 1967 1252 1995 1280
rect 2023 1252 2051 1280
rect 2079 1252 2107 1280
rect 2135 1252 2163 1280
rect -7 1196 21 1224
rect 49 1196 77 1224
rect 105 1196 133 1224
rect 161 1196 189 1224
rect 217 1196 245 1224
rect 273 1196 301 1224
rect 329 1196 357 1224
rect 385 1196 413 1224
rect 441 1196 469 1224
rect 497 1196 525 1224
rect 539 1196 567 1224
rect 595 1196 623 1224
rect 651 1196 679 1224
rect 707 1196 735 1224
rect 763 1196 791 1224
rect 819 1196 847 1224
rect 875 1196 903 1224
rect 931 1196 959 1224
rect 987 1196 1015 1224
rect 1043 1196 1071 1224
rect 1085 1196 1113 1224
rect 1141 1196 1169 1224
rect 1197 1196 1225 1224
rect 1253 1196 1281 1224
rect 1309 1196 1337 1224
rect 1365 1196 1393 1224
rect 1421 1196 1449 1224
rect 1477 1196 1505 1224
rect 1533 1196 1561 1224
rect 1589 1196 1617 1224
rect 1631 1196 1659 1224
rect 1687 1196 1715 1224
rect 1743 1196 1771 1224
rect 1799 1196 1827 1224
rect 1855 1196 1883 1224
rect 1911 1196 1939 1224
rect 1967 1196 1995 1224
rect 2023 1196 2051 1224
rect 2079 1196 2107 1224
rect 2135 1196 2163 1224
rect -7 1140 21 1168
rect 49 1140 77 1168
rect 105 1140 133 1168
rect 161 1140 189 1168
rect 217 1140 245 1168
rect 273 1140 301 1168
rect 329 1140 357 1168
rect 385 1140 413 1168
rect 441 1140 469 1168
rect 497 1140 525 1168
rect 539 1140 567 1168
rect 595 1140 623 1168
rect 651 1140 679 1168
rect 707 1140 735 1168
rect 763 1140 791 1168
rect 819 1140 847 1168
rect 875 1140 903 1168
rect 931 1140 959 1168
rect 987 1140 1015 1168
rect 1043 1140 1071 1168
rect 1085 1140 1113 1168
rect 1141 1140 1169 1168
rect 1197 1140 1225 1168
rect 1253 1140 1281 1168
rect 1309 1140 1337 1168
rect 1365 1140 1393 1168
rect 1421 1140 1449 1168
rect 1477 1140 1505 1168
rect 1533 1140 1561 1168
rect 1589 1140 1617 1168
rect 1631 1140 1659 1168
rect 1687 1140 1715 1168
rect 1743 1140 1771 1168
rect 1799 1140 1827 1168
rect 1855 1140 1883 1168
rect 1911 1140 1939 1168
rect 1967 1140 1995 1168
rect 2023 1140 2051 1168
rect 2079 1140 2107 1168
rect 2135 1140 2163 1168
rect -7 1098 21 1112
rect -21 1084 21 1098
rect 49 1084 77 1112
rect 105 1084 133 1112
rect 161 1084 189 1112
rect 217 1084 245 1112
rect 273 1084 301 1112
rect 329 1084 357 1112
rect 385 1084 413 1112
rect 441 1084 469 1112
rect 497 1098 525 1112
rect 539 1098 567 1112
rect 497 1084 567 1098
rect 595 1084 623 1112
rect 651 1084 679 1112
rect 707 1084 735 1112
rect 763 1084 791 1112
rect 819 1084 847 1112
rect 875 1084 903 1112
rect 931 1084 959 1112
rect 987 1084 1015 1112
rect 1043 1098 1071 1112
rect 1085 1098 1113 1112
rect 1043 1084 1113 1098
rect 1141 1084 1169 1112
rect 1197 1084 1225 1112
rect 1253 1084 1281 1112
rect 1309 1084 1337 1112
rect 1365 1084 1393 1112
rect 1421 1084 1449 1112
rect 1477 1084 1505 1112
rect 1533 1084 1561 1112
rect 1589 1098 1617 1112
rect 1631 1098 1659 1112
rect 1589 1084 1659 1098
rect 1687 1084 1715 1112
rect 1743 1084 1771 1112
rect 1799 1084 1827 1112
rect 1855 1084 1883 1112
rect 1911 1084 1939 1112
rect 1967 1084 1995 1112
rect 2023 1084 2051 1112
rect 2079 1084 2107 1112
rect 2135 1098 2163 1112
rect 2135 1084 2177 1098
rect -7 1070 7 1084
rect 511 1070 525 1084
rect 539 1070 553 1084
rect 1057 1070 1071 1084
rect 1085 1070 1099 1084
rect 1603 1070 1617 1084
rect 1631 1070 1645 1084
rect 2149 1070 2163 1084
rect -21 1056 21 1070
rect -7 1042 21 1056
rect 49 1042 77 1070
rect 105 1042 133 1070
rect 161 1042 189 1070
rect 217 1042 245 1070
rect 273 1042 301 1070
rect 329 1042 357 1070
rect 385 1042 413 1070
rect 441 1042 469 1070
rect 497 1056 567 1070
rect 497 1042 525 1056
rect 539 1042 567 1056
rect 595 1042 623 1070
rect 651 1042 679 1070
rect 707 1042 735 1070
rect 763 1042 791 1070
rect 819 1042 847 1070
rect 875 1042 903 1070
rect 931 1042 959 1070
rect 987 1042 1015 1070
rect 1043 1056 1113 1070
rect 1043 1042 1071 1056
rect 1085 1042 1113 1056
rect 1141 1042 1169 1070
rect 1197 1042 1225 1070
rect 1253 1042 1281 1070
rect 1309 1042 1337 1070
rect 1365 1042 1393 1070
rect 1421 1042 1449 1070
rect 1477 1042 1505 1070
rect 1533 1042 1561 1070
rect 1589 1056 1659 1070
rect 1589 1042 1617 1056
rect 1631 1042 1659 1056
rect 1687 1042 1715 1070
rect 1743 1042 1771 1070
rect 1799 1042 1827 1070
rect 1855 1042 1883 1070
rect 1911 1042 1939 1070
rect 1967 1042 1995 1070
rect 2023 1042 2051 1070
rect 2079 1042 2107 1070
rect 2135 1056 2177 1070
rect 2135 1042 2163 1056
rect -7 986 21 1014
rect 49 986 77 1014
rect 105 986 133 1014
rect 161 986 189 1014
rect 217 986 245 1014
rect 273 986 301 1014
rect 329 986 357 1014
rect 385 986 413 1014
rect 441 986 469 1014
rect 497 986 525 1014
rect 539 986 567 1014
rect 595 986 623 1014
rect 651 986 679 1014
rect 707 986 735 1014
rect 763 986 791 1014
rect 819 986 847 1014
rect 875 986 903 1014
rect 931 986 959 1014
rect 987 986 1015 1014
rect 1043 986 1071 1014
rect 1085 986 1113 1014
rect 1141 986 1169 1014
rect 1197 986 1225 1014
rect 1253 986 1281 1014
rect 1309 986 1337 1014
rect 1365 986 1393 1014
rect 1421 986 1449 1014
rect 1477 986 1505 1014
rect 1533 986 1561 1014
rect 1589 986 1617 1014
rect 1631 986 1659 1014
rect 1687 986 1715 1014
rect 1743 986 1771 1014
rect 1799 986 1827 1014
rect 1855 986 1883 1014
rect 1911 986 1939 1014
rect 1967 986 1995 1014
rect 2023 986 2051 1014
rect 2079 986 2107 1014
rect 2135 986 2163 1014
rect -7 930 21 958
rect 49 930 77 958
rect 105 930 133 958
rect 161 930 189 958
rect 217 930 245 958
rect 273 930 301 958
rect 329 930 357 958
rect 385 930 413 958
rect 441 930 469 958
rect 497 930 525 958
rect 539 930 567 958
rect 595 930 623 958
rect 651 930 679 958
rect 707 930 735 958
rect 763 930 791 958
rect 819 930 847 958
rect 875 930 903 958
rect 931 930 959 958
rect 987 930 1015 958
rect 1043 930 1071 958
rect 1085 930 1113 958
rect 1141 930 1169 958
rect 1197 930 1225 958
rect 1253 930 1281 958
rect 1309 930 1337 958
rect 1365 930 1393 958
rect 1421 930 1449 958
rect 1477 930 1505 958
rect 1533 930 1561 958
rect 1589 930 1617 958
rect 1631 930 1659 958
rect 1687 930 1715 958
rect 1743 930 1771 958
rect 1799 930 1827 958
rect 1855 930 1883 958
rect 1911 930 1939 958
rect 1967 930 1995 958
rect 2023 930 2051 958
rect 2079 930 2107 958
rect 2135 930 2163 958
rect -7 874 21 902
rect 49 874 77 902
rect 105 874 133 902
rect 161 874 189 902
rect 217 874 245 902
rect 273 874 301 902
rect 329 874 357 902
rect 385 874 413 902
rect 441 874 469 902
rect 497 874 525 902
rect 539 874 567 902
rect 595 874 623 902
rect 651 874 679 902
rect 707 874 735 902
rect 763 874 791 902
rect 819 874 847 902
rect 875 874 903 902
rect 931 874 959 902
rect 987 874 1015 902
rect 1043 874 1071 902
rect 1085 874 1113 902
rect 1141 874 1169 902
rect 1197 874 1225 902
rect 1253 874 1281 902
rect 1309 874 1337 902
rect 1365 874 1393 902
rect 1421 874 1449 902
rect 1477 874 1505 902
rect 1533 874 1561 902
rect 1589 874 1617 902
rect 1631 874 1659 902
rect 1687 874 1715 902
rect 1743 874 1771 902
rect 1799 874 1827 902
rect 1855 874 1883 902
rect 1911 874 1939 902
rect 1967 874 1995 902
rect 2023 874 2051 902
rect 2079 874 2107 902
rect 2135 874 2163 902
rect -7 818 21 846
rect 49 818 77 846
rect 105 818 133 846
rect 161 818 189 846
rect 217 818 245 846
rect 273 818 301 846
rect 329 818 357 846
rect 385 818 413 846
rect 441 818 469 846
rect 497 818 525 846
rect 539 818 567 846
rect 595 818 623 846
rect 651 818 679 846
rect 707 818 735 846
rect 763 818 791 846
rect 819 818 847 846
rect 875 818 903 846
rect 931 818 959 846
rect 987 818 1015 846
rect 1043 818 1071 846
rect 1085 818 1113 846
rect 1141 818 1169 846
rect 1197 818 1225 846
rect 1253 818 1281 846
rect 1309 818 1337 846
rect 1365 818 1393 846
rect 1421 818 1449 846
rect 1477 818 1505 846
rect 1533 818 1561 846
rect 1589 818 1617 846
rect 1631 818 1659 846
rect 1687 818 1715 846
rect 1743 818 1771 846
rect 1799 818 1827 846
rect 1855 818 1883 846
rect 1911 818 1939 846
rect 1967 818 1995 846
rect 2023 818 2051 846
rect 2079 818 2107 846
rect 2135 818 2163 846
rect -7 762 21 790
rect 49 762 77 790
rect 105 762 133 790
rect 161 762 189 790
rect 217 762 245 790
rect 273 762 301 790
rect 329 762 357 790
rect 385 762 413 790
rect 441 762 469 790
rect 497 762 525 790
rect 539 762 567 790
rect 595 762 623 790
rect 651 762 679 790
rect 707 762 735 790
rect 763 762 791 790
rect 819 762 847 790
rect 875 762 903 790
rect 931 762 959 790
rect 987 762 1015 790
rect 1043 762 1071 790
rect 1085 762 1113 790
rect 1141 762 1169 790
rect 1197 762 1225 790
rect 1253 762 1281 790
rect 1309 762 1337 790
rect 1365 762 1393 790
rect 1421 762 1449 790
rect 1477 762 1505 790
rect 1533 762 1561 790
rect 1589 762 1617 790
rect 1631 762 1659 790
rect 1687 762 1715 790
rect 1743 762 1771 790
rect 1799 762 1827 790
rect 1855 762 1883 790
rect 1911 762 1939 790
rect 1967 762 1995 790
rect 2023 762 2051 790
rect 2079 762 2107 790
rect 2135 762 2163 790
rect -7 706 21 734
rect 49 706 77 734
rect 105 706 133 734
rect 161 706 189 734
rect 217 706 245 734
rect 273 706 301 734
rect 329 706 357 734
rect 385 706 413 734
rect 441 706 469 734
rect 497 706 525 734
rect 539 706 567 734
rect 595 706 623 734
rect 651 706 679 734
rect 707 706 735 734
rect 763 706 791 734
rect 819 706 847 734
rect 875 706 903 734
rect 931 706 959 734
rect 987 706 1015 734
rect 1043 706 1071 734
rect 1085 706 1113 734
rect 1141 706 1169 734
rect 1197 706 1225 734
rect 1253 706 1281 734
rect 1309 706 1337 734
rect 1365 706 1393 734
rect 1421 706 1449 734
rect 1477 706 1505 734
rect 1533 706 1561 734
rect 1589 706 1617 734
rect 1631 706 1659 734
rect 1687 706 1715 734
rect 1743 706 1771 734
rect 1799 706 1827 734
rect 1855 706 1883 734
rect 1911 706 1939 734
rect 1967 706 1995 734
rect 2023 706 2051 734
rect 2079 706 2107 734
rect 2135 706 2163 734
rect -7 650 21 678
rect 49 650 77 678
rect 105 650 133 678
rect 161 650 189 678
rect 217 650 245 678
rect 273 650 301 678
rect 329 650 357 678
rect 385 650 413 678
rect 441 650 469 678
rect 497 650 525 678
rect 539 650 567 678
rect 595 650 623 678
rect 651 650 679 678
rect 707 650 735 678
rect 763 650 791 678
rect 819 650 847 678
rect 875 650 903 678
rect 931 650 959 678
rect 987 650 1015 678
rect 1043 650 1071 678
rect 1085 650 1113 678
rect 1141 650 1169 678
rect 1197 650 1225 678
rect 1253 650 1281 678
rect 1309 650 1337 678
rect 1365 650 1393 678
rect 1421 650 1449 678
rect 1477 650 1505 678
rect 1533 650 1561 678
rect 1589 650 1617 678
rect 1631 650 1659 678
rect 1687 650 1715 678
rect 1743 650 1771 678
rect 1799 650 1827 678
rect 1855 650 1883 678
rect 1911 650 1939 678
rect 1967 650 1995 678
rect 2023 650 2051 678
rect 2079 650 2107 678
rect 2135 650 2163 678
rect -7 594 21 622
rect 49 594 77 622
rect 105 594 133 622
rect 161 594 189 622
rect 217 594 245 622
rect 273 594 301 622
rect 329 594 357 622
rect 385 594 413 622
rect 441 594 469 622
rect 497 594 525 622
rect 539 594 567 622
rect 595 594 623 622
rect 651 594 679 622
rect 707 594 735 622
rect 763 594 791 622
rect 819 594 847 622
rect 875 594 903 622
rect 931 594 959 622
rect 987 594 1015 622
rect 1043 594 1071 622
rect 1085 594 1113 622
rect 1141 594 1169 622
rect 1197 594 1225 622
rect 1253 594 1281 622
rect 1309 594 1337 622
rect 1365 594 1393 622
rect 1421 594 1449 622
rect 1477 594 1505 622
rect 1533 594 1561 622
rect 1589 594 1617 622
rect 1631 594 1659 622
rect 1687 594 1715 622
rect 1743 594 1771 622
rect 1799 594 1827 622
rect 1855 594 1883 622
rect 1911 594 1939 622
rect 1967 594 1995 622
rect 2023 594 2051 622
rect 2079 594 2107 622
rect 2135 594 2163 622
rect -7 552 21 566
rect -21 538 21 552
rect 49 538 77 566
rect 105 538 133 566
rect 161 538 189 566
rect 217 538 245 566
rect 273 538 301 566
rect 329 538 357 566
rect 385 538 413 566
rect 441 538 469 566
rect 497 552 525 566
rect 539 552 567 566
rect 497 538 567 552
rect 595 538 623 566
rect 651 538 679 566
rect 707 538 735 566
rect 763 538 791 566
rect 819 538 847 566
rect 875 538 903 566
rect 931 538 959 566
rect 987 538 1015 566
rect 1043 552 1071 566
rect 1085 552 1113 566
rect 1043 538 1113 552
rect 1141 538 1169 566
rect 1197 538 1225 566
rect 1253 538 1281 566
rect 1309 538 1337 566
rect 1365 538 1393 566
rect 1421 538 1449 566
rect 1477 538 1505 566
rect 1533 538 1561 566
rect 1589 552 1617 566
rect 1631 552 1659 566
rect 1589 538 1659 552
rect 1687 538 1715 566
rect 1743 538 1771 566
rect 1799 538 1827 566
rect 1855 538 1883 566
rect 1911 538 1939 566
rect 1967 538 1995 566
rect 2023 538 2051 566
rect 2079 538 2107 566
rect 2135 552 2163 566
rect 2135 538 2177 552
rect -7 524 7 538
rect 511 524 525 538
rect 539 524 553 538
rect 1057 524 1071 538
rect 1085 524 1099 538
rect 1603 524 1617 538
rect 1631 524 1645 538
rect 2149 524 2163 538
rect -21 510 21 524
rect -7 496 21 510
rect 49 496 77 524
rect 105 496 133 524
rect 161 496 189 524
rect 217 496 245 524
rect 273 496 301 524
rect 329 496 357 524
rect 385 496 413 524
rect 441 496 469 524
rect 497 510 567 524
rect 497 496 525 510
rect 539 496 567 510
rect 595 496 623 524
rect 651 496 679 524
rect 707 496 735 524
rect 763 496 791 524
rect 819 496 847 524
rect 875 496 903 524
rect 931 496 959 524
rect 987 496 1015 524
rect 1043 510 1113 524
rect 1043 496 1071 510
rect 1085 496 1113 510
rect 1141 496 1169 524
rect 1197 496 1225 524
rect 1253 496 1281 524
rect 1309 496 1337 524
rect 1365 496 1393 524
rect 1421 496 1449 524
rect 1477 496 1505 524
rect 1533 496 1561 524
rect 1589 510 1659 524
rect 1589 496 1617 510
rect 1631 496 1659 510
rect 1687 496 1715 524
rect 1743 496 1771 524
rect 1799 496 1827 524
rect 1855 496 1883 524
rect 1911 496 1939 524
rect 1967 496 1995 524
rect 2023 496 2051 524
rect 2079 496 2107 524
rect 2135 510 2177 524
rect 2135 496 2163 510
rect -7 440 21 468
rect 49 440 77 468
rect 105 440 133 468
rect 161 440 189 468
rect 217 440 245 468
rect 273 440 301 468
rect 329 440 357 468
rect 385 440 413 468
rect 441 440 469 468
rect 497 440 525 468
rect 539 440 567 468
rect 595 440 623 468
rect 651 440 679 468
rect 707 440 735 468
rect 763 440 791 468
rect 819 440 847 468
rect 875 440 903 468
rect 931 440 959 468
rect 987 440 1015 468
rect 1043 440 1071 468
rect 1085 440 1113 468
rect 1141 440 1169 468
rect 1197 440 1225 468
rect 1253 440 1281 468
rect 1309 440 1337 468
rect 1365 440 1393 468
rect 1421 440 1449 468
rect 1477 440 1505 468
rect 1533 440 1561 468
rect 1589 440 1617 468
rect 1631 440 1659 468
rect 1687 440 1715 468
rect 1743 440 1771 468
rect 1799 440 1827 468
rect 1855 440 1883 468
rect 1911 440 1939 468
rect 1967 440 1995 468
rect 2023 440 2051 468
rect 2079 440 2107 468
rect 2135 440 2163 468
rect -7 384 21 412
rect 49 384 77 412
rect 105 384 133 412
rect 161 384 189 412
rect 217 384 245 412
rect 273 384 301 412
rect 329 384 357 412
rect 385 384 413 412
rect 441 384 469 412
rect 497 384 525 412
rect 539 384 567 412
rect 595 384 623 412
rect 651 384 679 412
rect 707 384 735 412
rect 763 384 791 412
rect 819 384 847 412
rect 875 384 903 412
rect 931 384 959 412
rect 987 384 1015 412
rect 1043 384 1071 412
rect 1085 384 1113 412
rect 1141 384 1169 412
rect 1197 384 1225 412
rect 1253 384 1281 412
rect 1309 384 1337 412
rect 1365 384 1393 412
rect 1421 384 1449 412
rect 1477 384 1505 412
rect 1533 384 1561 412
rect 1589 384 1617 412
rect 1631 384 1659 412
rect 1687 384 1715 412
rect 1743 384 1771 412
rect 1799 384 1827 412
rect 1855 384 1883 412
rect 1911 384 1939 412
rect 1967 384 1995 412
rect 2023 384 2051 412
rect 2079 384 2107 412
rect 2135 384 2163 412
rect -7 328 21 356
rect 49 328 77 356
rect 105 328 133 356
rect 161 328 189 356
rect 217 328 245 356
rect 273 328 301 356
rect 329 328 357 356
rect 385 328 413 356
rect 441 328 469 356
rect 497 328 525 356
rect 539 328 567 356
rect 595 328 623 356
rect 651 328 679 356
rect 707 328 735 356
rect 763 328 791 356
rect 819 328 847 356
rect 875 328 903 356
rect 931 328 959 356
rect 987 328 1015 356
rect 1043 328 1071 356
rect 1085 328 1113 356
rect 1141 328 1169 356
rect 1197 328 1225 356
rect 1253 328 1281 356
rect 1309 328 1337 356
rect 1365 328 1393 356
rect 1421 328 1449 356
rect 1477 328 1505 356
rect 1533 328 1561 356
rect 1589 328 1617 356
rect 1631 328 1659 356
rect 1687 328 1715 356
rect 1743 328 1771 356
rect 1799 328 1827 356
rect 1855 328 1883 356
rect 1911 328 1939 356
rect 1967 328 1995 356
rect 2023 328 2051 356
rect 2079 328 2107 356
rect 2135 328 2163 356
rect -7 272 21 300
rect 49 272 77 300
rect 105 272 133 300
rect 161 272 189 300
rect 217 272 245 300
rect 273 272 301 300
rect 329 272 357 300
rect 385 272 413 300
rect 441 272 469 300
rect 497 272 525 300
rect 539 272 567 300
rect 595 272 623 300
rect 651 272 679 300
rect 707 272 735 300
rect 763 272 791 300
rect 819 272 847 300
rect 875 272 903 300
rect 931 272 959 300
rect 987 272 1015 300
rect 1043 272 1071 300
rect 1085 272 1113 300
rect 1141 272 1169 300
rect 1197 272 1225 300
rect 1253 272 1281 300
rect 1309 272 1337 300
rect 1365 272 1393 300
rect 1421 272 1449 300
rect 1477 272 1505 300
rect 1533 272 1561 300
rect 1589 272 1617 300
rect 1631 272 1659 300
rect 1687 272 1715 300
rect 1743 272 1771 300
rect 1799 272 1827 300
rect 1855 272 1883 300
rect 1911 272 1939 300
rect 1967 272 1995 300
rect 2023 272 2051 300
rect 2079 272 2107 300
rect 2135 272 2163 300
rect -7 216 21 244
rect 49 216 77 244
rect 105 216 133 244
rect 161 216 189 244
rect 217 216 245 244
rect 273 216 301 244
rect 329 216 357 244
rect 385 216 413 244
rect 441 216 469 244
rect 497 216 525 244
rect 539 216 567 244
rect 595 216 623 244
rect 651 216 679 244
rect 707 216 735 244
rect 763 216 791 244
rect 819 216 847 244
rect 875 216 903 244
rect 931 216 959 244
rect 987 216 1015 244
rect 1043 216 1071 244
rect 1085 216 1113 244
rect 1141 216 1169 244
rect 1197 216 1225 244
rect 1253 216 1281 244
rect 1309 216 1337 244
rect 1365 216 1393 244
rect 1421 216 1449 244
rect 1477 216 1505 244
rect 1533 216 1561 244
rect 1589 216 1617 244
rect 1631 216 1659 244
rect 1687 216 1715 244
rect 1743 216 1771 244
rect 1799 216 1827 244
rect 1855 216 1883 244
rect 1911 216 1939 244
rect 1967 216 1995 244
rect 2023 216 2051 244
rect 2079 216 2107 244
rect 2135 216 2163 244
rect -7 160 21 188
rect 49 160 77 188
rect 105 160 133 188
rect 161 160 189 188
rect 217 160 245 188
rect 273 160 301 188
rect 329 160 357 188
rect 385 160 413 188
rect 441 160 469 188
rect 497 160 525 188
rect 539 160 567 188
rect 595 160 623 188
rect 651 160 679 188
rect 707 160 735 188
rect 763 160 791 188
rect 819 160 847 188
rect 875 160 903 188
rect 931 160 959 188
rect 987 160 1015 188
rect 1043 160 1071 188
rect 1085 160 1113 188
rect 1141 160 1169 188
rect 1197 160 1225 188
rect 1253 160 1281 188
rect 1309 160 1337 188
rect 1365 160 1393 188
rect 1421 160 1449 188
rect 1477 160 1505 188
rect 1533 160 1561 188
rect 1589 160 1617 188
rect 1631 160 1659 188
rect 1687 160 1715 188
rect 1743 160 1771 188
rect 1799 160 1827 188
rect 1855 160 1883 188
rect 1911 160 1939 188
rect 1967 160 1995 188
rect 2023 160 2051 188
rect 2079 160 2107 188
rect 2135 160 2163 188
rect -7 104 21 132
rect 49 104 77 132
rect 105 104 133 132
rect 161 104 189 132
rect 217 104 245 132
rect 273 104 301 132
rect 329 104 357 132
rect 385 104 413 132
rect 441 104 469 132
rect 497 104 525 132
rect 539 104 567 132
rect 595 104 623 132
rect 651 104 679 132
rect 707 104 735 132
rect 763 104 791 132
rect 819 104 847 132
rect 875 104 903 132
rect 931 104 959 132
rect 987 104 1015 132
rect 1043 104 1071 132
rect 1085 104 1113 132
rect 1141 104 1169 132
rect 1197 104 1225 132
rect 1253 104 1281 132
rect 1309 104 1337 132
rect 1365 104 1393 132
rect 1421 104 1449 132
rect 1477 104 1505 132
rect 1533 104 1561 132
rect 1589 104 1617 132
rect 1631 104 1659 132
rect 1687 104 1715 132
rect 1743 104 1771 132
rect 1799 104 1827 132
rect 1855 104 1883 132
rect 1911 104 1939 132
rect 1967 104 1995 132
rect 2023 104 2051 132
rect 2079 104 2107 132
rect 2135 104 2163 132
rect -7 48 21 76
rect 49 48 77 76
rect 105 48 133 76
rect 161 48 189 76
rect 217 48 245 76
rect 273 48 301 76
rect 329 48 357 76
rect 385 48 413 76
rect 441 48 469 76
rect 497 48 525 76
rect 539 48 567 76
rect 595 48 623 76
rect 651 48 679 76
rect 707 48 735 76
rect 763 48 791 76
rect 819 48 847 76
rect 875 48 903 76
rect 931 48 959 76
rect 987 48 1015 76
rect 1043 48 1071 76
rect 1085 48 1113 76
rect 1141 48 1169 76
rect 1197 48 1225 76
rect 1253 48 1281 76
rect 1309 48 1337 76
rect 1365 48 1393 76
rect 1421 48 1449 76
rect 1477 48 1505 76
rect 1533 48 1561 76
rect 1589 48 1617 76
rect 1631 48 1659 76
rect 1687 48 1715 76
rect 1743 48 1771 76
rect 1799 48 1827 76
rect 1855 48 1883 76
rect 1911 48 1939 76
rect 1967 48 1995 76
rect 2023 48 2051 76
rect 2079 48 2107 76
rect 2135 48 2163 76
rect -7 6 21 20
rect -21 -8 21 6
rect 49 -8 77 20
rect 105 -8 133 20
rect 161 -8 189 20
rect 217 -8 245 20
rect 273 -8 301 20
rect 329 -8 357 20
rect 385 -8 413 20
rect 441 -8 469 20
rect 497 6 525 20
rect 539 6 567 20
rect 497 -8 567 6
rect 595 -8 623 20
rect 651 -8 679 20
rect 707 -8 735 20
rect 763 -8 791 20
rect 819 -8 847 20
rect 875 -8 903 20
rect 931 -8 959 20
rect 987 -8 1015 20
rect 1043 6 1071 20
rect 1085 6 1113 20
rect 1043 -8 1113 6
rect 1141 -8 1169 20
rect 1197 -8 1225 20
rect 1253 -8 1281 20
rect 1309 -8 1337 20
rect 1365 -8 1393 20
rect 1421 -8 1449 20
rect 1477 -8 1505 20
rect 1533 -8 1561 20
rect 1589 6 1617 20
rect 1631 6 1659 20
rect 1589 -8 1659 6
rect 1687 -8 1715 20
rect 1743 -8 1771 20
rect 1799 -8 1827 20
rect 1855 -8 1883 20
rect 1911 -8 1939 20
rect 1967 -8 1995 20
rect 2023 -8 2051 20
rect 2079 -8 2107 20
rect 2135 6 2163 20
rect 2135 -8 2177 6
rect -7 -22 7 -8
rect 511 -22 525 -8
rect 539 -22 553 -8
rect 1057 -22 1071 -8
rect 1085 -22 1099 -8
rect 1603 -22 1617 -8
rect 1631 -22 1645 -8
rect 2149 -22 2163 -8
rect -21 -36 21 -22
rect -7 -50 21 -36
rect 49 -50 77 -22
rect 105 -50 133 -22
rect 161 -50 189 -22
rect 217 -50 245 -22
rect 273 -50 301 -22
rect 329 -50 357 -22
rect 385 -50 413 -22
rect 441 -50 469 -22
rect 497 -36 567 -22
rect 497 -50 525 -36
rect 539 -50 567 -36
rect 595 -50 623 -22
rect 651 -50 679 -22
rect 707 -50 735 -22
rect 763 -50 791 -22
rect 819 -50 847 -22
rect 875 -50 903 -22
rect 931 -50 959 -22
rect 987 -50 1015 -22
rect 1043 -36 1113 -22
rect 1043 -50 1071 -36
rect 1085 -50 1113 -36
rect 1141 -50 1169 -22
rect 1197 -50 1225 -22
rect 1253 -50 1281 -22
rect 1309 -50 1337 -22
rect 1365 -50 1393 -22
rect 1421 -50 1449 -22
rect 1477 -50 1505 -22
rect 1533 -50 1561 -22
rect 1589 -36 1659 -22
rect 1589 -50 1617 -36
rect 1631 -50 1659 -36
rect 1687 -50 1715 -22
rect 1743 -50 1771 -22
rect 1799 -50 1827 -22
rect 1855 -50 1883 -22
rect 1911 -50 1939 -22
rect 1967 -50 1995 -22
rect 2023 -50 2051 -22
rect 2079 -50 2107 -22
rect 2135 -36 2177 -22
rect 2135 -50 2163 -36
rect -7 -106 21 -78
rect 49 -106 77 -78
rect 105 -106 133 -78
rect 161 -106 189 -78
rect 217 -106 245 -78
rect 273 -106 301 -78
rect 329 -106 357 -78
rect 385 -106 413 -78
rect 441 -106 469 -78
rect 497 -106 525 -78
rect 539 -106 567 -78
rect 595 -106 623 -78
rect 651 -106 679 -78
rect 707 -106 735 -78
rect 763 -106 791 -78
rect 819 -106 847 -78
rect 875 -106 903 -78
rect 931 -106 959 -78
rect 987 -106 1015 -78
rect 1043 -106 1071 -78
rect 1085 -106 1113 -78
rect 1141 -106 1169 -78
rect 1197 -106 1225 -78
rect 1253 -106 1281 -78
rect 1309 -106 1337 -78
rect 1365 -106 1393 -78
rect 1421 -106 1449 -78
rect 1477 -106 1505 -78
rect 1533 -106 1561 -78
rect 1589 -106 1617 -78
rect 1631 -106 1659 -78
rect 1687 -106 1715 -78
rect 1743 -106 1771 -78
rect 1799 -106 1827 -78
rect 1855 -106 1883 -78
rect 1911 -106 1939 -78
rect 1967 -106 1995 -78
rect 2023 -106 2051 -78
rect 2079 -106 2107 -78
rect 2135 -106 2163 -78
rect -7 -162 21 -134
rect 49 -162 77 -134
rect 105 -162 133 -134
rect 161 -162 189 -134
rect 217 -162 245 -134
rect 273 -162 301 -134
rect 329 -162 357 -134
rect 385 -162 413 -134
rect 441 -162 469 -134
rect 497 -162 525 -134
rect 539 -162 567 -134
rect 595 -162 623 -134
rect 651 -162 679 -134
rect 707 -162 735 -134
rect 763 -162 791 -134
rect 819 -162 847 -134
rect 875 -162 903 -134
rect 931 -162 959 -134
rect 987 -162 1015 -134
rect 1043 -162 1071 -134
rect 1085 -162 1113 -134
rect 1141 -162 1169 -134
rect 1197 -162 1225 -134
rect 1253 -162 1281 -134
rect 1309 -162 1337 -134
rect 1365 -162 1393 -134
rect 1421 -162 1449 -134
rect 1477 -162 1505 -134
rect 1533 -162 1561 -134
rect 1589 -162 1617 -134
rect 1631 -162 1659 -134
rect 1687 -162 1715 -134
rect 1743 -162 1771 -134
rect 1799 -162 1827 -134
rect 1855 -162 1883 -134
rect 1911 -162 1939 -134
rect 1967 -162 1995 -134
rect 2023 -162 2051 -134
rect 2079 -162 2107 -134
rect 2135 -162 2163 -134
rect -7 -218 21 -190
rect 49 -218 77 -190
rect 105 -218 133 -190
rect 161 -218 189 -190
rect 217 -218 245 -190
rect 273 -218 301 -190
rect 329 -218 357 -190
rect 385 -218 413 -190
rect 441 -218 469 -190
rect 497 -218 525 -190
rect 539 -218 567 -190
rect 595 -218 623 -190
rect 651 -218 679 -190
rect 707 -218 735 -190
rect 763 -218 791 -190
rect 819 -218 847 -190
rect 875 -218 903 -190
rect 931 -218 959 -190
rect 987 -218 1015 -190
rect 1043 -218 1071 -190
rect 1085 -218 1113 -190
rect 1141 -218 1169 -190
rect 1197 -218 1225 -190
rect 1253 -218 1281 -190
rect 1309 -218 1337 -190
rect 1365 -218 1393 -190
rect 1421 -218 1449 -190
rect 1477 -218 1505 -190
rect 1533 -218 1561 -190
rect 1589 -218 1617 -190
rect 1631 -218 1659 -190
rect 1687 -218 1715 -190
rect 1743 -218 1771 -190
rect 1799 -218 1827 -190
rect 1855 -218 1883 -190
rect 1911 -218 1939 -190
rect 1967 -218 1995 -190
rect 2023 -218 2051 -190
rect 2079 -218 2107 -190
rect 2135 -218 2163 -190
rect -7 -274 21 -246
rect 49 -274 77 -246
rect 105 -274 133 -246
rect 161 -274 189 -246
rect 217 -274 245 -246
rect 273 -274 301 -246
rect 329 -274 357 -246
rect 385 -274 413 -246
rect 441 -274 469 -246
rect 497 -274 525 -246
rect 539 -274 567 -246
rect 595 -274 623 -246
rect 651 -274 679 -246
rect 707 -274 735 -246
rect 763 -274 791 -246
rect 819 -274 847 -246
rect 875 -274 903 -246
rect 931 -274 959 -246
rect 987 -274 1015 -246
rect 1043 -274 1071 -246
rect 1085 -274 1113 -246
rect 1141 -274 1169 -246
rect 1197 -274 1225 -246
rect 1253 -274 1281 -246
rect 1309 -274 1337 -246
rect 1365 -274 1393 -246
rect 1421 -274 1449 -246
rect 1477 -274 1505 -246
rect 1533 -274 1561 -246
rect 1589 -274 1617 -246
rect 1631 -274 1659 -246
rect 1687 -274 1715 -246
rect 1743 -274 1771 -246
rect 1799 -274 1827 -246
rect 1855 -274 1883 -246
rect 1911 -274 1939 -246
rect 1967 -274 1995 -246
rect 2023 -274 2051 -246
rect 2079 -274 2107 -246
rect 2135 -274 2163 -246
rect -7 -330 21 -302
rect 49 -330 77 -302
rect 105 -330 133 -302
rect 161 -330 189 -302
rect 217 -330 245 -302
rect 273 -330 301 -302
rect 329 -330 357 -302
rect 385 -330 413 -302
rect 441 -330 469 -302
rect 497 -330 525 -302
rect 539 -330 567 -302
rect 595 -330 623 -302
rect 651 -330 679 -302
rect 707 -330 735 -302
rect 763 -330 791 -302
rect 819 -330 847 -302
rect 875 -330 903 -302
rect 931 -330 959 -302
rect 987 -330 1015 -302
rect 1043 -330 1071 -302
rect 1085 -330 1113 -302
rect 1141 -330 1169 -302
rect 1197 -330 1225 -302
rect 1253 -330 1281 -302
rect 1309 -330 1337 -302
rect 1365 -330 1393 -302
rect 1421 -330 1449 -302
rect 1477 -330 1505 -302
rect 1533 -330 1561 -302
rect 1589 -330 1617 -302
rect 1631 -330 1659 -302
rect 1687 -330 1715 -302
rect 1743 -330 1771 -302
rect 1799 -330 1827 -302
rect 1855 -330 1883 -302
rect 1911 -330 1939 -302
rect 1967 -330 1995 -302
rect 2023 -330 2051 -302
rect 2079 -330 2107 -302
rect 2135 -330 2163 -302
rect -7 -386 21 -358
rect 49 -386 77 -358
rect 105 -386 133 -358
rect 161 -386 189 -358
rect 217 -386 245 -358
rect 273 -386 301 -358
rect 329 -386 357 -358
rect 385 -386 413 -358
rect 441 -386 469 -358
rect 497 -386 525 -358
rect 539 -386 567 -358
rect 595 -386 623 -358
rect 651 -386 679 -358
rect 707 -386 735 -358
rect 763 -386 791 -358
rect 819 -386 847 -358
rect 875 -386 903 -358
rect 931 -386 959 -358
rect 987 -386 1015 -358
rect 1043 -386 1071 -358
rect 1085 -386 1113 -358
rect 1141 -386 1169 -358
rect 1197 -386 1225 -358
rect 1253 -386 1281 -358
rect 1309 -386 1337 -358
rect 1365 -386 1393 -358
rect 1421 -386 1449 -358
rect 1477 -386 1505 -358
rect 1533 -386 1561 -358
rect 1589 -386 1617 -358
rect 1631 -386 1659 -358
rect 1687 -386 1715 -358
rect 1743 -386 1771 -358
rect 1799 -386 1827 -358
rect 1855 -386 1883 -358
rect 1911 -386 1939 -358
rect 1967 -386 1995 -358
rect 2023 -386 2051 -358
rect 2079 -386 2107 -358
rect 2135 -386 2163 -358
rect -7 -442 21 -414
rect 49 -442 77 -414
rect 105 -442 133 -414
rect 161 -442 189 -414
rect 217 -442 245 -414
rect 273 -442 301 -414
rect 329 -442 357 -414
rect 385 -442 413 -414
rect 441 -442 469 -414
rect 497 -442 525 -414
rect 539 -442 567 -414
rect 595 -442 623 -414
rect 651 -442 679 -414
rect 707 -442 735 -414
rect 763 -442 791 -414
rect 819 -442 847 -414
rect 875 -442 903 -414
rect 931 -442 959 -414
rect 987 -442 1015 -414
rect 1043 -442 1071 -414
rect 1085 -442 1113 -414
rect 1141 -442 1169 -414
rect 1197 -442 1225 -414
rect 1253 -442 1281 -414
rect 1309 -442 1337 -414
rect 1365 -442 1393 -414
rect 1421 -442 1449 -414
rect 1477 -442 1505 -414
rect 1533 -442 1561 -414
rect 1589 -442 1617 -414
rect 1631 -442 1659 -414
rect 1687 -442 1715 -414
rect 1743 -442 1771 -414
rect 1799 -442 1827 -414
rect 1855 -442 1883 -414
rect 1911 -442 1939 -414
rect 1967 -442 1995 -414
rect 2023 -442 2051 -414
rect 2079 -442 2107 -414
rect 2135 -442 2163 -414
rect -7 -498 21 -470
rect 49 -498 77 -470
rect 105 -498 133 -470
rect 161 -498 189 -470
rect 217 -498 245 -470
rect 273 -498 301 -470
rect 329 -498 357 -470
rect 385 -498 413 -470
rect 441 -498 469 -470
rect 497 -498 525 -470
rect 539 -498 567 -470
rect 595 -498 623 -470
rect 651 -498 679 -470
rect 707 -498 735 -470
rect 763 -498 791 -470
rect 819 -498 847 -470
rect 875 -498 903 -470
rect 931 -498 959 -470
rect 987 -498 1015 -470
rect 1043 -498 1071 -470
rect 1085 -498 1113 -470
rect 1141 -498 1169 -470
rect 1197 -498 1225 -470
rect 1253 -498 1281 -470
rect 1309 -498 1337 -470
rect 1365 -498 1393 -470
rect 1421 -498 1449 -470
rect 1477 -498 1505 -470
rect 1533 -498 1561 -470
rect 1589 -498 1617 -470
rect 1631 -498 1659 -470
rect 1687 -498 1715 -470
rect 1743 -498 1771 -470
rect 1799 -498 1827 -470
rect 1855 -498 1883 -470
rect 1911 -498 1939 -470
rect 1967 -498 1995 -470
rect 2023 -498 2051 -470
rect 2079 -498 2107 -470
rect 2135 -498 2163 -470
rect -7 -540 21 -526
rect -21 -554 21 -540
rect 49 -554 77 -526
rect 105 -554 133 -526
rect 161 -554 189 -526
rect 217 -554 245 -526
rect 273 -554 301 -526
rect 329 -554 357 -526
rect 385 -554 413 -526
rect 441 -554 469 -526
rect 497 -540 525 -526
rect 539 -540 567 -526
rect 497 -554 567 -540
rect 595 -554 623 -526
rect 651 -554 679 -526
rect 707 -554 735 -526
rect 763 -554 791 -526
rect 819 -554 847 -526
rect 875 -554 903 -526
rect 931 -554 959 -526
rect 987 -554 1015 -526
rect 1043 -540 1071 -526
rect 1085 -540 1113 -526
rect 1043 -554 1113 -540
rect 1141 -554 1169 -526
rect 1197 -554 1225 -526
rect 1253 -554 1281 -526
rect 1309 -554 1337 -526
rect 1365 -554 1393 -526
rect 1421 -554 1449 -526
rect 1477 -554 1505 -526
rect 1533 -554 1561 -526
rect 1589 -540 1617 -526
rect 1631 -540 1659 -526
rect 1589 -554 1659 -540
rect 1687 -554 1715 -526
rect 1743 -554 1771 -526
rect 1799 -554 1827 -526
rect 1855 -554 1883 -526
rect 1911 -554 1939 -526
rect 1967 -554 1995 -526
rect 2023 -554 2051 -526
rect 2079 -554 2107 -526
rect 2135 -540 2163 -526
rect 2135 -554 2177 -540
rect -7 -568 7 -554
rect 511 -568 525 -554
rect 539 -568 553 -554
rect 1057 -568 1071 -554
rect 1085 -568 1099 -554
rect 1603 -568 1617 -554
rect 1631 -568 1645 -554
rect 2149 -568 2163 -554
<< end >>
