** sch_path: /home/yohanes/10-bit-DAC/xschem/res_seg_3.sch
**.subckt res_seg_3 v8 v7 v6 v5 v4 v3 v2 v1 v0 body
*.opin v8
*.opin v7
*.opin v6
*.opin v5
*.opin v4
*.opin v3
*.opin v2
*.opin v1
*.opin v0
*.ipin body
XR1 v7 v8 body sky130_fd_pr__res_xhigh_po_0p35 L=0.9486 mult=1 m=1
XR2 v6 v7 body sky130_fd_pr__res_xhigh_po_0p35 L=0.8888 mult=1 m=1
XR3 v5 v6 body sky130_fd_pr__res_xhigh_po_0p35 L=0.8460 mult=1 m=1
XR4 v4 v5 body sky130_fd_pr__res_xhigh_po_0p35 L=0.8118 mult=1 m=1
XR5 v3 v4 body sky130_fd_pr__res_xhigh_po_0p35 L=0.7691 mult=1 m=1
XR6 v2 v3 body sky130_fd_pr__res_xhigh_po_0p35 L=0.7349 mult=1 m=1
XR7 v1 v2 body sky130_fd_pr__res_xhigh_po_0p35 L=0.7178 mult=1 m=1
XR8 v0 v1 body sky130_fd_pr__res_xhigh_po_0p35 L=0.6922 mult=1 m=1
**.ends
.end
