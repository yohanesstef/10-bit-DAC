magic
tech sky130A
magscale 1 2
timestamp 1750166469
<< nwell >>
rect 1803 1303 5043 3335
<< mvnsubdiff >>
rect 1869 3209 4977 3269
rect 1869 1429 1929 3209
rect 4917 1429 4977 3209
rect 1869 1369 4977 1429
<< locali >>
rect 1882 3222 4964 3256
rect 1882 1416 1916 3222
rect 4930 1416 4964 3222
rect 1882 1382 4964 1416
<< metal1 >>
rect 1859 3199 4987 3279
rect 1859 1439 1939 3199
rect 1967 2989 2027 2995
rect 1967 1621 2027 2929
rect 1967 1555 2027 1561
rect 2055 2901 2115 2907
rect 2143 2841 2447 3199
rect 2882 2929 2888 2989
rect 2948 2929 2954 2989
rect 3892 2929 3898 2989
rect 3958 2929 3964 2989
rect 2764 2841 2770 2901
rect 2830 2841 2836 2901
rect 2055 1533 2115 2841
rect 2777 2684 2823 2841
rect 2895 2672 2941 2929
rect 3017 2525 3077 2531
rect 2559 2408 2701 2468
rect 2512 2261 2572 2267
rect 2512 2195 2572 2201
rect 2641 2173 2701 2408
rect 3017 2230 3077 2465
rect 3146 2437 3206 2443
rect 3146 2371 3206 2377
rect 3271 2355 3317 2420
rect 3393 2355 3453 2813
rect 3905 2672 3951 2929
rect 4010 2841 4016 2901
rect 4076 2841 4082 2901
rect 4399 2841 4703 3199
rect 4819 2989 4879 2995
rect 4731 2901 4791 2907
rect 4023 2672 4069 2841
rect 3640 2525 3700 2531
rect 3640 2459 3700 2465
rect 3769 2437 3829 2443
rect 3529 2355 3575 2408
rect 3264 2349 3324 2355
rect 3264 2283 3324 2289
rect 3393 2349 3582 2355
rect 3393 2289 3522 2349
rect 3393 2283 3582 2289
rect 3271 2230 3317 2283
rect 3017 2170 3153 2230
rect 2641 2107 2701 2113
rect 2055 1467 2115 1473
rect 2143 1439 2447 1797
rect 2777 1709 2823 1954
rect 2895 1797 2941 1954
rect 3393 1825 3453 2283
rect 3529 2230 3575 2283
rect 3769 2230 3829 2377
rect 4145 2408 4281 2468
rect 4145 2261 4205 2408
rect 3693 2170 3829 2230
rect 3899 2170 3911 2230
rect 4145 2195 4205 2201
rect 4274 2173 4334 2179
rect 4274 2107 4334 2113
rect 2882 1737 2888 1797
rect 2948 1737 2954 1797
rect 2764 1649 2770 1709
rect 2830 1649 2836 1709
rect 3905 1621 3951 1954
rect 3892 1561 3898 1621
rect 3958 1561 3964 1621
rect 4023 1533 4069 1954
rect 4010 1473 4016 1533
rect 4076 1473 4082 1533
rect 4399 1439 4703 1797
rect 4731 1709 4791 2841
rect 4819 1797 4879 2929
rect 4819 1731 4879 1737
rect 4731 1643 4791 1649
rect 4907 1439 4987 3199
rect 1859 1359 4987 1439
<< via1 >>
rect 1967 2929 2027 2989
rect 1967 1561 2027 1621
rect 2055 2841 2115 2901
rect 2888 2929 2948 2989
rect 3898 2929 3958 2989
rect 2770 2841 2830 2901
rect 2512 2201 2572 2261
rect 2641 2113 2701 2173
rect 3017 2465 3077 2525
rect 3146 2377 3206 2437
rect 4016 2841 4076 2901
rect 4819 2929 4879 2989
rect 4731 2841 4791 2901
rect 3640 2465 3700 2525
rect 3769 2377 3829 2437
rect 3264 2289 3324 2349
rect 3522 2289 3582 2349
rect 2055 1473 2115 1533
rect 4145 2201 4205 2261
rect 4274 2113 4334 2173
rect 2888 1737 2948 1797
rect 2770 1649 2830 1709
rect 3898 1561 3958 1621
rect 4016 1473 4076 1533
rect 4819 1737 4879 1797
rect 4731 1649 4791 1709
<< metal2 >>
rect 1961 2929 1967 2989
rect 2027 2929 2888 2989
rect 2948 2929 2954 2989
rect 3892 2929 3898 2989
rect 3958 2929 4819 2989
rect 4879 2929 4885 2989
rect 2049 2841 2055 2901
rect 2115 2841 2770 2901
rect 2830 2841 2836 2901
rect 4010 2841 4016 2901
rect 4076 2841 4731 2901
rect 4791 2841 4797 2901
rect 3011 2465 3017 2525
rect 3077 2465 3640 2525
rect 3700 2465 3706 2525
rect 3140 2377 3146 2437
rect 3206 2377 3769 2437
rect 3829 2377 3835 2437
rect 3258 2289 3264 2349
rect 3324 2289 3330 2349
rect 3516 2289 3522 2349
rect 3582 2289 3588 2349
rect 2506 2201 2512 2261
rect 2572 2201 4145 2261
rect 4205 2201 4211 2261
rect 2635 2113 2641 2173
rect 2701 2113 4274 2173
rect 4334 2113 4340 2173
rect 2882 1737 2888 1797
rect 2948 1737 4819 1797
rect 4879 1737 4885 1797
rect 2764 1649 2770 1709
rect 2830 1649 4731 1709
rect 4791 1649 4797 1709
rect 1961 1561 1967 1621
rect 2027 1561 3898 1621
rect 3958 1561 3964 1621
rect 2027 1473 2055 1533
rect 2115 1473 4016 1533
rect 4076 1473 4082 1533
use cm2_pcell2_5  cm2_pcell2_5_0
timestamp 1750163329
transform 1 0 3325 0 1 2116
box -1254 184 1450 725
use cm2_pcell2_5  cm2_pcell2_5_1
timestamp 1750163329
transform 1 0 3325 0 -1 2522
box -1254 184 1450 725
<< labels >>
flabel metal1 s 3264 2289 3324 2349 0 FreeSans 480 0 0 0 S0
port 0 nsew
flabel metal2 s 3898 2929 3958 2989 0 FreeSans 480 0 0 0 S1
port 1 nsew
flabel metal2 s 2888 2929 2948 2989 0 FreeSans 480 0 0 0 S2
port 2 nsew
flabel metal2 s 4016 2841 4076 2901 0 FreeSans 480 0 0 0 S3
port 3 nsew
flabel metal2 s 2770 2841 2830 2901 0 FreeSans 480 0 0 0 S4
port 4 nsew
flabel metal2 s 3522 2289 3582 2349 0 FreeSans 480 0 0 0 D0
port 5 nsew
flabel metal2 s 3017 2465 3077 2525 0 FreeSans 480 0 0 0 D1
port 6 nsew
flabel metal2 s 3146 2377 3206 2437 0 FreeSans 480 0 0 0 D2
port 7 nsew
flabel metal2 s 2512 2201 2572 2261 0 FreeSans 480 0 0 0 D3
port 8 nsew
flabel metal2 s 2641 2113 2701 2173 0 FreeSans 480 0 0 0 D4
port 9 nsew
flabel locali s 1882 1382 1916 1416 0 FreeSans 480 0 0 0 VDDA
port 10 nsew
<< end >>
