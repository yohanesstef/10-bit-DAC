** sch_path: /home/yohanes/10-bit-DAC/xschem/diff_pair.sch
.subckt dp_nmos P_IN N_IN I_ONA I_ONB I_TAIL VNB
*.PININFO I_OPA:O I_OPB:O P_IN:I N_IN:I I_ONA:O I_ONB:O I_HEAD:I I_TAIL:I VPB:I VNB:I
XM3 I_ONA P_IN I_TAIL VNB sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=4
XM4 I_ONB N_IN I_TAIL VNB sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=4
.ends
