magic
tech sky130A
magscale 1 2
timestamp 1750900893
<< error_s >>
rect 2014 788 2020 794
rect 2068 788 2074 794
rect 2008 782 2014 788
rect 2074 782 2080 788
rect 2008 728 2014 734
rect 2074 728 2080 734
rect 2014 722 2020 728
rect 2068 722 2074 728
rect 1434 700 1440 706
rect 1488 700 1494 706
rect 1738 700 1744 706
rect 1792 700 1798 706
rect 1428 694 1434 700
rect 1494 694 1500 700
rect 1732 694 1738 700
rect 1798 694 1804 700
rect 1428 640 1434 646
rect 1494 640 1500 646
rect 1732 640 1738 646
rect 1798 640 1804 646
rect 1434 634 1440 640
rect 1488 634 1494 640
rect 1738 634 1744 640
rect 1792 634 1798 640
rect 854 612 860 618
rect 908 612 914 618
rect 1158 612 1164 618
rect 1212 612 1218 618
rect 848 606 854 612
rect 914 606 920 612
rect 1152 606 1158 612
rect 1218 606 1224 612
rect 848 552 854 558
rect 914 552 920 558
rect 1152 552 1158 558
rect 1218 552 1224 558
rect 854 546 860 552
rect 908 546 914 552
rect 1158 546 1164 552
rect 1212 546 1218 552
rect 274 524 280 530
rect 328 524 334 530
rect 578 524 584 530
rect 632 524 638 530
rect 268 518 274 524
rect 334 518 340 524
rect 572 518 578 524
rect 638 518 644 524
rect 268 464 274 470
rect 334 464 340 470
rect 572 464 578 470
rect 638 464 644 470
rect 274 458 280 464
rect 328 458 334 464
rect 578 458 584 464
rect 632 458 638 464
rect -2 436 4 442
rect 52 436 58 442
rect -8 430 -2 436
rect 58 430 64 436
rect -8 376 -2 382
rect 58 376 64 382
rect -2 370 4 376
rect 52 370 58 376
<< pwell >>
rect -156 -189 2416 349
<< mvpsubdiff >>
rect -120 301 2380 313
rect -120 267 -12 301
rect 2272 267 2380 301
rect -120 255 2380 267
rect -120 205 -62 255
rect -120 -45 -108 205
rect -74 -45 -62 205
rect -120 -95 -62 -45
rect 2322 205 2380 255
rect 2322 -45 2334 205
rect 2368 -45 2380 205
rect 2322 -95 2380 -45
rect -120 -107 2380 -95
rect -120 -141 -12 -107
rect 2272 -141 2380 -107
rect -120 -153 2380 -141
<< mvpsubdiffcont >>
rect -12 267 2272 301
rect -108 -45 -74 205
rect 2334 -45 2368 205
rect -12 -141 2272 -107
<< locali >>
rect -108 267 -12 301
rect 2272 267 2368 301
rect -108 205 -74 267
rect -108 -107 -74 -45
rect 2334 205 2368 267
rect 2334 -107 2368 -45
rect -108 -141 -12 -107
rect 2272 -141 2368 -107
<< metal1 >>
rect 2014 788 2074 794
rect 1434 700 1494 706
rect 854 612 914 618
rect 274 524 334 530
rect -2 436 58 442
rect -2 197 58 376
rect 186 436 246 442
rect 186 197 246 376
rect -2 95 48 197
rect 196 95 246 197
rect -2 7 58 95
rect 186 7 246 95
rect 274 197 334 464
rect 578 524 638 530
rect 462 348 522 354
rect 462 197 522 288
rect 274 95 324 197
rect 472 95 522 197
rect 274 7 334 95
rect 462 7 522 95
rect 578 197 638 464
rect 766 436 826 442
rect 766 197 826 376
rect 578 95 628 197
rect 776 95 826 197
rect 578 7 638 95
rect 766 7 826 95
rect 854 198 914 552
rect 1158 612 1218 618
rect 1042 524 1102 530
rect 1042 348 1102 464
rect 854 96 904 198
rect 1042 197 1102 288
rect 854 7 914 96
rect 1052 95 1102 197
rect 1042 7 1102 95
rect 1158 197 1218 552
rect 1346 436 1406 442
rect 1346 197 1406 376
rect 1158 95 1208 197
rect 1356 95 1406 197
rect 1158 7 1218 95
rect 1346 7 1406 95
rect 1434 197 1494 640
rect 1738 700 1798 706
rect 1622 524 1682 530
rect 1622 197 1682 464
rect 1434 95 1484 197
rect 1632 95 1682 197
rect 1434 7 1494 95
rect 1622 7 1682 95
rect 1738 197 1798 640
rect 1926 436 1986 442
rect 1926 197 1986 376
rect 1738 95 1788 197
rect 1936 95 1986 197
rect 1738 7 1798 95
rect 1926 7 1986 95
rect 2014 197 2074 728
rect 2202 524 2262 530
rect 2202 197 2262 464
rect 2014 95 2064 197
rect 2212 95 2262 197
rect 2014 7 2074 95
rect 2202 7 2262 95
<< via1 >>
rect 2014 728 2074 788
rect 1434 640 1494 700
rect 854 552 914 612
rect 274 464 334 524
rect -2 376 58 436
rect 186 376 246 436
rect 578 464 638 524
rect 462 288 522 348
rect 766 376 826 436
rect 1158 552 1218 612
rect 1042 464 1102 524
rect 1042 288 1102 348
rect 1346 376 1406 436
rect 1738 640 1798 700
rect 1622 464 1682 524
rect 1926 376 1986 436
rect 2202 464 2262 524
<< metal2 >>
rect 1036 464 1042 524
rect 1102 464 1622 524
rect 1682 464 2202 524
rect 2262 464 2268 524
rect 180 376 186 436
rect 246 376 766 436
rect 826 376 1346 436
rect 1406 376 1926 436
rect 1986 376 1992 436
rect 455 288 462 348
rect 522 288 1042 348
rect 1102 288 1108 348
use hnmos_2  hnmos_2_0
timestamp 1750900893
transform 1 0 -12 0 1 -20
box -4 1 548 199
use hnmos_2  hnmos_2_1
timestamp 1750900893
transform 1 0 568 0 1 -20
box -4 1 548 199
use hnmos_2  hnmos_2_2
timestamp 1750900893
transform 1 0 1148 0 1 -20
box -4 1 548 199
use hnmos_2  hnmos_2_3
timestamp 1750900893
transform 1 0 1728 0 1 -20
box -4 1 548 199
<< end >>
