magic
tech sky130A
magscale 1 2
timestamp 1749834095
<< magnet >>
rect 1829 4813 1857 4841
rect 2653 4813 2681 4841
rect 2709 4813 2737 4841
rect 3533 4813 3561 4841
rect 1801 4785 1889 4813
rect 1829 4753 1889 4785
rect 1917 4753 1977 4813
rect 2005 4753 2065 4813
rect 2093 4753 2153 4813
rect 2181 4753 2241 4813
rect 2269 4753 2329 4813
rect 2357 4753 2417 4813
rect 2445 4753 2505 4813
rect 2533 4753 2593 4813
rect 2621 4785 2769 4813
rect 2621 4753 2681 4785
rect 2709 4753 2769 4785
rect 2797 4753 2857 4813
rect 2885 4753 2945 4813
rect 2973 4753 3033 4813
rect 3061 4753 3121 4813
rect 3149 4753 3209 4813
rect 3237 4753 3297 4813
rect 3325 4753 3385 4813
rect 3413 4753 3473 4813
rect 3501 4785 3589 4813
rect 3501 4753 3561 4785
rect 1829 4665 1889 4725
rect 1917 4665 1977 4725
rect 2005 4665 2065 4725
rect 2093 4665 2153 4725
rect 2181 4665 2241 4725
rect 2269 4665 2329 4725
rect 2357 4665 2417 4725
rect 2445 4665 2505 4725
rect 2533 4665 2593 4725
rect 2621 4665 2681 4725
rect 2709 4665 2769 4725
rect 2797 4665 2857 4725
rect 2885 4665 2945 4725
rect 2973 4665 3033 4725
rect 3061 4665 3121 4725
rect 3149 4665 3209 4725
rect 3237 4665 3297 4725
rect 3325 4665 3385 4725
rect 3413 4665 3473 4725
rect 3501 4665 3561 4725
rect 1829 4577 1889 4637
rect 1917 4577 1977 4637
rect 2005 4577 2065 4637
rect 2093 4577 2153 4637
rect 2181 4577 2241 4637
rect 2269 4577 2329 4637
rect 2357 4577 2417 4637
rect 2445 4577 2505 4637
rect 2533 4577 2593 4637
rect 2621 4577 2681 4637
rect 2709 4577 2769 4637
rect 2797 4577 2857 4637
rect 2885 4577 2945 4637
rect 2973 4577 3033 4637
rect 3061 4577 3121 4637
rect 3149 4577 3209 4637
rect 3237 4577 3297 4637
rect 3325 4577 3385 4637
rect 3413 4577 3473 4637
rect 3501 4577 3561 4637
rect 1829 4489 1889 4549
rect 1917 4489 1977 4549
rect 2005 4489 2065 4549
rect 2093 4489 2153 4549
rect 2181 4489 2241 4549
rect 2269 4489 2329 4549
rect 2357 4489 2417 4549
rect 2445 4489 2505 4549
rect 2533 4489 2593 4549
rect 2621 4489 2681 4549
rect 2709 4489 2769 4549
rect 2797 4489 2857 4549
rect 2885 4489 2945 4549
rect 2973 4489 3033 4549
rect 3061 4489 3121 4549
rect 3149 4489 3209 4549
rect 3237 4489 3297 4549
rect 3325 4489 3385 4549
rect 3413 4489 3473 4549
rect 3501 4489 3561 4549
rect 1829 4401 1889 4461
rect 1917 4401 1977 4461
rect 2005 4401 2065 4461
rect 2093 4401 2153 4461
rect 2181 4401 2241 4461
rect 2269 4401 2329 4461
rect 2357 4401 2417 4461
rect 2445 4401 2505 4461
rect 2533 4401 2593 4461
rect 2621 4401 2681 4461
rect 2709 4401 2769 4461
rect 2797 4401 2857 4461
rect 2885 4401 2945 4461
rect 2973 4401 3033 4461
rect 3061 4401 3121 4461
rect 3149 4401 3209 4461
rect 3237 4401 3297 4461
rect 3325 4401 3385 4461
rect 3413 4401 3473 4461
rect 3501 4401 3561 4461
rect 1829 4313 1889 4373
rect 1917 4313 1977 4373
rect 2005 4313 2065 4373
rect 2093 4313 2153 4373
rect 2181 4313 2241 4373
rect 2269 4313 2329 4373
rect 2357 4313 2417 4373
rect 2445 4313 2505 4373
rect 2533 4313 2593 4373
rect 2621 4313 2681 4373
rect 2709 4313 2769 4373
rect 2797 4313 2857 4373
rect 2885 4313 2945 4373
rect 2973 4313 3033 4373
rect 3061 4313 3121 4373
rect 3149 4313 3209 4373
rect 3237 4313 3297 4373
rect 3325 4313 3385 4373
rect 3413 4313 3473 4373
rect 3501 4313 3561 4373
rect 1829 4225 1889 4285
rect 1917 4225 1977 4285
rect 2005 4225 2065 4285
rect 2093 4225 2153 4285
rect 2181 4225 2241 4285
rect 2269 4225 2329 4285
rect 2357 4225 2417 4285
rect 2445 4225 2505 4285
rect 2533 4225 2593 4285
rect 2621 4225 2681 4285
rect 2709 4225 2769 4285
rect 2797 4225 2857 4285
rect 2885 4225 2945 4285
rect 2973 4225 3033 4285
rect 3061 4225 3121 4285
rect 3149 4225 3209 4285
rect 3237 4225 3297 4285
rect 3325 4225 3385 4285
rect 3413 4225 3473 4285
rect 3501 4225 3561 4285
rect 1829 4137 1889 4197
rect 1917 4137 1977 4197
rect 2005 4137 2065 4197
rect 2093 4137 2153 4197
rect 2181 4137 2241 4197
rect 2269 4137 2329 4197
rect 2357 4137 2417 4197
rect 2445 4137 2505 4197
rect 2533 4137 2593 4197
rect 2621 4137 2681 4197
rect 2709 4137 2769 4197
rect 2797 4137 2857 4197
rect 2885 4137 2945 4197
rect 2973 4137 3033 4197
rect 3061 4137 3121 4197
rect 3149 4137 3209 4197
rect 3237 4137 3297 4197
rect 3325 4137 3385 4197
rect 3413 4137 3473 4197
rect 3501 4137 3561 4197
rect 1829 4049 1889 4109
rect 1917 4049 1977 4109
rect 2005 4049 2065 4109
rect 2093 4049 2153 4109
rect 2181 4049 2241 4109
rect 2269 4049 2329 4110
rect 2357 4049 2417 4109
rect 2445 4049 2505 4109
rect 2533 4049 2593 4109
rect 2621 4049 2681 4110
rect 2709 4049 2769 4110
rect 2797 4049 2857 4109
rect 2885 4049 2945 4109
rect 2973 4049 3033 4109
rect 3061 4049 3121 4109
rect 3149 4049 3209 4110
rect 3237 4049 3297 4109
rect 3325 4049 3385 4109
rect 3413 4049 3473 4109
rect 3501 4048 3561 4109
rect 1829 3989 1889 4021
rect 1801 3961 1889 3989
rect 1917 3961 1977 4021
rect 2005 3961 2065 4021
rect 2093 3961 2153 4021
rect 2181 3961 2241 4021
rect 2269 3961 2329 4021
rect 2357 3961 2417 4021
rect 2445 3961 2505 4021
rect 2533 3961 2593 4021
rect 2621 3989 2681 4021
rect 2709 3989 2769 4021
rect 2621 3961 2769 3989
rect 2797 3961 2857 4021
rect 2885 3961 2945 4021
rect 2973 3961 3033 4021
rect 3061 3961 3121 4021
rect 3149 3961 3209 4021
rect 3237 3961 3297 4021
rect 3325 3961 3385 4021
rect 3413 3961 3473 4021
rect 3501 3989 3561 4021
rect 3501 3961 3589 3989
rect 1829 3933 1857 3961
rect 2653 3933 2681 3961
rect 2709 3933 2737 3961
rect 3533 3933 3561 3961
rect 1801 3905 1889 3933
rect 1829 3873 1889 3905
rect 1917 3873 1977 3933
rect 2005 3873 2065 3933
rect 2093 3873 2153 3933
rect 2181 3873 2241 3933
rect 2269 3873 2329 3933
rect 2357 3873 2417 3933
rect 2445 3873 2505 3933
rect 2533 3873 2593 3933
rect 2621 3905 2769 3933
rect 2621 3873 2681 3905
rect 2709 3873 2769 3905
rect 2797 3873 2857 3933
rect 2885 3873 2945 3933
rect 2973 3873 3033 3933
rect 3061 3873 3121 3933
rect 3149 3873 3209 3933
rect 3237 3873 3297 3933
rect 3325 3873 3385 3933
rect 3413 3873 3473 3933
rect 3501 3905 3589 3933
rect 3501 3873 3561 3905
rect 1829 3785 1889 3845
rect 1917 3785 1977 3845
rect 2005 3785 2065 3845
rect 2093 3785 2153 3845
rect 2181 3785 2241 3845
rect 2269 3785 2329 3845
rect 2357 3785 2417 3845
rect 2445 3785 2505 3845
rect 2533 3785 2593 3845
rect 2621 3785 2681 3845
rect 2709 3785 2769 3845
rect 2797 3785 2857 3845
rect 2885 3785 2945 3845
rect 2973 3785 3033 3845
rect 3061 3785 3121 3845
rect 3149 3785 3209 3845
rect 3237 3785 3297 3845
rect 3325 3785 3385 3845
rect 3413 3785 3473 3845
rect 3501 3785 3561 3845
rect 1829 3697 1889 3757
rect 1917 3697 1977 3757
rect 2005 3697 2065 3757
rect 2093 3697 2153 3757
rect 2181 3697 2241 3757
rect 2269 3697 2329 3757
rect 2357 3697 2417 3757
rect 2445 3697 2505 3757
rect 2533 3697 2593 3757
rect 2621 3697 2681 3757
rect 2709 3697 2769 3757
rect 2797 3697 2857 3757
rect 2885 3697 2945 3757
rect 2973 3697 3033 3757
rect 3061 3697 3121 3757
rect 3149 3697 3209 3757
rect 3237 3697 3297 3757
rect 3325 3697 3385 3757
rect 3413 3697 3473 3757
rect 3501 3697 3561 3757
rect 1829 3609 1889 3669
rect 1917 3609 1977 3669
rect 2005 3609 2065 3669
rect 2093 3609 2153 3669
rect 2181 3609 2241 3669
rect 2269 3609 2329 3669
rect 2357 3609 2417 3669
rect 2445 3609 2505 3669
rect 2533 3609 2593 3669
rect 2621 3609 2681 3669
rect 2709 3609 2769 3669
rect 2797 3609 2857 3669
rect 2885 3609 2945 3669
rect 2973 3609 3033 3669
rect 3061 3609 3121 3669
rect 3149 3609 3209 3669
rect 3237 3609 3297 3669
rect 3325 3609 3385 3669
rect 3413 3609 3473 3669
rect 3501 3609 3561 3669
rect 1829 3521 1889 3581
rect 1917 3521 1977 3581
rect 2005 3521 2065 3581
rect 2093 3521 2153 3581
rect 2181 3521 2241 3581
rect 2269 3521 2329 3581
rect 2357 3521 2417 3581
rect 2445 3521 2505 3581
rect 2533 3521 2593 3581
rect 2621 3521 2681 3581
rect 2709 3521 2769 3581
rect 2797 3521 2857 3581
rect 2885 3521 2945 3581
rect 2973 3521 3033 3581
rect 3061 3521 3121 3581
rect 3149 3521 3209 3581
rect 3237 3521 3297 3581
rect 3325 3521 3385 3581
rect 3413 3521 3473 3581
rect 3501 3521 3561 3581
rect 1829 3433 1889 3493
rect 1917 3433 1977 3493
rect 2005 3433 2065 3493
rect 2093 3433 2153 3493
rect 2181 3433 2241 3493
rect 2269 3433 2329 3493
rect 2357 3433 2417 3493
rect 2445 3433 2505 3493
rect 2533 3433 2593 3493
rect 2621 3433 2681 3493
rect 2709 3433 2769 3493
rect 2797 3433 2857 3493
rect 2885 3433 2945 3493
rect 2973 3433 3033 3493
rect 3061 3433 3121 3493
rect 3149 3433 3209 3493
rect 3237 3433 3297 3493
rect 3325 3433 3385 3493
rect 3413 3433 3473 3493
rect 3501 3433 3561 3493
rect 1829 3345 1889 3405
rect 1917 3345 1977 3405
rect 2005 3345 2065 3405
rect 2093 3345 2153 3405
rect 2181 3345 2241 3405
rect 2269 3345 2329 3405
rect 2357 3345 2417 3405
rect 2445 3345 2505 3405
rect 2533 3345 2593 3405
rect 2621 3345 2681 3405
rect 2709 3345 2769 3405
rect 2797 3345 2857 3405
rect 2885 3345 2945 3405
rect 2973 3345 3033 3405
rect 3061 3345 3121 3405
rect 3149 3345 3209 3405
rect 3237 3345 3297 3405
rect 3325 3345 3385 3405
rect 3413 3345 3473 3405
rect 3501 3345 3561 3405
rect 1829 3257 1889 3317
rect 1917 3257 1977 3317
rect 2005 3257 2065 3317
rect 2093 3257 2153 3317
rect 2181 3257 2241 3317
rect 2269 3257 2329 3317
rect 2357 3257 2417 3317
rect 2445 3257 2505 3317
rect 2533 3257 2593 3317
rect 2621 3257 2681 3317
rect 2709 3257 2769 3317
rect 2797 3257 2857 3317
rect 2885 3257 2945 3317
rect 2973 3257 3033 3317
rect 3061 3257 3121 3317
rect 3149 3257 3209 3317
rect 3237 3257 3297 3317
rect 3325 3257 3385 3317
rect 3413 3257 3473 3317
rect 3501 3257 3561 3317
rect 1829 3169 1889 3229
rect 1917 3168 1977 3228
rect 2005 3168 2065 3228
rect 2093 3168 2153 3228
rect 2181 3168 2241 3228
rect 2269 3168 2329 3229
rect 2357 3168 2417 3228
rect 2445 3168 2505 3228
rect 2533 3168 2593 3228
rect 2621 3168 2681 3229
rect 2709 3168 2769 3229
rect 2797 3168 2857 3228
rect 2885 3168 2945 3228
rect 2973 3168 3033 3228
rect 3061 3168 3121 3228
rect 3149 3168 3209 3229
rect 3237 3168 3297 3228
rect 3325 3168 3385 3228
rect 3413 3168 3473 3228
rect 3501 3168 3561 3229
rect 1829 3109 1889 3141
rect 1801 3081 1889 3109
rect 1917 3081 1977 3141
rect 2005 3081 2065 3141
rect 2093 3081 2153 3141
rect 2181 3081 2241 3141
rect 2269 3081 2329 3141
rect 2357 3081 2417 3141
rect 2445 3081 2505 3141
rect 2533 3081 2593 3141
rect 2621 3109 2681 3141
rect 2709 3109 2769 3141
rect 2621 3081 2769 3109
rect 2797 3081 2857 3141
rect 2885 3081 2945 3141
rect 2973 3081 3033 3141
rect 3061 3081 3121 3141
rect 3149 3081 3209 3141
rect 3237 3081 3297 3141
rect 3325 3081 3385 3141
rect 3413 3081 3473 3141
rect 3501 3109 3561 3141
rect 3501 3081 3589 3109
rect 1829 3053 1857 3081
rect 2653 3053 2681 3081
rect 2709 3053 2737 3081
rect 3533 3053 3561 3081
<< end >>
