magic
tech sky130A
magscale 1 2
timestamp 1749890363
<< error_s >>
rect 11 8 41 496
rect 77 74 107 430
rect 1491 74 1521 430
rect 77 70 393 74
rect 453 70 769 74
rect 829 70 1145 74
rect 1205 70 1521 74
rect 1557 8 1587 496
rect 11 4 1587 8
<< metal2 >>
rect 47 457 1551 517
use cm_pcell1_2  cm_pcell1_2_0
timestamp 1749889584
transform 1 0 13 0 1 22
box -2 -18 822 508
use cm_pcell1_2  cm_pcell1_2_1
timestamp 1749889584
transform 1 0 765 0 1 22
box -2 -18 822 508
<< end >>
