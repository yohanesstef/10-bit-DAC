magic
tech sky130A
magscale 1 2
timestamp 1749399058
<< error_p >>
rect 240 4692 270 4904
rect 306 4758 336 4838
rect 4632 4758 4662 4838
rect 306 4754 522 4758
rect 582 4754 798 4758
rect 858 4754 1074 4758
rect 1134 4754 1188 4758
rect 3780 4754 3834 4758
rect 3894 4754 4110 4758
rect 4170 4754 4386 4758
rect 4446 4754 4662 4758
rect 4698 4692 4728 4904
rect 240 4688 1188 4692
rect 3780 4688 4728 4692
<< error_s >>
rect 1188 4754 1350 4758
rect 1410 4754 1626 4758
rect 1686 4754 1902 4758
rect 1962 4754 2178 4758
rect 2238 4754 2454 4758
rect 2514 4754 2730 4758
rect 2790 4754 3006 4758
rect 3066 4754 3282 4758
rect 3342 4754 3558 4758
rect 3618 4754 3780 4758
rect 1188 4688 3780 4692
use hpmos_8  hpmos_8_0
timestamp 1749386853
transform 1 0 -121 0 1 4700
box 361 -12 2641 238
use hpmos_8  hpmos_8_1
timestamp 1749386853
transform 1 0 2087 0 1 4700
box 361 -12 2641 238
<< end >>
