* PEX produced on Fri Jun  6 20:48:16 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from rseg_1_v3.ext - technology: sky130A

.subckt rseg_1_v3 v0 v1 v2 v3 v4 v5 v6 v7 v8 v9 v10 v11 v12 v13 v14 v15 v16 v17 v18
+ v19 v20 v21 v22 v23 v24 v25 v26 v27 v28 v29 v30 v31 v32 v33 v34 v35 v36 v37 v38
+ v39 v40 v41 v42 v43 v44 v45 v46 v47 v48 v49 v50 v51 v52 v53 v54 v55 v56 v57 v58
+ v59 v60 v61 v62 v63 v64 gnd
X0 gnd.t1 gnd.t2 gnd.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X1 v49.t1 v50.t1 gnd.t10 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X2 gnd.t30 gnd.t31 gnd.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X3 gnd.t38 gnd.t39 gnd.t0 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X4 v49.t0 v48.t1 gnd.t10 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X5 v3.t1 v4.t1 gnd.t7 sky130_fd_pr__res_xhigh_po_1p41 l=3.37
X6 v27.t0 v28.t1 gnd.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X7 v23.t0 v22.t0 gnd.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X8 gnd.t26 gnd.t27 gnd.t10 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X9 v47.t0 v48.t0 gnd.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X10 v55.t1 v54.t0 gnd.t10 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X11 v33.t1 v32.t1 gnd.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X12 v63.t1 v62.t1 gnd.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X13 gnd.t36 gnd.t37 gnd.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X14 v25.t1 v24.t1 gnd.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X15 gnd.t24 gnd.t25 gnd.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X16 v27.t1 v26.t1 gnd.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X17 gnd.t13 gnd.t14 gnd.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X18 v17.t1 v18.t0 gnd.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X19 v37.t0 v36.t1 gnd.t0 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X20 v23.t1 v24.t0 gnd.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X21 v39.t0 v40.t1 gnd.t0 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X22 v63.t0 v64.t0 gnd.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X23 v21.t1 v20.t0 gnd.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X24 v5.t0 v6.t0 gnd.t7 sky130_fd_pr__res_xhigh_po_1p41 l=2.86
X25 v55.t0 v56.t0 gnd.t10 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X26 v9.t1 v10.t0 gnd.t17 sky130_fd_pr__res_xhigh_po_1p41 l=2.19
X27 gnd.t22 gnd.t23 gnd.t17 sky130_fd_pr__res_xhigh_po_1p41 l=1.68
X28 v29.t0 v28.t0 gnd.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X29 v41.t1 v42.t0 gnd.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X30 v17.t0 v16.t0 gnd.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X31 v21.t0 v22.t1 gnd.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X32 v41.t0 v40.t0 gnd.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X33 v57.t1 v58.t1 gnd.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X34 v31.t1 v30.t1 gnd.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X35 v11.t0 v12.t1 gnd.t17 sky130_fd_pr__res_xhigh_po_1p41 l=1.99
X36 v53.t0 v52.t0 gnd.t10 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X37 gnd.t15 gnd.t16 gnd.t7 sky130_fd_pr__res_xhigh_po_1p41 l=2.5
X38 gnd.t28 gnd.t29 gnd.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X39 v15.t1 v16.t1 gnd.t17 sky130_fd_pr__res_xhigh_po_1p41 l=1.68
X40 v13.t0 v12.t0 gnd.t17 sky130_fd_pr__res_xhigh_po_1p41 l=1.89
X41 v5.t1 v4.t0 gnd.t7 sky130_fd_pr__res_xhigh_po_1p41 l=3.12
X42 v1.t0 v2.t0 gnd.t7 sky130_fd_pr__res_xhigh_po_1p41 l=4.24
X43 gnd.t34 gnd.t35 gnd.t17 sky130_fd_pr__res_xhigh_po_1p41 l=2.35
X44 v29.t1 v30.t0 gnd.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X45 v43.t1 v42.t1 gnd.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X46 v53.t1 v54.t1 gnd.t10 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X47 v15.t0 v14.t1 gnd.t17 sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X48 v45.t0 v44.t1 gnd.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X49 v31.t0 v32.t0 gnd.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X50 v37.t1 v38.t1 gnd.t0 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X51 gnd.t18 gnd.t19 gnd.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X52 v35.t0 v36.t0 gnd.t0 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X53 v11.t1 v10.t1 gnd.t17 sky130_fd_pr__res_xhigh_po_1p41 l=2.09
X54 v7.t1 v8.t1 gnd.t7 sky130_fd_pr__res_xhigh_po_1p41 l=2.5
X55 gnd.t8 gnd.t9 gnd.t7 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X56 v3.t0 v2.t1 gnd.t7 sky130_fd_pr__res_xhigh_po_1p41 l=3.73
X57 v43.t0 v44.t0 gnd.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X58 v7.t0 v6.t1 gnd.t7 sky130_fd_pr__res_xhigh_po_1p41 l=2.66
X59 v9.t0 v8.t0 gnd.t17 sky130_fd_pr__res_xhigh_po_1p41 l=2.35
X60 v19.t1 v20.t1 gnd.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X61 v59.t0 v60.t1 gnd.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X62 v1.t1 v0.t0 gnd.t7 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X63 v45.t1 v46.t1 gnd.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X64 v51.t0 v50.t0 gnd.t10 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X65 v13.t1 v14.t0 gnd.t17 sky130_fd_pr__res_xhigh_po_1p41 l=1.84
X66 v51.t1 v52.t1 gnd.t10 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X67 v57.t0 v56.t1 gnd.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X68 v61.t0 v60.t0 gnd.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X69 v59.t1 v58.t0 gnd.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X70 v47.t1 v46.t0 gnd.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X71 v19.t0 v18.t1 gnd.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X72 v35.t1 v34.t1 gnd.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X73 gnd.t11 gnd.t12 gnd.t10 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X74 v39.t1 v38.t0 gnd.t0 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X75 gnd.t32 gnd.t33 gnd.t5 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X76 v25.t0 v26.t0 gnd.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X77 gnd.t20 gnd.t21 gnd.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X78 v33.t0 v34.t0 gnd.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X79 v61.t1 v62.t0 gnd.t4 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
R0 gnd.n30 gnd.n2 28676.6
R1 gnd.n32 gnd.n2 28676.6
R2 gnd.n30 gnd.n3 28673.3
R3 gnd.n32 gnd.n3 28673.3
R4 gnd.t17 gnd.t7 2422.51
R5 gnd.t3 gnd.t6 1972.93
R6 gnd.t6 gnd.t17 1942.12
R7 gnd.t0 gnd.t5 1879.36
R8 gnd.t10 gnd.t4 1838.28
R9 gnd.t5 gnd.t10 1749.27
R10 gnd.n31 gnd.t0 1582.68
R11 gnd.t7 gnd.n3 1480.72
R12 gnd.t4 gnd.n2 995.764
R13 gnd.n13 gnd.n12 461.243
R14 gnd.n22 gnd.n0 461.243
R15 gnd.n12 gnd.n11 459.111
R16 gnd.n41 gnd.n0 361.601
R17 gnd.n23 gnd.n22 235.98
R18 gnd.n31 gnd.t3 225.935
R19 gnd.n39 gnd.n38 207.393
R20 gnd.n35 gnd.n34 172.619
R21 gnd.n6 gnd.n5 171.554
R22 gnd.n10 gnd.n9 171.339
R23 gnd.n15 gnd.n14 171.339
R24 gnd.n19 gnd.n18 171.339
R25 gnd.n24 gnd.n23 171.339
R26 gnd.n28 gnd.n27 170.274
R27 gnd.n4 gnd.n1 151.714
R28 gnd.n17 gnd.n16 151.5
R29 gnd.n21 gnd.n20 151.5
R30 gnd.n26 gnd.n25 151.5
R31 gnd.n8 gnd.n7 150.434
R32 gnd.n41 gnd.n40 149.99
R33 gnd.n37 gnd.n36 142.754
R34 gnd.n40 gnd.n39 135.286
R35 gnd.n38 gnd.n37 128.887
R36 gnd.n25 gnd.n24 100.299
R37 gnd.n27 gnd.n26 96.0333
R38 gnd.n36 gnd.n35 84.94
R39 gnd.n20 gnd.n19 72.14
R40 gnd.n34 gnd.n33 70.499
R41 gnd.n7 gnd.n6 67.4467
R42 gnd.n29 gnd.n28 65.3297
R43 gnd.n5 gnd.n4 65.3133
R44 gnd.n16 gnd.n15 63.18
R45 gnd.n18 gnd.n17 61.0467
R46 gnd.n9 gnd.n8 58.9133
R47 gnd.n11 gnd.n10 58.9133
R48 gnd.n14 gnd.n13 54.6467
R49 gnd.n40 gnd.t16 39.3159
R50 gnd.n39 gnd.t15 39.3159
R51 gnd.n38 gnd.t35 39.3159
R52 gnd.n37 gnd.t34 39.3159
R53 gnd.n36 gnd.t31 39.3159
R54 gnd.n35 gnd.t30 39.3159
R55 gnd.n34 gnd.t21 39.3159
R56 gnd.n1 gnd.t20 39.3159
R57 gnd.n4 gnd.t39 39.3159
R58 gnd.n5 gnd.t38 39.3159
R59 gnd.n6 gnd.t25 39.3159
R60 gnd.n7 gnd.t24 39.3159
R61 gnd.n8 gnd.t27 39.3159
R62 gnd.n9 gnd.t26 39.3159
R63 gnd.n10 gnd.t19 39.3159
R64 gnd.n11 gnd.t18 39.3159
R65 gnd.n13 gnd.t36 39.3159
R66 gnd.n14 gnd.t37 39.3159
R67 gnd.n15 gnd.t11 39.3159
R68 gnd.n16 gnd.t12 39.3159
R69 gnd.n17 gnd.t32 39.3159
R70 gnd.n18 gnd.t33 39.3159
R71 gnd.n19 gnd.t1 39.3159
R72 gnd.n20 gnd.t2 39.3159
R73 gnd.n21 gnd.t28 39.3159
R74 gnd.n28 gnd.t29 39.3159
R75 gnd.n27 gnd.t13 39.3159
R76 gnd.n26 gnd.t14 39.3159
R77 gnd.n25 gnd.t22 39.3159
R78 gnd.n24 gnd.t23 39.3159
R79 gnd.n23 gnd.t8 39.3159
R80 gnd.n22 gnd.t9 39.3159
R81 gnd.n12 gnd.n2 13.296
R82 gnd.n3 gnd.n0 13.296
R83 gnd.n33 gnd.n1 10.1749
R84 gnd.n29 gnd.n21 8.94409
R85 gnd gnd.n41 6.4005
R86 gnd.n33 gnd.n32 2.9255
R87 gnd.n32 gnd.n31 2.9255
R88 gnd.n30 gnd.n29 2.9255
R89 gnd.n31 gnd.n30 2.9255
R90 v49.n0 v49.t1 10.6136
R91 v49.n0 v49.t0 10.5739
R92 v49 v49.n0 1.70606
R93 v50.n0 v50.t0 10.5296
R94 v50.n0 v50.t1 10.5285
R95 v50 v50.n0 2.5532
R96 v48.n0 v48.t1 13.5958
R97 v48.n0 v48.t0 10.612
R98 v48 v48.n0 1.67003
R99 v3.n0 v3.t1 10.5816
R100 v3.n0 v3.t0 10.5739
R101 v3 v3.n0 3.15304
R102 v4.n0 v4.t0 10.5339
R103 v4.n0 v4.t1 10.5285
R104 v4 v4.n0 3.88451
R105 v27.n0 v27.t1 10.6701
R106 v27.n0 v27.t0 10.5739
R107 v27 v27.n0 4.43205
R108 v28.n0 v28.t0 10.5296
R109 v28.n0 v28.t1 10.5285
R110 v28 v28.n0 3.80338
R111 v23.n0 v23.t1 10.6701
R112 v23.n0 v23.t0 10.5739
R113 v23 v23.n0 5.84121
R114 v22.n0 v22.t0 10.5296
R115 v22.n0 v22.t1 10.5285
R116 v22 v22.n0 5.21015
R117 v47.n0 v47.t1 10.5751
R118 v47.n0 v47.t0 10.5749
R119 v47 v47.n0 1.75448
R120 v55.n0 v55.t0 10.6701
R121 v55.n0 v55.t1 10.5739
R122 v55 v55.n0 5.83358
R123 v54.n0 v54.t0 10.6247
R124 v54.n0 v54.t1 10.5285
R125 v54 v54.n0 5.15858
R126 v33.n0 v33.t0 10.6155
R127 v33.n0 v33.t1 10.5739
R128 v33 v33.n0 1.70606
R129 v32.n0 v32.t1 13.6159
R130 v32.n0 v32.t0 10.612
R131 v32 v32.n0 1.67003
R132 v63.n0 v63.t1 10.5751
R133 v63.n0 v63.t0 10.5749
R134 v63 v63.n0 1.75448
R135 v62.n0 v62.t0 10.6247
R136 v62.n0 v62.t1 10.5285
R137 v62 v62.n0 2.53946
R138 v25.n0 v25.t1 10.6701
R139 v25.n0 v25.t0 10.5739
R140 v25 v25.n0 5.82165
R141 v24.n0 v24.t1 13.5018
R142 v24.n0 v24.t0 10.7924
R143 v24 v24.n0 6.39503
R144 v26.n0 v26.t1 10.5296
R145 v26.n0 v26.t0 10.5285
R146 v26 v26.n0 5.19298
R147 v17.n0 v17.t1 10.6701
R148 v17.n0 v17.t0 10.5739
R149 v17 v17.n0 1.70606
R150 v18.n0 v18.t1 10.5307
R151 v18.n0 v18.t0 10.5285
R152 v18 v18.n0 2.55213
R153 v37.n0 v37.t0 10.575
R154 v37.n0 v37.t1 10.5739
R155 v37 v37.n0 4.4858
R156 v36.n0 v36.t1 10.5296
R157 v36.n0 v36.t0 10.5285
R158 v36 v36.n0 3.82368
R159 v39.n0 v39.t0 10.575
R160 v39.n0 v39.t1 10.5739
R161 v39 v39.n0 5.88017
R162 v40.n0 v40.t0 13.4746
R163 v40.n0 v40.t1 10.7876
R164 v40 v40.n0 6.39503
R165 v64 v64.t0 12.2816
R166 v21.n0 v21.t0 10.6701
R167 v21.n0 v21.t1 10.5739
R168 v21 v21.n0 4.44684
R169 v20.n0 v20.t0 10.5309
R170 v20.n0 v20.t1 10.5285
R171 v20 v20.n0 3.8145
R172 v5.n0 v5.t0 10.5795
R173 v5.n0 v5.t1 10.5739
R174 v5 v5.n0 4.57149
R175 v6.n0 v6.t1 10.5328
R176 v6.n0 v6.t0 10.5285
R177 v6 v6.n0 5.29951
R178 v56.n0 v56.t1 13.4579
R179 v56.n0 v56.t0 10.7848
R180 v56 v56.n0 6.39503
R181 v9.n0 v9.t1 10.5773
R182 v9.n0 v9.t0 10.5739
R183 v9 v9.n0 5.84824
R184 v10.n0 v10.t1 10.5307
R185 v10.n0 v10.t0 10.5285
R186 v10 v10.n0 5.17712
R187 v29.n0 v29.t0 10.6701
R188 v29.n0 v29.t1 10.5739
R189 v29 v29.n0 3.21446
R190 v41.n0 v41.t1 10.575
R191 v41.n0 v41.t0 10.5739
R192 v41 v41.n0 5.87015
R193 v42.n0 v42.t1 10.5296
R194 v42.n0 v42.t0 10.5285
R195 v42 v42.n0 5.19536
R196 v16.n0 v16.t0 13.6693
R197 v16.n0 v16.t1 10.612
R198 v16 v16.n0 1.67003
R199 v57.n0 v57.t1 10.575
R200 v57.n0 v57.t0 10.5739
R201 v57 v57.n0 5.87254
R202 v58.n0 v58.t1 10.6247
R203 v58.n0 v58.t0 10.5285
R204 v58 v58.n0 5.15142
R205 v31.n0 v31.t1 10.6701
R206 v31.n0 v31.t0 10.5739
R207 v31 v31.n0 1.70606
R208 v30.n0 v30.t1 10.5296
R209 v30.n0 v30.t0 10.5285
R210 v30 v30.n0 2.57219
R211 v11.n0 v11.t0 10.5761
R212 v11.n0 v11.t1 10.5739
R213 v11 v11.n0 4.51275
R214 v12.n0 v12.t0 10.5307
R215 v12.n0 v12.t1 10.5285
R216 v12 v12.n0 3.84069
R217 v53.n0 v53.t1 10.6701
R218 v53.n0 v53.t0 10.5739
R219 v53 v53.n0 4.44159
R220 v52.n0 v52.t0 10.5296
R221 v52.n0 v52.t1 10.5285
R222 v52 v52.n0 3.81054
R223 v15.n0 v15.t0 10.6713
R224 v15.n0 v15.t1 10.5739
R225 v15 v15.n0 1.70653
R226 v13.n0 v13.t1 10.575
R227 v13.n0 v13.t0 10.5739
R228 v13 v13.n0 3.27356
R229 v1.n0 v1.t0 10.5871
R230 v1.n0 v1.t1 10.5739
R231 v1 v1.n0 1.91746
R232 v2.n0 v2.t1 10.5394
R233 v2.n0 v2.t0 10.5285
R234 v2 v2.n0 2.45788
R235 v43.n0 v43.t1 10.575
R236 v43.n0 v43.t0 10.5739
R237 v43 v43.n0 4.48055
R238 v14.n0 v14.t1 10.5309
R239 v14.n0 v14.t0 10.5285
R240 v14 v14.n0 2.58212
R241 v45.n0 v45.t0 10.6671
R242 v45.n0 v45.t1 10.5769
R243 v45 v45.n0 3.21745
R244 v44.n0 v44.t1 10.5296
R245 v44.n0 v44.t0 10.5285
R246 v44 v44.n0 3.80338
R247 v38.n0 v38.t0 10.5296
R248 v38.n0 v38.t1 10.5285
R249 v38 v38.n0 5.203
R250 v35.n0 v35.t0 10.5752
R251 v35.n0 v35.t1 10.5739
R252 v35 v35.n0 3.21923
R253 v7.n0 v7.t1 10.5773
R254 v7.n0 v7.t0 10.5739
R255 v7 v7.n0 5.98279
R256 v8.n0 v8.t0 13.5844
R257 v8.n0 v8.t1 10.8954
R258 v8 v8.n0 6.39217
R259 v19.n0 v19.t1 10.6701
R260 v19.n0 v19.t0 10.5739
R261 v19 v19.n0 3.18426
R262 v59.n0 v59.t1 10.6701
R263 v59.n0 v59.t0 10.5739
R264 v59 v59.n0 4.43682
R265 v60.n0 v60.t1 10.6247
R266 v60.n0 v60.t0 10.5285
R267 v60 v60.n0 3.75944
R268 v0 v0.t0 12.7924
R269 v46.n0 v46.t1 10.6247
R270 v46.n0 v46.t0 10.5285
R271 v46 v46.n0 2.53946
R272 v51.n0 v51.t0 10.575
R273 v51.n0 v51.t1 10.5739
R274 v51 v51.n0 3.22926
R275 v61.n0 v61.t0 10.6701
R276 v61.n0 v61.t1 10.5739
R277 v61 v61.n0 3.20325
R278 v34.n0 v34.t1 10.6247
R279 v34.n0 v34.t0 10.5285
R280 v34 v34.n0 2.52825
C0 v10 v21 0.02605f
C1 v44 v48 0.12056f
C2 v13 v4 0.01814f
C3 v0 v4 0.01508f
C4 v48 v53 0.12271f
C5 v59 v58 0.13601f
C6 v18 v16 0.73858f
C7 v1 v0 0.60526f
C8 v8 v23 0.05167f
C9 v46 v51 0.02493f
C10 v36 v34 1.36923f
C11 v20 v19 0.0646f
C12 v50 v48 0.73678f
C13 v63 v64 0.1865f
C14 v17 v18 0.0917f
C15 v58 v64 0.15411f
C16 v4 v2 1.32227f
C17 v18 v31 0.02179f
C18 v59 v57 1.89898f
C19 v19 v12 0.02564f
C20 v59 v56 0.01311f
C21 v28 v37 0.0251f
C22 v1 v2 0.02376f
C23 v47 v32 0.02425f
C24 v59 v54 0.02147f
C25 v0 v7 0.15367f
C26 v9 v10 0.04456f
C27 v32 v37 0.12272f
C28 v13 v2 0.01887f
C29 v44 v53 0.02514f
C30 v0 v2 1.16018f
C31 v40 v39 0.10723f
C32 v24 v25 2.49563f
C33 v4 v6 1.6918f
C34 v50 v49 0.15573f
C35 v50 v63 0.02163f
C36 v62 v64 1.21931f
C37 v35 v37 1.55046f
C38 v45 v46 0.11369f
C39 v62 v63 0.13703f
C40 v20 v16 0.01378f
C41 v57 v58 0.13595f
C42 v36 v43 0.02159f
C43 v19 v21 1.54419f
C44 v56 v58 0.55116f
C45 v52 v48 0.01369f
C46 v59 v61 1.55555f
C47 v30 v31 0.08794f
C48 v15 v16 0.08905f
C49 v20 v27 0.02143f
C50 v22 v23 0.07152f
C51 v21 v23 1.89384f
C52 v24 v22 2.07533f
C53 v32 v39 0.11987f
C54 v16 v12 0.12063f
C55 v53 v54 0.1272f
C56 v8 v11 0.01311f
C57 v47 v45 1.27985f
C58 v38 v37 0.09637f
C59 v25 v26 0.07716f
C60 v5 v3 1.51072f
C61 v59 v52 0.02147f
C62 v48 v51 0.13156f
C63 v56 v57 2.5376f
C64 v61 v63 1.27985f
C65 v14 v15 0.05614f
C66 v28 v26 1.71746f
C67 v25 v27 1.89543f
C68 v57 v54 0.02147f
C69 v14 v12 1.37455f
C70 v48 v55 0.11987f
C71 v36 v32 0.01377f
C72 v56 v54 2.07551f
C73 v27 v28 0.08057f
C74 v7 v6 0.03657f
C75 v10 v23 1.58849f
C76 v9 v6 0.01724f
C77 v32 v26 0.12029f
C78 v44 v43 0.10714f
C79 v21 v16 0.12277f
C80 v47 v46 0.11373f
C81 v36 v35 0.09669f
C82 v33 v34 0.12582f
C83 v20 v18 1.36887f
C84 v11 v12 0.04901f
C85 v38 v39 0.10121f
C86 v42 v48 0.1203f
C87 v32 v31 0.12374f
C88 v5 v4 0.03159f
C89 v27 v22 0.02143f
C90 v29 v27 1.5529f
C91 v52 v53 0.12756f
C92 v49 v51 1.2717f
C93 v50 v61 0.02147f
C94 v29 v31 1.27963f
C95 v61 v62 0.137f
C96 v10 v16 0.1203f
C97 v36 v38 1.71154f
C98 v44 v51 0.02514f
C99 v36 v45 0.02159f
C100 v53 v51 1.55159f
C101 v50 v52 1.36553f
C102 v0 v5 0.1233f
C103 v11 v4 0.0178f
C104 v60 v59 0.13643f
C105 v13 v14 0.05301f
C106 v55 v53 1.89779f
C107 v52 v54 1.71504f
C108 v30 v33 0.02514f
C109 v32 v34 0.73825f
C110 v29 v18 0.02163f
C111 v48 v46 1.21914f
C112 v50 v51 0.12805f
C113 v13 v11 1.55225f
C114 v60 v64 0.12057f
C115 v11 v10 0.04656f
C116 v44 v42 1.71627f
C117 v35 v34 0.09194f
C118 v5 v7 1.87971f
C119 v42 v53 0.02493f
C120 v56 v55 0.12772f
C121 v40 v43 0.01313f
C122 v39 v37 1.89634f
C123 v60 v58 1.71687f
C124 v61 v52 0.02163f
C125 v55 v54 0.1272f
C126 v44 v45 0.11317f
C127 v47 v48 0.1586f
C128 v30 v28 1.37467f
C129 v24 v23 0.07226f
C130 v41 v43 1.89463f
C131 v9 v11 1.89368f
C132 v30 v32 1.22402f
C133 v32 v33 0.68843f
C134 v36 v37 0.10155f
C135 v49 v46 0.02514f
C136 v24 v39 0.04779f
C137 v45 v34 0.02179f
C138 v5 v6 0.03415f
C139 v40 v41 2.51611f
C140 v26 v37 0.02532f
C141 v19 v16 0.13162f
C142 v29 v30 0.08433f
C143 v30 v35 0.02537f
C144 v35 v33 1.28018f
C145 v60 v62 1.37506f
C146 v20 v22 1.71403f
C147 v44 v46 1.37506f
C148 v20 v21 0.06935f
C149 v20 v29 0.02163f
C150 v52 v51 0.11996f
C151 v16 v23 0.11987f
C152 v40 v55 0.04831f
C153 v17 v19 1.27804f
C154 v19 v14 0.02541f
C155 v8 v10 0.5416f
C156 v24 v26 0.55405f
C157 v11 v6 0.01745f
C158 v42 v43 0.11271f
C159 v32 v28 0.12053f
C160 v3 v4 0.02937f
C161 v21 v12 0.02559f
C162 v39 v26 1.58219f
C163 v25 v22 0.02143f
C164 v24 v27 0.0131f
C165 v40 v42 0.5513f
C166 v60 v61 0.13646f
C167 v29 v28 0.08388f
C168 v38 v43 0.02159f
C169 v35 v28 0.0251f
C170 v1 v3 1.17004f
C171 v45 v43 1.55772f
C172 v47 v34 0.02179f
C173 v8 v7 0.03886f
C174 v9 v8 2.45916f
C175 v40 v38 2.07259f
C176 v13 v15 1.26142f
C177 v0 v15 0.02431f
C178 v42 v41 0.10671f
C179 v0 v3 0.13391f
C180 v35 v32 0.13136f
C181 v13 v12 0.05141f
C182 v10 v12 1.70992f
C183 v18 v19 0.06489f
C184 v21 v22 0.06911f
C185 v17 v16 0.66585f
C186 v14 v16 1.21926f
C187 v38 v41 0.02159f
C188 v27 v26 0.08021f
C189 v16 v31 0.0245f
C190 v42 v55 1.58135f
C191 v49 v48 0.70728f
C192 v48 v63 0.02425f
C193 v8 v6 2.07017f
C194 v17 v14 0.02537f
C195 v15 v2 0.01992f
C196 v3 v2 0.0268f
C197 v56 gnd 2.40728f
C198 v40 gnd 2.38733f
C199 v24 gnd 2.43442f
C200 v8 gnd 2.65358f
C201 v57 gnd 1.39148f
C202 v55 gnd 1.19815f
C203 v41 gnd 1.4031f
C204 v39 gnd 1.21716f
C205 v25 gnd 1.41361f
C206 v23 gnd 1.2439f
C207 v9 gnd 1.4726f
C208 v7 gnd 2.14783f
C209 v58 gnd 1.38404f
C210 v54 gnd 0.87085f
C211 v42 gnd 0.72721f
C212 v38 gnd 0.89685f
C213 v26 gnd 0.74725f
C214 v22 gnd 0.92937f
C215 v10 gnd 0.78548f
C216 v6 gnd 1.11471f
C217 v59 gnd 0.62935f
C218 v53 gnd 0.63067f
C219 v43 gnd 0.64688f
C220 v37 gnd 0.65203f
C221 v27 gnd 0.66618f
C222 v21 gnd 0.68556f
C223 v11 gnd 0.72239f
C224 v5 gnd 0.90863f
C225 v60 gnd 0.63372f
C226 v52 gnd 0.6245f
C227 v44 gnd 0.61524f
C228 v36 gnd 0.64138f
C229 v28 gnd 0.63761f
C230 v20 gnd 0.67978f
C231 v12 gnd 0.67997f
C232 v4 gnd 0.86121f
C233 v61 gnd 0.54421f
C234 v51 gnd 0.55425f
C235 v45 gnd 0.55722f
C236 v35 gnd 0.57001f
C237 v29 gnd 0.58306f
C238 v19 gnd 0.60577f
C239 v13 gnd 0.63366f
C240 v3 gnd 0.82192f
C241 v62 gnd 0.5485f
C242 v50 gnd 0.69419f
C243 v46 gnd 0.53164f
C244 v34 gnd 0.71027f
C245 v30 gnd 0.55486f
C246 v18 gnd 0.75344f
C247 v14 gnd 0.59918f
C248 v2 gnd 0.78256f
C249 v64 gnd 1.09738f
C250 v63 gnd 1.07065f
C251 v49 gnd 1.08211f
C252 v48 gnd 1.82764f
C253 v47 gnd 1.08423f
C254 v33 gnd 1.09674f
C255 v32 gnd 1.87488f
C256 v31 gnd 1.10867f
C257 v17 gnd 1.13778f
C258 v16 gnd 1.97001f
C259 v15 gnd 1.15716f
C260 v0 gnd 1.74573f
C261 v1 gnd 1.3571f
C262 v8.t0 gnd 0.49372f
C263 v8.t1 gnd 0.16832f
C264 v8.n0 gnd 3.64859f
C265 v38.t0 gnd 0.09206f
C266 v38.t1 gnd 0.09199f
C267 v38.n0 gnd 1.74551f
C268 v57.t1 gnd 0.10808f
C269 v57.t0 gnd 0.10799f
C270 v57.n0 gnd 2.06002f
C271 v41.t1 gnd 0.10823f
C272 v41.t0 gnd 0.10814f
C273 v41.n0 gnd 2.0596f
C274 v9.t1 gnd 0.11106f
C275 v9.t0 gnd 0.11079f
C276 v9.n0 gnd 2.05043f
C277 v56.t0 gnd 0.16999f
C278 v56.t1 gnd 0.50347f
C279 v56.n0 gnd 3.60881f
C280 v6.t1 gnd 0.08835f
C281 v6.t0 gnd 0.08808f
C282 v6.n0 gnd 1.7531f
C283 v40.t1 gnd 0.16901f
C284 v40.t0 gnd 0.50442f
C285 v40.n0 gnd 3.61131f
C286 v24.t0 gnd 0.16742f
C287 v24.t1 gnd 0.50594f
C288 v24.n0 gnd 3.61546f
C289 v25.t0 gnd 0.10781f
C290 v25.t1 gnd 0.11542f
C291 v25.n0 gnd 2.05772f
C292 v54.t1 gnd 0.09161f
C293 v54.t0 gnd 0.09812f
C294 v54.n0 gnd 1.74436f
C295 v22.t0 gnd 0.09168f
C296 v22.t1 gnd 0.09161f
C297 v22.n0 gnd 1.74647f
.ends

