magic
tech sky130A
magscale 1 2
timestamp 1749289931
<< metal1 >>
rect 9957 -17093 10017 -15149
rect 10045 -16445 10105 -15149
rect 10133 -15797 10193 -15149
rect 10133 -16383 10206 -15797
rect 10045 -17031 10180 -16445
rect 9957 -17679 10139 -17093
<< end >>
