magic
tech sky130A
magscale 1 2
timestamp 1750079478
<< error_s >>
rect 1533 1475 1539 1481
rect 1587 1475 1593 1481
rect 1651 1475 1657 1481
rect 1705 1475 1711 1481
rect 3037 1475 3043 1481
rect 3091 1475 3097 1481
rect 3155 1475 3161 1481
rect 3209 1475 3215 1481
rect 1527 1469 1533 1475
rect 1593 1469 1599 1475
rect 1645 1469 1651 1475
rect 1711 1469 1717 1475
rect 3031 1469 3037 1475
rect 3097 1469 3103 1475
rect 3149 1469 3155 1475
rect 3215 1469 3221 1475
rect 1527 1415 1533 1421
rect 1593 1415 1599 1421
rect 1645 1415 1651 1421
rect 1711 1415 1717 1421
rect 3031 1415 3037 1421
rect 3097 1415 3103 1421
rect 3149 1415 3155 1421
rect 3215 1415 3221 1421
rect 1533 1409 1539 1415
rect 1587 1409 1593 1415
rect 1651 1409 1657 1415
rect 1705 1409 1711 1415
rect 3037 1409 3043 1415
rect 3091 1409 3097 1415
rect 3155 1409 3161 1415
rect 3209 1409 3215 1415
rect 781 1387 787 1393
rect 835 1387 841 1393
rect 899 1387 905 1393
rect 953 1387 959 1393
rect 2285 1387 2291 1393
rect 2339 1387 2345 1393
rect 2403 1387 2409 1393
rect 2457 1387 2463 1393
rect 775 1381 781 1387
rect 841 1381 847 1387
rect 893 1381 899 1387
rect 959 1381 965 1387
rect 2279 1381 2285 1387
rect 2345 1381 2351 1387
rect 2397 1381 2403 1387
rect 2463 1381 2469 1387
rect 775 1327 781 1333
rect 841 1327 847 1333
rect 893 1327 899 1333
rect 959 1327 965 1333
rect 2279 1327 2285 1333
rect 2345 1327 2351 1333
rect 2397 1327 2403 1333
rect 2463 1327 2469 1333
rect 781 1321 787 1327
rect 835 1321 841 1327
rect 899 1321 905 1327
rect 953 1321 959 1327
rect 2285 1321 2291 1327
rect 2339 1321 2345 1327
rect 2403 1321 2409 1327
rect 2457 1321 2463 1327
rect 1275 1299 1281 1305
rect 1329 1299 1335 1305
rect 1909 1299 1915 1305
rect 1963 1299 1969 1305
rect 2779 1299 2785 1305
rect 2833 1299 2839 1305
rect 3413 1299 3419 1305
rect 3467 1299 3473 1305
rect 1269 1293 1275 1299
rect 1335 1293 1341 1299
rect 1903 1293 1909 1299
rect 1969 1293 1975 1299
rect 2773 1293 2779 1299
rect 2839 1293 2845 1299
rect 3407 1293 3413 1299
rect 3473 1293 3479 1299
rect 1269 1239 1275 1245
rect 1335 1239 1341 1245
rect 1903 1239 1909 1245
rect 1969 1239 1975 1245
rect 2773 1239 2779 1245
rect 2839 1239 2845 1245
rect 3407 1239 3413 1245
rect 3473 1239 3479 1245
rect 1275 1233 1281 1239
rect 1329 1233 1335 1239
rect 1909 1233 1915 1239
rect 1963 1233 1969 1239
rect 2779 1233 2785 1239
rect 2833 1233 2839 1239
rect 3413 1233 3419 1239
rect 3467 1233 3473 1239
rect 523 1211 529 1217
rect 577 1211 583 1217
rect 1157 1211 1163 1217
rect 1211 1211 1217 1217
rect 2027 1211 2033 1217
rect 2081 1211 2087 1217
rect 2661 1211 2667 1217
rect 2715 1211 2721 1217
rect 517 1205 523 1211
rect 583 1205 589 1211
rect 1151 1205 1157 1211
rect 1217 1205 1223 1211
rect 2021 1205 2027 1211
rect 2087 1205 2093 1211
rect 2655 1205 2661 1211
rect 2721 1205 2727 1211
rect 517 1151 523 1157
rect 583 1151 589 1157
rect 1151 1151 1157 1157
rect 1217 1151 1223 1157
rect 2021 1151 2027 1157
rect 2087 1151 2093 1157
rect 2655 1151 2661 1157
rect 2721 1151 2727 1157
rect 523 1145 529 1151
rect 577 1145 583 1151
rect 1157 1145 1163 1151
rect 1211 1145 1217 1151
rect 2027 1145 2033 1151
rect 2081 1145 2087 1151
rect 2661 1145 2667 1151
rect 2715 1145 2721 1151
rect 2490 1035 2496 1041
rect 2544 1035 2550 1041
rect 2950 1035 2956 1041
rect 3004 1035 3010 1041
rect 2484 1029 2490 1035
rect 2550 1029 2556 1035
rect 2944 1029 2950 1035
rect 3010 1029 3016 1035
rect 2484 975 2490 981
rect 2550 975 2556 981
rect 2944 975 2950 981
rect 3010 975 3016 981
rect 2490 969 2496 975
rect 2544 969 2550 975
rect 2950 969 2956 975
rect 3004 969 3010 975
rect 2574 947 2580 953
rect 2628 947 2634 953
rect 2866 947 2872 953
rect 2920 947 2926 953
rect 2568 941 2574 947
rect 2634 941 2640 947
rect 2860 941 2866 947
rect 2926 941 2932 947
rect 2568 887 2574 893
rect 2634 887 2640 893
rect 2860 887 2866 893
rect 2926 887 2932 893
rect 2574 881 2580 887
rect 2628 881 2634 887
rect 2866 881 2872 887
rect 2920 881 2926 887
rect 1908 859 1914 865
rect 1962 859 1968 865
rect 2026 859 2032 865
rect 2080 859 2086 865
rect 1902 853 1908 859
rect 1968 853 1974 859
rect 2020 853 2026 859
rect 2086 853 2092 859
rect 1902 799 1908 805
rect 1968 799 1974 805
rect 2020 799 2026 805
rect 2086 799 2092 805
rect 1908 793 1914 799
rect 1962 793 1968 799
rect 2026 793 2032 799
rect 2080 793 2086 799
rect 1157 771 1163 777
rect 1211 771 1217 777
rect 1275 771 1281 777
rect 1329 771 1335 777
rect 1151 765 1157 771
rect 1217 765 1223 771
rect 1269 765 1275 771
rect 1335 765 1341 771
rect 1151 711 1157 717
rect 1217 711 1223 717
rect 1269 711 1275 717
rect 1335 711 1341 717
rect 1157 705 1163 711
rect 1211 705 1217 711
rect 1275 705 1281 711
rect 1329 705 1335 711
rect 1651 683 1657 689
rect 1705 683 1711 689
rect 2285 683 2291 689
rect 2339 683 2345 689
rect 1645 677 1651 683
rect 1711 677 1717 683
rect 2279 677 2285 683
rect 2345 677 2351 683
rect 1645 623 1651 629
rect 1711 623 1717 629
rect 2279 623 2285 629
rect 2345 623 2351 629
rect 1651 617 1657 623
rect 1705 617 1711 623
rect 2285 617 2291 623
rect 2339 617 2345 623
rect 899 595 905 601
rect 953 595 959 601
rect 1533 595 1539 601
rect 1587 595 1593 601
rect 893 589 899 595
rect 959 589 965 595
rect 1527 589 1533 595
rect 1593 589 1599 595
rect 893 535 899 541
rect 959 535 965 541
rect 1527 535 1533 541
rect 1593 535 1599 541
rect 899 529 905 535
rect 953 529 959 535
rect 1533 529 1539 535
rect 1587 529 1593 535
rect 3155 419 3161 425
rect 3209 419 3215 425
rect 3149 413 3155 419
rect 3215 413 3221 419
rect 3149 359 3155 365
rect 3215 359 3221 365
rect 3155 353 3161 359
rect 3209 353 3215 359
rect 3413 243 3419 249
rect 3467 243 3473 249
rect 3407 237 3413 243
rect 3473 237 3479 243
rect 3407 183 3413 189
rect 3473 183 3479 189
rect 3413 177 3419 183
rect 3467 177 3473 183
<< metal1 >>
rect 1527 1415 1533 1475
rect 1593 1415 1599 1475
rect 1645 1415 1651 1475
rect 1711 1415 1717 1475
rect 3031 1415 3037 1475
rect 3097 1415 3103 1475
rect 3149 1415 3155 1475
rect 3215 1415 3221 1475
rect 775 1327 781 1387
rect 841 1327 847 1387
rect 893 1327 899 1387
rect 959 1327 965 1387
rect 517 1151 523 1211
rect 583 1151 589 1211
rect 530 1033 576 1151
rect 788 925 834 1327
rect 906 925 952 1327
rect 1269 1239 1275 1299
rect 1335 1239 1341 1299
rect 1151 1151 1157 1211
rect 1217 1151 1223 1211
rect 1164 1033 1210 1151
rect 1282 1033 1328 1239
rect 1540 925 1586 1415
rect 1658 925 1704 1415
rect 2279 1327 2285 1387
rect 2345 1327 2351 1387
rect 2397 1327 2403 1387
rect 2463 1327 2469 1387
rect 1903 1239 1909 1299
rect 1969 1239 1975 1299
rect 1916 1033 1962 1239
rect 2021 1151 2027 1211
rect 2087 1151 2093 1211
rect 2034 1033 2080 1151
rect 2292 925 2338 1327
rect 2410 925 2456 1327
rect 2773 1239 2779 1299
rect 2839 1239 2845 1299
rect 2655 1151 2661 1211
rect 2721 1151 2727 1211
rect 2484 975 2490 1035
rect 2550 975 2556 1035
rect 2668 1033 2714 1151
rect 2786 1033 2832 1239
rect 2944 975 2950 1035
rect 3010 975 3016 1035
rect 1902 799 1908 859
rect 1968 799 1974 859
rect 2020 799 2026 859
rect 2086 799 2092 859
rect 1151 711 1157 771
rect 1217 711 1223 771
rect 1269 711 1275 771
rect 1335 711 1341 771
rect 1164 645 1210 711
rect 893 535 899 595
rect 959 535 965 595
rect 1282 525 1328 711
rect 1645 623 1651 683
rect 1711 623 1717 683
rect 1916 645 1962 799
rect 1527 535 1533 595
rect 1593 535 1599 595
rect 2034 525 2080 799
rect 2279 623 2285 683
rect 2345 623 2351 683
rect 2484 645 2530 975
rect 2568 887 2574 947
rect 2634 887 2640 947
rect 2410 633 2530 645
rect 2449 599 2530 633
rect 2594 645 2640 887
rect 2860 887 2866 947
rect 2926 887 2932 947
rect 2860 645 2906 887
rect 2594 599 2675 645
rect 2832 599 2906 645
rect 2970 645 3016 975
rect 3044 925 3090 1415
rect 3162 925 3208 1415
rect 3407 1239 3413 1299
rect 3473 1239 3479 1299
rect 3420 1033 3466 1239
rect 2970 599 3051 645
rect 3162 419 3208 525
rect 3149 359 3155 419
rect 3215 359 3221 419
rect 3420 243 3466 535
rect 3407 183 3413 243
rect 3473 183 3479 243
<< via1 >>
rect 1533 1415 1593 1475
rect 1651 1415 1711 1475
rect 3037 1415 3097 1475
rect 3155 1415 3215 1475
rect 781 1327 841 1387
rect 899 1327 959 1387
rect 523 1151 583 1211
rect 1275 1239 1335 1299
rect 1157 1151 1217 1211
rect 2285 1327 2345 1387
rect 2403 1327 2463 1387
rect 1909 1239 1969 1299
rect 2027 1151 2087 1211
rect 2779 1239 2839 1299
rect 2661 1151 2721 1211
rect 2490 975 2550 1035
rect 2950 975 3010 1035
rect 1908 799 1968 859
rect 2026 799 2086 859
rect 1157 711 1217 771
rect 1275 711 1335 771
rect 899 535 959 595
rect 1651 623 1711 683
rect 1533 535 1593 595
rect 2285 623 2345 683
rect 2574 887 2634 947
rect 2866 887 2926 947
rect 3413 1239 3473 1299
rect 3155 359 3215 419
rect 3413 183 3473 243
use cm_ncell2_cell  cm_ncell2_cell_0
timestamp 1750079478
transform -1 0 3498 0 1 -5
box -4 -8 3506 1588
<< end >>
