magic
tech sky130A
magscale 1 2
timestamp 1749548291
<< error_s >>
rect 1074 684 1080 690
rect 1128 684 1134 690
rect 1068 678 1074 684
rect 1134 678 1140 684
rect 1068 624 1074 630
rect 1134 624 1140 630
rect 1074 618 1080 624
rect 1128 618 1134 624
rect 798 596 804 602
rect 852 596 858 602
rect 792 590 798 596
rect 858 590 864 596
rect 792 536 798 542
rect 858 536 864 542
rect 798 530 804 536
rect 852 530 858 536
rect 522 508 528 514
rect 576 508 582 514
rect 516 502 522 508
rect 582 502 588 508
rect 516 448 522 454
rect 582 448 588 454
rect 522 442 528 448
rect 576 442 582 448
rect 246 420 252 426
rect 300 420 306 426
rect 240 414 246 420
rect 306 414 312 420
rect 240 360 246 366
rect 306 360 312 366
rect 246 354 252 360
rect 300 354 306 360
rect 891 -397 897 -391
rect 945 -397 951 -391
rect 885 -403 891 -397
rect 951 -403 957 -397
rect 885 -457 891 -451
rect 951 -457 957 -451
rect 891 -463 897 -457
rect 945 -463 951 -457
rect 615 -485 621 -479
rect 669 -485 675 -479
rect 609 -491 615 -485
rect 675 -491 681 -485
rect 609 -545 615 -539
rect 675 -545 681 -539
rect 615 -551 621 -545
rect 669 -551 675 -545
rect 339 -573 345 -567
rect 393 -573 399 -567
rect 333 -579 339 -573
rect 399 -579 405 -573
rect 333 -633 339 -627
rect 399 -633 405 -627
rect 339 -639 345 -633
rect 393 -639 399 -633
rect 63 -661 69 -655
rect 117 -661 123 -655
rect 57 -667 63 -661
rect 123 -667 129 -661
rect 57 -721 63 -715
rect 123 -721 129 -715
rect 63 -727 69 -721
rect 117 -727 123 -721
<< metal1 >>
rect 1074 684 1134 690
rect 798 596 858 602
rect 522 508 582 514
rect 246 420 306 426
rect 246 70 306 360
rect 522 70 582 448
rect 63 -661 123 70
rect 339 -573 399 70
rect 615 -485 675 71
rect 798 70 858 536
rect 1074 70 1134 624
rect 891 -397 951 70
rect 891 -463 951 -457
rect 615 -551 675 -545
rect 339 -639 399 -633
rect 63 -727 123 -721
<< via1 >>
rect 1074 624 1134 684
rect 798 536 858 596
rect 522 448 582 508
rect 246 360 306 420
rect 891 -457 951 -397
rect 615 -545 675 -485
rect 339 -633 399 -573
rect 63 -721 123 -661
use hnmos_4  hnmos_4_0
timestamp 1749548291
transform 1 0 42 0 1 44
box -8 0 1096 198
<< end >>
