.subckt rseg_2_v3 v0 v1 v2 v3 v4 v5 v6 v7 v8 v9 v10 v11 v12 v13 v14 v15 v16 v17 v18 v19 v20 v21 v22 v23 v24 v25 v26 v27 v28 v29 v30 v31 v32 v33 v34 v35 v36 v37 v38 v39 v40 v41 v42 v43 v44 v45 v46 v47 v48 gnd
XR1 v0 v1 gnd sky130_fd_pr__res_xhigh_po_0p35 L=2.0389 mult=1 m=1
XR2 v1 v2 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.7967 mult=1 m=1
XR3 v2 v3 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.6105 mult=1 m=1
XR4 v3 v4 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.4802 mult=1 m=1
XR5 v4 v5 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.3684 mult=1 m=1
XR6 v5 v6 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.2845 mult=1 m=1
XR7 v6 v7 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.2101 mult=1 m=1
XR8 v7 v8 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.1449 mult=1 m=1
XR9 v8 v9 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.0890 mult=1 m=1
XR10 v9 v10 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.0518 mult=1 m=1
XR11 v10 v11 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.0146 mult=1 m=1
XR12 v11 v12 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.0066 mult=1 m=1
XR13 v12 v13 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.9294 mult=1 m=1
XR14 v13 v14 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.8927 mult=1 m=1
XR15 v14 v15 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.8376 mult=1 m=1
XR16 v15 v16 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.7826 mult=1 m=1
XR17 v16 v17 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.7642 mult=1 m=1
XR18 v17 v18 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.7459 mult=1 m=1
XR19 v18 v19 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.7091 mult=1 m=1
XR20 v19 v20 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6724 mult=1 m=1
XR21 v20 v21 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6724 mult=1 m=1
XR22 v21 v22 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6540 mult=1 m=1
XR23 v22 v23 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6357 mult=1 m=1
XR24 v23 v24 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6173 mult=1 m=1
XR25 v24 v25 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6173 mult=1 m=1
XR26 v25 v26 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6173 mult=1 m=1
XR27 v26 v27 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.5989 mult=1 m=1
XR28 v27 v28 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6173 mult=1 m=1
XR29 v28 v29 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.5989 mult=1 m=1
XR30 v29 v30 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.5989 mult=1 m=1
XR31 v30 v31 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6173 mult=1 m=1
XR32 v31 v32 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6173 mult=1 m=1
XR33 v32 v33 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6357 mult=1 m=1
XR34 v33 v34 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6357 mult=1 m=1
XR35 v34 v35 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6540 mult=1 m=1
XR36 v35 v36 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6724 mult=1 m=1
XR37 v36 v37 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.6907 mult=1 m=1
XR38 v37 v38 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.7275 mult=1 m=1
XR39 v38 v39 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.7275 mult=1 m=1
XR40 v39 v40 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.7826 mult=1 m=1
XR41 v40 v41 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.8009 mult=1 m=1
XR42 v41 v42 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.8376 mult=1 m=1
XR43 v42 v43 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.8927 mult=1 m=1
XR44 v43 v44 gnd sky130_fd_pr__res_xhigh_po_0p69 L=1.9294 mult=1 m=1
XR45 v44 v45 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.0066 mult=1 m=1
XR46 v45 v46 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.0052 mult=1 m=1
XR47 v46 v47 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.0424 mult=1 m=1
XR48 v47 v48 gnd sky130_fd_pr__res_xhigh_po_0p35 L=1.0890 mult=1 m=1
.ends