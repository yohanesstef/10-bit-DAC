.model dac_buff dac_bridge(out_low=0 out_high=1.8
  +out_undef=0.9 input_load=10e-15 t_rise=100e-9 t_fall=100e-9)
  
.model adc_buff adc_bridge(in_low=0 in_high=1.8)