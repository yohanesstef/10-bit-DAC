magic
tech sky130A
magscale 1 2
timestamp 1749382774
<< metal1 >>
rect 2907 3395 2967 3401
rect 2907 2955 2967 3335
rect 3083 3307 3143 3313
rect 2995 3219 3055 3225
rect 2995 2955 3055 3159
rect 3083 2955 3143 3247
<< via1 >>
rect 2907 3335 2967 3395
rect 3083 3247 3143 3307
rect 2995 3159 3055 3219
<< metal2 >>
rect 2721 3335 2907 3395
rect 2967 3335 2973 3395
rect 2721 3247 3083 3307
rect 3143 3247 3149 3307
rect 2721 3159 2995 3219
rect 3055 3159 3061 3219
<< end >>
