magic
tech sky130A
magscale 1 2
timestamp 1750134470
<< metal3 >>
rect -2916 2372 -2144 2400
rect -2916 1948 -2228 2372
rect -2164 1948 -2144 2372
rect -2916 1920 -2144 1948
rect -1904 2372 -1132 2400
rect -1904 1948 -1216 2372
rect -1152 1948 -1132 2372
rect -1904 1920 -1132 1948
rect -892 2372 -120 2400
rect -892 1948 -204 2372
rect -140 1948 -120 2372
rect -892 1920 -120 1948
rect 120 2372 892 2400
rect 120 1948 808 2372
rect 872 1948 892 2372
rect 120 1920 892 1948
rect 1132 2372 1904 2400
rect 1132 1948 1820 2372
rect 1884 1948 1904 2372
rect 1132 1920 1904 1948
rect 2144 2372 2916 2400
rect 2144 1948 2832 2372
rect 2896 1948 2916 2372
rect 2144 1920 2916 1948
rect -2916 1652 -2144 1680
rect -2916 1228 -2228 1652
rect -2164 1228 -2144 1652
rect -2916 1200 -2144 1228
rect -1904 1652 -1132 1680
rect -1904 1228 -1216 1652
rect -1152 1228 -1132 1652
rect -1904 1200 -1132 1228
rect -892 1652 -120 1680
rect -892 1228 -204 1652
rect -140 1228 -120 1652
rect -892 1200 -120 1228
rect 120 1652 892 1680
rect 120 1228 808 1652
rect 872 1228 892 1652
rect 120 1200 892 1228
rect 1132 1652 1904 1680
rect 1132 1228 1820 1652
rect 1884 1228 1904 1652
rect 1132 1200 1904 1228
rect 2144 1652 2916 1680
rect 2144 1228 2832 1652
rect 2896 1228 2916 1652
rect 2144 1200 2916 1228
rect -2916 932 -2144 960
rect -2916 508 -2228 932
rect -2164 508 -2144 932
rect -2916 480 -2144 508
rect -1904 932 -1132 960
rect -1904 508 -1216 932
rect -1152 508 -1132 932
rect -1904 480 -1132 508
rect -892 932 -120 960
rect -892 508 -204 932
rect -140 508 -120 932
rect -892 480 -120 508
rect 120 932 892 960
rect 120 508 808 932
rect 872 508 892 932
rect 120 480 892 508
rect 1132 932 1904 960
rect 1132 508 1820 932
rect 1884 508 1904 932
rect 1132 480 1904 508
rect 2144 932 2916 960
rect 2144 508 2832 932
rect 2896 508 2916 932
rect 2144 480 2916 508
rect -2916 212 -2144 240
rect -2916 -212 -2228 212
rect -2164 -212 -2144 212
rect -2916 -240 -2144 -212
rect -1904 212 -1132 240
rect -1904 -212 -1216 212
rect -1152 -212 -1132 212
rect -1904 -240 -1132 -212
rect -892 212 -120 240
rect -892 -212 -204 212
rect -140 -212 -120 212
rect -892 -240 -120 -212
rect 120 212 892 240
rect 120 -212 808 212
rect 872 -212 892 212
rect 120 -240 892 -212
rect 1132 212 1904 240
rect 1132 -212 1820 212
rect 1884 -212 1904 212
rect 1132 -240 1904 -212
rect 2144 212 2916 240
rect 2144 -212 2832 212
rect 2896 -212 2916 212
rect 2144 -240 2916 -212
rect -2916 -508 -2144 -480
rect -2916 -932 -2228 -508
rect -2164 -932 -2144 -508
rect -2916 -960 -2144 -932
rect -1904 -508 -1132 -480
rect -1904 -932 -1216 -508
rect -1152 -932 -1132 -508
rect -1904 -960 -1132 -932
rect -892 -508 -120 -480
rect -892 -932 -204 -508
rect -140 -932 -120 -508
rect -892 -960 -120 -932
rect 120 -508 892 -480
rect 120 -932 808 -508
rect 872 -932 892 -508
rect 120 -960 892 -932
rect 1132 -508 1904 -480
rect 1132 -932 1820 -508
rect 1884 -932 1904 -508
rect 1132 -960 1904 -932
rect 2144 -508 2916 -480
rect 2144 -932 2832 -508
rect 2896 -932 2916 -508
rect 2144 -960 2916 -932
rect -2916 -1228 -2144 -1200
rect -2916 -1652 -2228 -1228
rect -2164 -1652 -2144 -1228
rect -2916 -1680 -2144 -1652
rect -1904 -1228 -1132 -1200
rect -1904 -1652 -1216 -1228
rect -1152 -1652 -1132 -1228
rect -1904 -1680 -1132 -1652
rect -892 -1228 -120 -1200
rect -892 -1652 -204 -1228
rect -140 -1652 -120 -1228
rect -892 -1680 -120 -1652
rect 120 -1228 892 -1200
rect 120 -1652 808 -1228
rect 872 -1652 892 -1228
rect 120 -1680 892 -1652
rect 1132 -1228 1904 -1200
rect 1132 -1652 1820 -1228
rect 1884 -1652 1904 -1228
rect 1132 -1680 1904 -1652
rect 2144 -1228 2916 -1200
rect 2144 -1652 2832 -1228
rect 2896 -1652 2916 -1228
rect 2144 -1680 2916 -1652
rect -2916 -1948 -2144 -1920
rect -2916 -2372 -2228 -1948
rect -2164 -2372 -2144 -1948
rect -2916 -2400 -2144 -2372
rect -1904 -1948 -1132 -1920
rect -1904 -2372 -1216 -1948
rect -1152 -2372 -1132 -1948
rect -1904 -2400 -1132 -2372
rect -892 -1948 -120 -1920
rect -892 -2372 -204 -1948
rect -140 -2372 -120 -1948
rect -892 -2400 -120 -2372
rect 120 -1948 892 -1920
rect 120 -2372 808 -1948
rect 872 -2372 892 -1948
rect 120 -2400 892 -2372
rect 1132 -1948 1904 -1920
rect 1132 -2372 1820 -1948
rect 1884 -2372 1904 -1948
rect 1132 -2400 1904 -2372
rect 2144 -1948 2916 -1920
rect 2144 -2372 2832 -1948
rect 2896 -2372 2916 -1948
rect 2144 -2400 2916 -2372
<< via3 >>
rect -2228 1948 -2164 2372
rect -1216 1948 -1152 2372
rect -204 1948 -140 2372
rect 808 1948 872 2372
rect 1820 1948 1884 2372
rect 2832 1948 2896 2372
rect -2228 1228 -2164 1652
rect -1216 1228 -1152 1652
rect -204 1228 -140 1652
rect 808 1228 872 1652
rect 1820 1228 1884 1652
rect 2832 1228 2896 1652
rect -2228 508 -2164 932
rect -1216 508 -1152 932
rect -204 508 -140 932
rect 808 508 872 932
rect 1820 508 1884 932
rect 2832 508 2896 932
rect -2228 -212 -2164 212
rect -1216 -212 -1152 212
rect -204 -212 -140 212
rect 808 -212 872 212
rect 1820 -212 1884 212
rect 2832 -212 2896 212
rect -2228 -932 -2164 -508
rect -1216 -932 -1152 -508
rect -204 -932 -140 -508
rect 808 -932 872 -508
rect 1820 -932 1884 -508
rect 2832 -932 2896 -508
rect -2228 -1652 -2164 -1228
rect -1216 -1652 -1152 -1228
rect -204 -1652 -140 -1228
rect 808 -1652 872 -1228
rect 1820 -1652 1884 -1228
rect 2832 -1652 2896 -1228
rect -2228 -2372 -2164 -1948
rect -1216 -2372 -1152 -1948
rect -204 -2372 -140 -1948
rect 808 -2372 872 -1948
rect 1820 -2372 1884 -1948
rect 2832 -2372 2896 -1948
<< mimcap >>
rect -2876 2320 -2476 2360
rect -2876 2000 -2836 2320
rect -2516 2000 -2476 2320
rect -2876 1960 -2476 2000
rect -1864 2320 -1464 2360
rect -1864 2000 -1824 2320
rect -1504 2000 -1464 2320
rect -1864 1960 -1464 2000
rect -852 2320 -452 2360
rect -852 2000 -812 2320
rect -492 2000 -452 2320
rect -852 1960 -452 2000
rect 160 2320 560 2360
rect 160 2000 200 2320
rect 520 2000 560 2320
rect 160 1960 560 2000
rect 1172 2320 1572 2360
rect 1172 2000 1212 2320
rect 1532 2000 1572 2320
rect 1172 1960 1572 2000
rect 2184 2320 2584 2360
rect 2184 2000 2224 2320
rect 2544 2000 2584 2320
rect 2184 1960 2584 2000
rect -2876 1600 -2476 1640
rect -2876 1280 -2836 1600
rect -2516 1280 -2476 1600
rect -2876 1240 -2476 1280
rect -1864 1600 -1464 1640
rect -1864 1280 -1824 1600
rect -1504 1280 -1464 1600
rect -1864 1240 -1464 1280
rect -852 1600 -452 1640
rect -852 1280 -812 1600
rect -492 1280 -452 1600
rect -852 1240 -452 1280
rect 160 1600 560 1640
rect 160 1280 200 1600
rect 520 1280 560 1600
rect 160 1240 560 1280
rect 1172 1600 1572 1640
rect 1172 1280 1212 1600
rect 1532 1280 1572 1600
rect 1172 1240 1572 1280
rect 2184 1600 2584 1640
rect 2184 1280 2224 1600
rect 2544 1280 2584 1600
rect 2184 1240 2584 1280
rect -2876 880 -2476 920
rect -2876 560 -2836 880
rect -2516 560 -2476 880
rect -2876 520 -2476 560
rect -1864 880 -1464 920
rect -1864 560 -1824 880
rect -1504 560 -1464 880
rect -1864 520 -1464 560
rect -852 880 -452 920
rect -852 560 -812 880
rect -492 560 -452 880
rect -852 520 -452 560
rect 160 880 560 920
rect 160 560 200 880
rect 520 560 560 880
rect 160 520 560 560
rect 1172 880 1572 920
rect 1172 560 1212 880
rect 1532 560 1572 880
rect 1172 520 1572 560
rect 2184 880 2584 920
rect 2184 560 2224 880
rect 2544 560 2584 880
rect 2184 520 2584 560
rect -2876 160 -2476 200
rect -2876 -160 -2836 160
rect -2516 -160 -2476 160
rect -2876 -200 -2476 -160
rect -1864 160 -1464 200
rect -1864 -160 -1824 160
rect -1504 -160 -1464 160
rect -1864 -200 -1464 -160
rect -852 160 -452 200
rect -852 -160 -812 160
rect -492 -160 -452 160
rect -852 -200 -452 -160
rect 160 160 560 200
rect 160 -160 200 160
rect 520 -160 560 160
rect 160 -200 560 -160
rect 1172 160 1572 200
rect 1172 -160 1212 160
rect 1532 -160 1572 160
rect 1172 -200 1572 -160
rect 2184 160 2584 200
rect 2184 -160 2224 160
rect 2544 -160 2584 160
rect 2184 -200 2584 -160
rect -2876 -560 -2476 -520
rect -2876 -880 -2836 -560
rect -2516 -880 -2476 -560
rect -2876 -920 -2476 -880
rect -1864 -560 -1464 -520
rect -1864 -880 -1824 -560
rect -1504 -880 -1464 -560
rect -1864 -920 -1464 -880
rect -852 -560 -452 -520
rect -852 -880 -812 -560
rect -492 -880 -452 -560
rect -852 -920 -452 -880
rect 160 -560 560 -520
rect 160 -880 200 -560
rect 520 -880 560 -560
rect 160 -920 560 -880
rect 1172 -560 1572 -520
rect 1172 -880 1212 -560
rect 1532 -880 1572 -560
rect 1172 -920 1572 -880
rect 2184 -560 2584 -520
rect 2184 -880 2224 -560
rect 2544 -880 2584 -560
rect 2184 -920 2584 -880
rect -2876 -1280 -2476 -1240
rect -2876 -1600 -2836 -1280
rect -2516 -1600 -2476 -1280
rect -2876 -1640 -2476 -1600
rect -1864 -1280 -1464 -1240
rect -1864 -1600 -1824 -1280
rect -1504 -1600 -1464 -1280
rect -1864 -1640 -1464 -1600
rect -852 -1280 -452 -1240
rect -852 -1600 -812 -1280
rect -492 -1600 -452 -1280
rect -852 -1640 -452 -1600
rect 160 -1280 560 -1240
rect 160 -1600 200 -1280
rect 520 -1600 560 -1280
rect 160 -1640 560 -1600
rect 1172 -1280 1572 -1240
rect 1172 -1600 1212 -1280
rect 1532 -1600 1572 -1280
rect 1172 -1640 1572 -1600
rect 2184 -1280 2584 -1240
rect 2184 -1600 2224 -1280
rect 2544 -1600 2584 -1280
rect 2184 -1640 2584 -1600
rect -2876 -2000 -2476 -1960
rect -2876 -2320 -2836 -2000
rect -2516 -2320 -2476 -2000
rect -2876 -2360 -2476 -2320
rect -1864 -2000 -1464 -1960
rect -1864 -2320 -1824 -2000
rect -1504 -2320 -1464 -2000
rect -1864 -2360 -1464 -2320
rect -852 -2000 -452 -1960
rect -852 -2320 -812 -2000
rect -492 -2320 -452 -2000
rect -852 -2360 -452 -2320
rect 160 -2000 560 -1960
rect 160 -2320 200 -2000
rect 520 -2320 560 -2000
rect 160 -2360 560 -2320
rect 1172 -2000 1572 -1960
rect 1172 -2320 1212 -2000
rect 1532 -2320 1572 -2000
rect 1172 -2360 1572 -2320
rect 2184 -2000 2584 -1960
rect 2184 -2320 2224 -2000
rect 2544 -2320 2584 -2000
rect 2184 -2360 2584 -2320
<< mimcapcontact >>
rect -2836 2000 -2516 2320
rect -1824 2000 -1504 2320
rect -812 2000 -492 2320
rect 200 2000 520 2320
rect 1212 2000 1532 2320
rect 2224 2000 2544 2320
rect -2836 1280 -2516 1600
rect -1824 1280 -1504 1600
rect -812 1280 -492 1600
rect 200 1280 520 1600
rect 1212 1280 1532 1600
rect 2224 1280 2544 1600
rect -2836 560 -2516 880
rect -1824 560 -1504 880
rect -812 560 -492 880
rect 200 560 520 880
rect 1212 560 1532 880
rect 2224 560 2544 880
rect -2836 -160 -2516 160
rect -1824 -160 -1504 160
rect -812 -160 -492 160
rect 200 -160 520 160
rect 1212 -160 1532 160
rect 2224 -160 2544 160
rect -2836 -880 -2516 -560
rect -1824 -880 -1504 -560
rect -812 -880 -492 -560
rect 200 -880 520 -560
rect 1212 -880 1532 -560
rect 2224 -880 2544 -560
rect -2836 -1600 -2516 -1280
rect -1824 -1600 -1504 -1280
rect -812 -1600 -492 -1280
rect 200 -1600 520 -1280
rect 1212 -1600 1532 -1280
rect 2224 -1600 2544 -1280
rect -2836 -2320 -2516 -2000
rect -1824 -2320 -1504 -2000
rect -812 -2320 -492 -2000
rect 200 -2320 520 -2000
rect 1212 -2320 1532 -2000
rect 2224 -2320 2544 -2000
<< metal4 >>
rect -2244 2372 -2148 2388
rect -2837 2320 -2515 2321
rect -2837 2000 -2836 2320
rect -2516 2000 -2515 2320
rect -2837 1999 -2515 2000
rect -2244 1948 -2228 2372
rect -2164 1948 -2148 2372
rect -1232 2372 -1136 2388
rect -1825 2320 -1503 2321
rect -1825 2000 -1824 2320
rect -1504 2000 -1503 2320
rect -1825 1999 -1503 2000
rect -2244 1932 -2148 1948
rect -1232 1948 -1216 2372
rect -1152 1948 -1136 2372
rect -220 2372 -124 2388
rect -813 2320 -491 2321
rect -813 2000 -812 2320
rect -492 2000 -491 2320
rect -813 1999 -491 2000
rect -1232 1932 -1136 1948
rect -220 1948 -204 2372
rect -140 1948 -124 2372
rect 792 2372 888 2388
rect 199 2320 521 2321
rect 199 2000 200 2320
rect 520 2000 521 2320
rect 199 1999 521 2000
rect -220 1932 -124 1948
rect 792 1948 808 2372
rect 872 1948 888 2372
rect 1804 2372 1900 2388
rect 1211 2320 1533 2321
rect 1211 2000 1212 2320
rect 1532 2000 1533 2320
rect 1211 1999 1533 2000
rect 792 1932 888 1948
rect 1804 1948 1820 2372
rect 1884 1948 1900 2372
rect 2816 2372 2912 2388
rect 2223 2320 2545 2321
rect 2223 2000 2224 2320
rect 2544 2000 2545 2320
rect 2223 1999 2545 2000
rect 1804 1932 1900 1948
rect 2816 1948 2832 2372
rect 2896 1948 2912 2372
rect 2816 1932 2912 1948
rect -2244 1652 -2148 1668
rect -2837 1600 -2515 1601
rect -2837 1280 -2836 1600
rect -2516 1280 -2515 1600
rect -2837 1279 -2515 1280
rect -2244 1228 -2228 1652
rect -2164 1228 -2148 1652
rect -1232 1652 -1136 1668
rect -1825 1600 -1503 1601
rect -1825 1280 -1824 1600
rect -1504 1280 -1503 1600
rect -1825 1279 -1503 1280
rect -2244 1212 -2148 1228
rect -1232 1228 -1216 1652
rect -1152 1228 -1136 1652
rect -220 1652 -124 1668
rect -813 1600 -491 1601
rect -813 1280 -812 1600
rect -492 1280 -491 1600
rect -813 1279 -491 1280
rect -1232 1212 -1136 1228
rect -220 1228 -204 1652
rect -140 1228 -124 1652
rect 792 1652 888 1668
rect 199 1600 521 1601
rect 199 1280 200 1600
rect 520 1280 521 1600
rect 199 1279 521 1280
rect -220 1212 -124 1228
rect 792 1228 808 1652
rect 872 1228 888 1652
rect 1804 1652 1900 1668
rect 1211 1600 1533 1601
rect 1211 1280 1212 1600
rect 1532 1280 1533 1600
rect 1211 1279 1533 1280
rect 792 1212 888 1228
rect 1804 1228 1820 1652
rect 1884 1228 1900 1652
rect 2816 1652 2912 1668
rect 2223 1600 2545 1601
rect 2223 1280 2224 1600
rect 2544 1280 2545 1600
rect 2223 1279 2545 1280
rect 1804 1212 1900 1228
rect 2816 1228 2832 1652
rect 2896 1228 2912 1652
rect 2816 1212 2912 1228
rect -2244 932 -2148 948
rect -2837 880 -2515 881
rect -2837 560 -2836 880
rect -2516 560 -2515 880
rect -2837 559 -2515 560
rect -2244 508 -2228 932
rect -2164 508 -2148 932
rect -1232 932 -1136 948
rect -1825 880 -1503 881
rect -1825 560 -1824 880
rect -1504 560 -1503 880
rect -1825 559 -1503 560
rect -2244 492 -2148 508
rect -1232 508 -1216 932
rect -1152 508 -1136 932
rect -220 932 -124 948
rect -813 880 -491 881
rect -813 560 -812 880
rect -492 560 -491 880
rect -813 559 -491 560
rect -1232 492 -1136 508
rect -220 508 -204 932
rect -140 508 -124 932
rect 792 932 888 948
rect 199 880 521 881
rect 199 560 200 880
rect 520 560 521 880
rect 199 559 521 560
rect -220 492 -124 508
rect 792 508 808 932
rect 872 508 888 932
rect 1804 932 1900 948
rect 1211 880 1533 881
rect 1211 560 1212 880
rect 1532 560 1533 880
rect 1211 559 1533 560
rect 792 492 888 508
rect 1804 508 1820 932
rect 1884 508 1900 932
rect 2816 932 2912 948
rect 2223 880 2545 881
rect 2223 560 2224 880
rect 2544 560 2545 880
rect 2223 559 2545 560
rect 1804 492 1900 508
rect 2816 508 2832 932
rect 2896 508 2912 932
rect 2816 492 2912 508
rect -2244 212 -2148 228
rect -2837 160 -2515 161
rect -2837 -160 -2836 160
rect -2516 -160 -2515 160
rect -2837 -161 -2515 -160
rect -2244 -212 -2228 212
rect -2164 -212 -2148 212
rect -1232 212 -1136 228
rect -1825 160 -1503 161
rect -1825 -160 -1824 160
rect -1504 -160 -1503 160
rect -1825 -161 -1503 -160
rect -2244 -228 -2148 -212
rect -1232 -212 -1216 212
rect -1152 -212 -1136 212
rect -220 212 -124 228
rect -813 160 -491 161
rect -813 -160 -812 160
rect -492 -160 -491 160
rect -813 -161 -491 -160
rect -1232 -228 -1136 -212
rect -220 -212 -204 212
rect -140 -212 -124 212
rect 792 212 888 228
rect 199 160 521 161
rect 199 -160 200 160
rect 520 -160 521 160
rect 199 -161 521 -160
rect -220 -228 -124 -212
rect 792 -212 808 212
rect 872 -212 888 212
rect 1804 212 1900 228
rect 1211 160 1533 161
rect 1211 -160 1212 160
rect 1532 -160 1533 160
rect 1211 -161 1533 -160
rect 792 -228 888 -212
rect 1804 -212 1820 212
rect 1884 -212 1900 212
rect 2816 212 2912 228
rect 2223 160 2545 161
rect 2223 -160 2224 160
rect 2544 -160 2545 160
rect 2223 -161 2545 -160
rect 1804 -228 1900 -212
rect 2816 -212 2832 212
rect 2896 -212 2912 212
rect 2816 -228 2912 -212
rect -2244 -508 -2148 -492
rect -2837 -560 -2515 -559
rect -2837 -880 -2836 -560
rect -2516 -880 -2515 -560
rect -2837 -881 -2515 -880
rect -2244 -932 -2228 -508
rect -2164 -932 -2148 -508
rect -1232 -508 -1136 -492
rect -1825 -560 -1503 -559
rect -1825 -880 -1824 -560
rect -1504 -880 -1503 -560
rect -1825 -881 -1503 -880
rect -2244 -948 -2148 -932
rect -1232 -932 -1216 -508
rect -1152 -932 -1136 -508
rect -220 -508 -124 -492
rect -813 -560 -491 -559
rect -813 -880 -812 -560
rect -492 -880 -491 -560
rect -813 -881 -491 -880
rect -1232 -948 -1136 -932
rect -220 -932 -204 -508
rect -140 -932 -124 -508
rect 792 -508 888 -492
rect 199 -560 521 -559
rect 199 -880 200 -560
rect 520 -880 521 -560
rect 199 -881 521 -880
rect -220 -948 -124 -932
rect 792 -932 808 -508
rect 872 -932 888 -508
rect 1804 -508 1900 -492
rect 1211 -560 1533 -559
rect 1211 -880 1212 -560
rect 1532 -880 1533 -560
rect 1211 -881 1533 -880
rect 792 -948 888 -932
rect 1804 -932 1820 -508
rect 1884 -932 1900 -508
rect 2816 -508 2912 -492
rect 2223 -560 2545 -559
rect 2223 -880 2224 -560
rect 2544 -880 2545 -560
rect 2223 -881 2545 -880
rect 1804 -948 1900 -932
rect 2816 -932 2832 -508
rect 2896 -932 2912 -508
rect 2816 -948 2912 -932
rect -2244 -1228 -2148 -1212
rect -2837 -1280 -2515 -1279
rect -2837 -1600 -2836 -1280
rect -2516 -1600 -2515 -1280
rect -2837 -1601 -2515 -1600
rect -2244 -1652 -2228 -1228
rect -2164 -1652 -2148 -1228
rect -1232 -1228 -1136 -1212
rect -1825 -1280 -1503 -1279
rect -1825 -1600 -1824 -1280
rect -1504 -1600 -1503 -1280
rect -1825 -1601 -1503 -1600
rect -2244 -1668 -2148 -1652
rect -1232 -1652 -1216 -1228
rect -1152 -1652 -1136 -1228
rect -220 -1228 -124 -1212
rect -813 -1280 -491 -1279
rect -813 -1600 -812 -1280
rect -492 -1600 -491 -1280
rect -813 -1601 -491 -1600
rect -1232 -1668 -1136 -1652
rect -220 -1652 -204 -1228
rect -140 -1652 -124 -1228
rect 792 -1228 888 -1212
rect 199 -1280 521 -1279
rect 199 -1600 200 -1280
rect 520 -1600 521 -1280
rect 199 -1601 521 -1600
rect -220 -1668 -124 -1652
rect 792 -1652 808 -1228
rect 872 -1652 888 -1228
rect 1804 -1228 1900 -1212
rect 1211 -1280 1533 -1279
rect 1211 -1600 1212 -1280
rect 1532 -1600 1533 -1280
rect 1211 -1601 1533 -1600
rect 792 -1668 888 -1652
rect 1804 -1652 1820 -1228
rect 1884 -1652 1900 -1228
rect 2816 -1228 2912 -1212
rect 2223 -1280 2545 -1279
rect 2223 -1600 2224 -1280
rect 2544 -1600 2545 -1280
rect 2223 -1601 2545 -1600
rect 1804 -1668 1900 -1652
rect 2816 -1652 2832 -1228
rect 2896 -1652 2912 -1228
rect 2816 -1668 2912 -1652
rect -2244 -1948 -2148 -1932
rect -2837 -2000 -2515 -1999
rect -2837 -2320 -2836 -2000
rect -2516 -2320 -2515 -2000
rect -2837 -2321 -2515 -2320
rect -2244 -2372 -2228 -1948
rect -2164 -2372 -2148 -1948
rect -1232 -1948 -1136 -1932
rect -1825 -2000 -1503 -1999
rect -1825 -2320 -1824 -2000
rect -1504 -2320 -1503 -2000
rect -1825 -2321 -1503 -2320
rect -2244 -2388 -2148 -2372
rect -1232 -2372 -1216 -1948
rect -1152 -2372 -1136 -1948
rect -220 -1948 -124 -1932
rect -813 -2000 -491 -1999
rect -813 -2320 -812 -2000
rect -492 -2320 -491 -2000
rect -813 -2321 -491 -2320
rect -1232 -2388 -1136 -2372
rect -220 -2372 -204 -1948
rect -140 -2372 -124 -1948
rect 792 -1948 888 -1932
rect 199 -2000 521 -1999
rect 199 -2320 200 -2000
rect 520 -2320 521 -2000
rect 199 -2321 521 -2320
rect -220 -2388 -124 -2372
rect 792 -2372 808 -1948
rect 872 -2372 888 -1948
rect 1804 -1948 1900 -1932
rect 1211 -2000 1533 -1999
rect 1211 -2320 1212 -2000
rect 1532 -2320 1533 -2000
rect 1211 -2321 1533 -2320
rect 792 -2388 888 -2372
rect 1804 -2372 1820 -1948
rect 1884 -2372 1900 -1948
rect 2816 -1948 2912 -1932
rect 2223 -2000 2545 -1999
rect 2223 -2320 2224 -2000
rect 2544 -2320 2545 -2000
rect 2223 -2321 2545 -2320
rect 1804 -2388 1900 -2372
rect 2816 -2372 2832 -1948
rect 2896 -2372 2912 -1948
rect 2816 -2388 2912 -2372
<< properties >>
string FIXED_BBOX 2144 1920 2624 2400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 6 ny 7 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
