magic
tech sky130A
magscale 1 2
timestamp 1749624948
<< error_p >>
rect -531 198 531 202
rect -531 -130 -501 198
rect -465 132 465 136
rect -465 -64 -435 132
rect 435 -64 465 132
rect 501 -130 531 198
<< nwell >>
rect -501 -164 501 198
<< mvpmos >>
rect -407 -64 -247 136
rect -189 -64 -29 136
rect 29 -64 189 136
rect 247 -64 407 136
<< mvpdiff >>
rect -465 124 -407 136
rect -465 -52 -453 124
rect -419 -52 -407 124
rect -465 -64 -407 -52
rect -247 124 -189 136
rect -247 -52 -235 124
rect -201 -52 -189 124
rect -247 -64 -189 -52
rect -29 124 29 136
rect -29 -52 -17 124
rect 17 -52 29 124
rect -29 -64 29 -52
rect 189 124 247 136
rect 189 -52 201 124
rect 235 -52 247 124
rect 189 -64 247 -52
rect 407 124 465 136
rect 407 -52 419 124
rect 453 -52 465 124
rect 407 -64 465 -52
<< mvpdiffc >>
rect -453 -52 -419 124
rect -235 -52 -201 124
rect -17 -52 17 124
rect 201 -52 235 124
rect 419 -52 453 124
<< poly >>
rect -407 136 -247 162
rect -189 136 -29 162
rect 29 136 189 162
rect 247 136 407 162
rect -407 -111 -247 -64
rect -407 -145 -391 -111
rect -263 -145 -247 -111
rect -407 -161 -247 -145
rect -189 -111 -29 -64
rect -189 -145 -173 -111
rect -45 -145 -29 -111
rect -189 -161 -29 -145
rect 29 -111 189 -64
rect 29 -145 45 -111
rect 173 -145 189 -111
rect 29 -161 189 -145
rect 247 -111 407 -64
rect 247 -145 263 -111
rect 391 -145 407 -111
rect 247 -161 407 -145
<< polycont >>
rect -391 -145 -263 -111
rect -173 -145 -45 -111
rect 45 -145 173 -111
rect 263 -145 391 -111
<< locali >>
rect -453 124 -419 140
rect -453 -68 -419 -52
rect -235 124 -201 140
rect -235 -68 -201 -52
rect -17 124 17 140
rect -17 -68 17 -52
rect 201 124 235 140
rect 201 -68 235 -52
rect 419 124 453 140
rect 419 -68 453 -52
rect -407 -145 -391 -111
rect -263 -145 -247 -111
rect -189 -145 -173 -111
rect -45 -145 -29 -111
rect 29 -145 45 -111
rect 173 -145 189 -111
rect 247 -145 263 -111
rect 391 -145 407 -111
<< viali >>
rect -453 -52 -419 124
rect -235 -52 -201 124
rect -17 -52 17 124
rect 201 -52 235 124
rect 419 -52 453 124
rect -391 -145 -263 -111
rect -173 -145 -45 -111
rect 45 -145 173 -111
rect 263 -145 391 -111
<< metal1 >>
rect -459 124 -413 136
rect -459 -52 -453 124
rect -419 -52 -413 124
rect -459 -64 -413 -52
rect -241 124 -195 136
rect -241 -52 -235 124
rect -201 -52 -195 124
rect -241 -64 -195 -52
rect -23 124 23 136
rect -23 -52 -17 124
rect 17 -52 23 124
rect -23 -64 23 -52
rect 195 124 241 136
rect 195 -52 201 124
rect 235 -52 241 124
rect 195 -64 241 -52
rect 413 124 459 136
rect 413 -52 419 124
rect 453 -52 459 124
rect 413 -64 459 -52
rect -403 -111 -251 -105
rect -403 -145 -391 -111
rect -263 -145 -251 -111
rect -403 -151 -251 -145
rect -185 -111 -33 -105
rect -185 -145 -173 -111
rect -45 -145 -33 -111
rect -185 -151 -33 -145
rect 33 -111 185 -105
rect 33 -145 45 -111
rect 173 -145 185 -111
rect 33 -151 185 -145
rect 251 -111 403 -105
rect 251 -145 263 -111
rect 391 -145 403 -111
rect 251 -151 403 -145
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 0.8 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
