magic
tech sky130A
magscale 1 2
timestamp 1748204885
<< checkpaint >>
rect -615 -23377 2375 -23351
rect -1313 -23440 2375 -23377
rect -1313 -23517 2792 -23440
rect -1313 -23596 3209 -23517
rect -1313 -23669 3626 -23596
rect -1313 -23738 4043 -23669
rect -1313 -23805 4460 -23738
rect -1313 -23874 4877 -23805
rect -1313 -23916 5294 -23874
rect -1313 -23989 7106 -23916
rect -1313 -24052 7667 -23989
rect -1313 -24125 8228 -24052
rect -1313 -24178 8789 -24125
rect -1313 -24253 9350 -24178
rect -1313 -24306 9911 -24253
rect -1313 -24379 10472 -24306
rect -1313 -24432 11033 -24379
rect -1313 -24495 11594 -24432
rect -1313 -24548 12155 -24495
rect -1313 -24623 12716 -24548
rect -1313 -24676 13277 -24623
rect -1313 -24739 13838 -24676
rect -1313 -24792 14399 -24739
rect -1313 -24855 14960 -24792
rect -1313 -24908 15521 -24855
rect -1313 -24971 16082 -24908
rect -1313 -25024 16643 -24971
rect -1313 -25087 17204 -25024
rect -1313 -25140 17765 -25087
rect -1313 -25193 18326 -25140
rect -1313 -25256 18887 -25193
rect -1313 -25319 19448 -25256
rect -1313 -25362 20009 -25319
rect -1313 -25425 20570 -25362
rect -1313 -25459 21131 -25425
rect -1313 -25565 23663 -25459
rect -1313 -25618 25073 -25565
rect -1313 -25671 25922 -25618
rect -1313 -25744 26771 -25671
rect -1313 -25777 27620 -25744
rect -1313 -25850 28469 -25777
rect -1313 -25923 29318 -25850
rect -1313 -25956 30167 -25923
rect -1313 -26029 31016 -25956
rect -1313 -26082 31865 -26029
rect -1313 -26135 32714 -26082
rect -1313 -26188 33563 -26135
rect -1313 -26241 34412 -26188
rect -1313 -26316 35261 -26241
rect -1313 -26369 36110 -26316
rect -1313 -26422 36959 -26369
rect -1313 -26475 37808 -26422
rect -1313 -26528 38657 -26475
rect -1313 -26581 39506 -26528
rect -1313 -26654 40355 -26581
rect -1313 -27313 41204 -26654
rect -964 -27366 41204 -27313
rect -615 -27419 41204 -27366
rect -198 -27472 41204 -27419
rect 219 -27525 41204 -27472
rect 636 -27578 41204 -27525
rect 1053 -27631 41204 -27578
rect 1470 -27684 41204 -27631
rect 1887 -27737 41204 -27684
rect 2304 -27790 41204 -27737
rect 2721 -27843 41204 -27790
rect 3138 -27896 41204 -27843
rect 3555 -27949 41204 -27896
rect 3972 -28002 41204 -27949
rect 4533 -28055 41204 -28002
rect 5094 -28108 41204 -28055
rect 5655 -28161 41204 -28108
rect 6216 -28214 41204 -28161
rect 6777 -28267 41204 -28214
rect 7338 -28320 41204 -28267
rect 7899 -28373 41204 -28320
rect 8460 -28426 41204 -28373
rect 9021 -28479 41204 -28426
rect 9582 -28532 41204 -28479
rect 10143 -28585 41204 -28532
rect 10704 -28638 41204 -28585
rect 11265 -28691 41204 -28638
rect 11826 -28744 41204 -28691
rect 12387 -28797 41204 -28744
rect 12948 -28850 41204 -28797
rect 13509 -28903 41204 -28850
rect 14070 -28956 41204 -28903
rect 14631 -29009 41204 -28956
rect 15192 -29062 41204 -29009
rect 15753 -29115 41204 -29062
rect 16314 -29168 41204 -29115
rect 16875 -29221 41204 -29168
rect 17436 -29274 41204 -29221
rect 17997 -29327 41204 -29274
rect 18558 -29380 41204 -29327
rect 19119 -29433 41204 -29380
rect 19680 -29486 41204 -29433
rect 20241 -29539 41204 -29486
rect 21090 -29592 41204 -29539
rect 21651 -29645 41204 -29592
rect 22500 -29698 41204 -29645
rect 23349 -29751 41204 -29698
rect 24198 -29804 41204 -29751
rect 25047 -29857 41204 -29804
rect 25896 -29910 41204 -29857
rect 26745 -29963 41204 -29910
rect 27594 -30016 41204 -29963
rect 28443 -30069 41204 -30016
rect 29292 -30122 41204 -30069
rect 30141 -30175 41204 -30122
rect 30990 -30228 41204 -30175
rect 31839 -30281 41204 -30228
rect 32688 -30334 41204 -30281
rect 33537 -30387 41204 -30334
rect 34386 -30440 41204 -30387
rect 35235 -30493 41204 -30440
rect 36084 -30546 41204 -30493
rect 36933 -30599 41204 -30546
rect 37782 -30652 41204 -30599
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
rect 0 -8400 200 -8200
rect 0 -8800 200 -8600
rect 0 -9200 200 -9000
rect 0 -9600 200 -9400
rect 0 -10000 200 -9800
rect 0 -10400 200 -10200
rect 0 -10800 200 -10600
rect 0 -11200 200 -11000
rect 0 -11600 200 -11400
rect 0 -12000 200 -11800
rect 0 -12400 200 -12200
rect 0 -12800 200 -12600
rect 0 -13200 200 -13000
rect 0 -13600 200 -13400
rect 0 -14000 200 -13800
rect 0 -14400 200 -14200
rect 0 -14800 200 -14600
rect 0 -15200 200 -15000
rect 0 -15600 200 -15400
rect 0 -16000 200 -15800
rect 0 -16400 200 -16200
rect 0 -16800 200 -16600
rect 0 -17200 200 -17000
rect 0 -17600 200 -17400
rect 0 -18000 200 -17800
rect 0 -18400 200 -18200
rect 0 -18800 200 -18600
rect 0 -19200 200 -19000
rect 0 -19600 200 -19400
rect 0 -20000 200 -19800
rect 0 -20400 200 -20200
rect 0 -20800 200 -20600
rect 0 -21200 200 -21000
rect 0 -21600 200 -21400
rect 0 -22000 200 -21800
rect 0 -22400 200 -22200
rect 0 -22800 200 -22600
rect 0 -23200 200 -23000
rect 0 -23600 200 -23400
rect 0 -24000 200 -23800
rect 0 -24400 200 -24200
rect 0 -24800 200 -24600
rect 0 -25200 200 -25000
rect 0 -25600 200 -25400
rect 0 -26000 200 -25800
use sky130_fd_pr__res_xhigh_po_0p35_RL62MD  XR1
timestamp 0
transform 1 0 148 0 1 -25345
box -201 -708 201 708
use sky130_fd_pr__res_xhigh_po_0p35_WTBJYY  XR2
timestamp 0
transform 1 0 497 0 1 -25414
box -201 -692 201 692
use sky130_fd_pr__res_xhigh_po_0p69_5QPZKM  XR3
timestamp 0
transform 1 0 880 0 1 -25385
box -235 -774 235 774
use sky130_fd_pr__res_xhigh_po_0p69_MKRCVN  XR4
timestamp 0
transform 1 0 1297 0 1 -25456
box -235 -756 235 756
use sky130_fd_pr__res_xhigh_po_0p69_BWLLCM  XR5
timestamp 0
transform 1 0 1714 0 1 -25521
box -235 -744 235 744
use sky130_fd_pr__res_xhigh_po_0p69_RP95CT  XR6
timestamp 0
transform 1 0 2131 0 1 -25587
box -235 -731 235 731
use sky130_fd_pr__res_xhigh_po_0p69_B9L8UC  XR7
timestamp 0
transform 1 0 2548 0 1 -25650
box -235 -721 235 721
use sky130_fd_pr__res_xhigh_po_0p69_3HJCGF  XR8
timestamp 0
transform 1 0 2965 0 1 -25711
box -235 -713 235 713
use sky130_fd_pr__res_xhigh_po_0p69_4KUEG2  XR9
timestamp 0
transform 1 0 3382 0 1 -25771
box -235 -706 235 706
use sky130_fd_pr__res_xhigh_po_0p69_THP23T  XR10
timestamp 0
transform 1 0 3799 0 1 -25832
box -235 -698 235 698
use sky130_fd_pr__res_xhigh_po_0p69_UCJEAS  XR11
timestamp 0
transform 1 0 4216 0 1 -25890
box -235 -693 235 693
use sky130_fd_pr__res_xhigh_po_0p69_PH3F3P  XR12
timestamp 0
transform 1 0 4633 0 1 -25948
box -235 -688 235 688
use sky130_fd_pr__res_xhigh_po_0p69_73P63X  XR13
timestamp 0
transform 1 0 5050 0 1 -26006
box -235 -683 235 683
use sky130_fd_pr__res_xhigh_po_1p41_J3VGEN  XR14
timestamp 0
transform 1 0 5539 0 1 -25959
box -307 -783 307 783
use sky130_fd_pr__res_xhigh_po_1p41_FMVSM8  XR15
timestamp 0
transform 1 0 6100 0 1 -26022
box -307 -773 307 773
use sky130_fd_pr__res_xhigh_po_1p41_TSKUDA  XR16
timestamp 0
transform 1 0 6661 0 1 -26080
box -307 -768 307 768
use sky130_fd_pr__res_xhigh_po_1p41_S5LQAA  XR17
timestamp 0
transform 1 0 7222 0 1 -26143
box -307 -758 307 758
use sky130_fd_pr__res_xhigh_po_1p41_S5LQAA  XR18
timestamp 0
transform 1 0 7783 0 1 -26196
box -307 -758 307 758
use sky130_fd_pr__res_xhigh_po_1p41_HUF2GN  XR19
timestamp 0
transform 1 0 8344 0 1 -26260
box -307 -747 307 747
use sky130_fd_pr__res_xhigh_po_1p41_HUF2GN  XR20
timestamp 0
transform 1 0 8905 0 1 -26313
box -307 -747 307 747
use sky130_fd_pr__res_xhigh_po_1p41_9HH8QQ  XR21
timestamp 0
transform 1 0 9466 0 1 -26376
box -307 -737 307 737
use sky130_fd_pr__res_xhigh_po_1p41_9HH8QQ  XR22
timestamp 0
transform 1 0 10027 0 1 -26429
box -307 -737 307 737
use sky130_fd_pr__res_xhigh_po_1p41_X2L423  XR23
timestamp 0
transform 1 0 10588 0 1 -26487
box -307 -732 307 732
use sky130_fd_pr__res_xhigh_po_1p41_X2L423  XR24
timestamp 0
transform 1 0 11149 0 1 -26540
box -307 -732 307 732
use sky130_fd_pr__res_xhigh_po_1p41_QEVKRF  XR25
timestamp 0
transform 1 0 11710 0 1 -26604
box -307 -721 307 721
use sky130_fd_pr__res_xhigh_po_1p41_QEVKRF  XR26
timestamp 0
transform 1 0 12271 0 1 -26657
box -307 -721 307 721
use sky130_fd_pr__res_xhigh_po_1p41_7FPTVH  XR27
timestamp 0
transform 1 0 12832 0 1 -26715
box -307 -716 307 716
use sky130_fd_pr__res_xhigh_po_1p41_7FPTVH  XR28
timestamp 0
transform 1 0 13393 0 1 -26768
box -307 -716 307 716
use sky130_fd_pr__res_xhigh_po_1p41_4MEUZY  XR29
timestamp 0
transform 1 0 13954 0 1 -26826
box -307 -711 307 711
use sky130_fd_pr__res_xhigh_po_1p41_4MEUZY  XR30
timestamp 0
transform 1 0 14515 0 1 -26879
box -307 -711 307 711
use sky130_fd_pr__res_xhigh_po_1p41_YPFF3H  XR31
timestamp 0
transform 1 0 15076 0 1 -26937
box -307 -706 307 706
use sky130_fd_pr__res_xhigh_po_1p41_YPFF3H  XR32
timestamp 0
transform 1 0 15637 0 1 -26990
box -307 -706 307 706
use sky130_fd_pr__res_xhigh_po_1p41_MWY8WZ  XR33
timestamp 0
transform 1 0 16198 0 1 -27048
box -307 -701 307 701
use sky130_fd_pr__res_xhigh_po_1p41_MWY8WZ  XR34
timestamp 0
transform 1 0 16759 0 1 -27101
box -307 -701 307 701
use sky130_fd_pr__res_xhigh_po_1p41_MWY8WZ  XR35
timestamp 0
transform 1 0 17320 0 1 -27154
box -307 -701 307 701
use sky130_fd_pr__res_xhigh_po_1p41_LSX63M  XR36
timestamp 0
transform 1 0 17881 0 1 -27212
box -307 -696 307 696
use sky130_fd_pr__res_xhigh_po_1p41_27TN7E  XR37
timestamp 0
transform 1 0 18442 0 1 -27270
box -307 -691 307 691
use sky130_fd_pr__res_xhigh_po_1p41_LSX63M  XR38
timestamp 0
transform 1 0 19003 0 1 -27318
box -307 -696 307 696
use sky130_fd_pr__res_xhigh_po_1p41_27TN7E  XR39
timestamp 0
transform 1 0 19564 0 1 -27376
box -307 -691 307 691
use sky130_fd_pr__res_xhigh_po_1p41_N3JE47  XR40
timestamp 0
transform 1 0 20125 0 1 -27435
box -307 -685 307 685
use sky130_fd_pr__res_xhigh_po_1p41_27TN7E  XR41
timestamp 0
transform 1 0 20686 0 1 -27482
box -307 -691 307 691
use sky130_fd_pr__res_xhigh_po_1p41_N3JE47  XR42
timestamp 0
transform 1 0 21247 0 1 -27541
box -307 -685 307 685
use sky130_fd_pr__res_xhigh_po_2p85_3C9AJP  XR43
timestamp 0
transform 1 0 21952 0 1 -27499
box -451 -780 451 780
use sky130_fd_pr__res_xhigh_po_1p41_N3JE47  XR44
timestamp 0
transform 1 0 22657 0 1 -27647
box -307 -685 307 685
use sky130_fd_pr__res_xhigh_po_2p85_3C9AJP  XR45
timestamp 0
transform 1 0 23362 0 1 -27605
box -451 -780 451 780
use sky130_fd_pr__res_xhigh_po_2p85_3C9AJP  XR46
timestamp 0
transform 1 0 24211 0 1 -27658
box -451 -780 451 780
use sky130_fd_pr__res_xhigh_po_2p85_3C9AJP  XR47
timestamp 0
transform 1 0 25060 0 1 -27711
box -451 -780 451 780
use sky130_fd_pr__res_xhigh_po_2p85_R7UNSU  XR48
timestamp 0
transform 1 0 25909 0 1 -27774
box -451 -770 451 770
use sky130_fd_pr__res_xhigh_po_2p85_3C9AJP  XR49
timestamp 0
transform 1 0 26758 0 1 -27817
box -451 -780 451 780
use sky130_fd_pr__res_xhigh_po_2p85_R7UNSU  XR50
timestamp 0
transform 1 0 27607 0 1 -27880
box -451 -770 451 770
use sky130_fd_pr__res_xhigh_po_2p85_YV8936  XR51
timestamp 0
transform 1 0 28456 0 1 -27943
box -451 -760 451 760
use sky130_fd_pr__res_xhigh_po_2p85_R7UNSU  XR52
timestamp 0
transform 1 0 29305 0 1 -27986
box -451 -770 451 770
use sky130_fd_pr__res_xhigh_po_2p85_YV8936  XR53
timestamp 0
transform 1 0 30154 0 1 -28049
box -451 -760 451 760
use sky130_fd_pr__res_xhigh_po_2p85_YV8936  XR54
timestamp 0
transform 1 0 31003 0 1 -28102
box -451 -760 451 760
use sky130_fd_pr__res_xhigh_po_2p85_YV8936  XR55
timestamp 0
transform 1 0 31852 0 1 -28155
box -451 -760 451 760
use sky130_fd_pr__res_xhigh_po_2p85_YV8936  XR56
timestamp 0
transform 1 0 32701 0 1 -28208
box -451 -760 451 760
use sky130_fd_pr__res_xhigh_po_2p85_YV8936  XR57
timestamp 0
transform 1 0 33550 0 1 -28261
box -451 -760 451 760
use sky130_fd_pr__res_xhigh_po_2p85_ZW9B2M  XR58
timestamp 0
transform 1 0 34399 0 1 -28325
box -451 -749 451 749
use sky130_fd_pr__res_xhigh_po_2p85_ZW9B2M  XR59
timestamp 0
transform 1 0 35248 0 1 -28378
box -451 -749 451 749
use sky130_fd_pr__res_xhigh_po_2p85_ZW9B2M  XR60
timestamp 0
transform 1 0 36097 0 1 -28431
box -451 -749 451 749
use sky130_fd_pr__res_xhigh_po_2p85_ZW9B2M  XR61
timestamp 0
transform 1 0 36946 0 1 -28484
box -451 -749 451 749
use sky130_fd_pr__res_xhigh_po_2p85_ZW9B2M  XR62
timestamp 0
transform 1 0 37795 0 1 -28537
box -451 -749 451 749
use sky130_fd_pr__res_xhigh_po_2p85_ZW9B2M  XR63
timestamp 0
transform 1 0 38644 0 1 -28590
box -451 -749 451 749
use sky130_fd_pr__res_xhigh_po_2p85_UG8474  XR64
timestamp 0
transform 1 0 39493 0 1 -28653
box -451 -739 451 739
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 v0
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 v1
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 v2
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 v3
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 v4
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 v5
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 v6
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 v7
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 v8
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 v9
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 v10
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 v11
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 v12
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 v13
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 v14
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 v15
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 v16
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 v17
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 v18
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 v19
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 v20
port 20 nsew
flabel metal1 0 -8400 200 -8200 0 FreeSans 256 0 0 0 v21
port 21 nsew
flabel metal1 0 -8800 200 -8600 0 FreeSans 256 0 0 0 v22
port 22 nsew
flabel metal1 0 -9200 200 -9000 0 FreeSans 256 0 0 0 v23
port 23 nsew
flabel metal1 0 -9600 200 -9400 0 FreeSans 256 0 0 0 v24
port 24 nsew
flabel metal1 0 -10000 200 -9800 0 FreeSans 256 0 0 0 v25
port 25 nsew
flabel metal1 0 -10400 200 -10200 0 FreeSans 256 0 0 0 v26
port 26 nsew
flabel metal1 0 -10800 200 -10600 0 FreeSans 256 0 0 0 v27
port 27 nsew
flabel metal1 0 -11200 200 -11000 0 FreeSans 256 0 0 0 v28
port 28 nsew
flabel metal1 0 -11600 200 -11400 0 FreeSans 256 0 0 0 v29
port 29 nsew
flabel metal1 0 -12000 200 -11800 0 FreeSans 256 0 0 0 v30
port 30 nsew
flabel metal1 0 -12400 200 -12200 0 FreeSans 256 0 0 0 v31
port 31 nsew
flabel metal1 0 -12800 200 -12600 0 FreeSans 256 0 0 0 v32
port 32 nsew
flabel metal1 0 -13200 200 -13000 0 FreeSans 256 0 0 0 v33
port 33 nsew
flabel metal1 0 -13600 200 -13400 0 FreeSans 256 0 0 0 v34
port 34 nsew
flabel metal1 0 -14000 200 -13800 0 FreeSans 256 0 0 0 v35
port 35 nsew
flabel metal1 0 -14400 200 -14200 0 FreeSans 256 0 0 0 v36
port 36 nsew
flabel metal1 0 -14800 200 -14600 0 FreeSans 256 0 0 0 v37
port 37 nsew
flabel metal1 0 -15200 200 -15000 0 FreeSans 256 0 0 0 v38
port 38 nsew
flabel metal1 0 -15600 200 -15400 0 FreeSans 256 0 0 0 v39
port 39 nsew
flabel metal1 0 -16000 200 -15800 0 FreeSans 256 0 0 0 v40
port 40 nsew
flabel metal1 0 -16400 200 -16200 0 FreeSans 256 0 0 0 v41
port 41 nsew
flabel metal1 0 -16800 200 -16600 0 FreeSans 256 0 0 0 v42
port 42 nsew
flabel metal1 0 -17200 200 -17000 0 FreeSans 256 0 0 0 v43
port 43 nsew
flabel metal1 0 -17600 200 -17400 0 FreeSans 256 0 0 0 v44
port 44 nsew
flabel metal1 0 -18000 200 -17800 0 FreeSans 256 0 0 0 v45
port 45 nsew
flabel metal1 0 -18400 200 -18200 0 FreeSans 256 0 0 0 v46
port 46 nsew
flabel metal1 0 -18800 200 -18600 0 FreeSans 256 0 0 0 v47
port 47 nsew
flabel metal1 0 -19200 200 -19000 0 FreeSans 256 0 0 0 v48
port 48 nsew
flabel metal1 0 -19600 200 -19400 0 FreeSans 256 0 0 0 v49
port 49 nsew
flabel metal1 0 -20000 200 -19800 0 FreeSans 256 0 0 0 v50
port 50 nsew
flabel metal1 0 -20400 200 -20200 0 FreeSans 256 0 0 0 v51
port 51 nsew
flabel metal1 0 -20800 200 -20600 0 FreeSans 256 0 0 0 v52
port 52 nsew
flabel metal1 0 -21200 200 -21000 0 FreeSans 256 0 0 0 v53
port 53 nsew
flabel metal1 0 -21600 200 -21400 0 FreeSans 256 0 0 0 v54
port 54 nsew
flabel metal1 0 -22000 200 -21800 0 FreeSans 256 0 0 0 v55
port 55 nsew
flabel metal1 0 -22400 200 -22200 0 FreeSans 256 0 0 0 v56
port 56 nsew
flabel metal1 0 -22800 200 -22600 0 FreeSans 256 0 0 0 v57
port 57 nsew
flabel metal1 0 -23200 200 -23000 0 FreeSans 256 0 0 0 v58
port 58 nsew
flabel metal1 0 -23600 200 -23400 0 FreeSans 256 0 0 0 v59
port 59 nsew
flabel metal1 0 -24000 200 -23800 0 FreeSans 256 0 0 0 v60
port 60 nsew
flabel metal1 0 -24400 200 -24200 0 FreeSans 256 0 0 0 v61
port 61 nsew
flabel metal1 0 -24800 200 -24600 0 FreeSans 256 0 0 0 v62
port 62 nsew
flabel metal1 0 -25200 200 -25000 0 FreeSans 256 0 0 0 v63
port 63 nsew
flabel metal1 0 -25600 200 -25400 0 FreeSans 256 0 0 0 v64
port 64 nsew
flabel metal1 0 -26000 200 -25800 0 FreeSans 256 0 0 0 gnd
port 65 nsew
<< end >>
