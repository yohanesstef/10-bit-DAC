magic
tech sky130A
magscale 1 2
timestamp 1749376058
<< metal1 >>
rect 1487 3483 1547 3489
rect 1399 3307 1459 3313
rect 1311 3131 1371 3137
rect 1311 2955 1371 3071
rect 1399 2955 1459 3247
rect 1487 2955 1547 3423
<< via1 >>
rect 1487 3423 1547 3483
rect 1399 3247 1459 3307
rect 1311 3071 1371 3131
<< metal2 >>
rect 1057 3423 1487 3483
rect 1547 3423 1553 3483
rect 1057 3247 1399 3307
rect 1459 3247 1465 3307
rect 1057 3071 1311 3131
rect 1371 3071 1377 3131
<< end >>
