magic
tech sky130A
magscale 1 2
timestamp 1750825354
<< viali >>
rect 184 3714 218 3748
rect 364 3713 398 3747
rect 525 3711 559 3745
rect 700 3714 734 3748
rect 866 3712 900 3746
rect 1045 3711 1079 3745
rect 1214 3712 1248 3746
rect 1387 3713 1421 3747
<< metal1 >>
rect 44 3954 1468 4102
rect 262 3760 322 3766
rect 170 3748 262 3760
rect 170 3714 184 3748
rect 218 3714 262 3748
rect 170 3700 262 3714
rect 262 3694 322 3700
rect 350 3760 410 3766
rect 604 3760 664 3766
rect 513 3745 604 3760
rect 513 3711 525 3745
rect 559 3711 604 3745
rect 513 3700 604 3711
rect 350 3694 410 3700
rect 604 3694 664 3700
rect 692 3760 752 3766
rect 946 3760 1006 3766
rect 853 3746 946 3760
rect 853 3712 866 3746
rect 900 3712 946 3746
rect 853 3700 946 3712
rect 692 3694 752 3700
rect 946 3694 1006 3700
rect 1034 3760 1094 3766
rect 1288 3760 1348 3766
rect 1203 3746 1288 3760
rect 1203 3712 1214 3746
rect 1248 3712 1288 3746
rect 1203 3700 1288 3712
rect 1034 3694 1094 3700
rect 1288 3694 1348 3700
rect 1376 3760 1436 3766
rect 1376 3694 1436 3700
rect 44 3230 1468 3390
<< via1 >>
rect 262 3700 322 3760
rect 350 3747 410 3760
rect 350 3713 364 3747
rect 364 3713 398 3747
rect 398 3713 410 3747
rect 350 3700 410 3713
rect 604 3700 664 3760
rect 692 3748 752 3760
rect 692 3714 700 3748
rect 700 3714 734 3748
rect 734 3714 752 3748
rect 692 3700 752 3714
rect 946 3700 1006 3760
rect 1034 3745 1094 3760
rect 1034 3711 1045 3745
rect 1045 3711 1079 3745
rect 1079 3711 1094 3745
rect 1034 3700 1094 3711
rect 1288 3700 1348 3760
rect 1376 3747 1436 3760
rect 1376 3713 1387 3747
rect 1387 3713 1421 3747
rect 1421 3713 1436 3747
rect 1376 3700 1436 3713
<< metal2 >>
rect 262 3760 322 4102
rect 262 3694 322 3700
rect 350 3760 410 4102
rect 350 3260 410 3700
rect 604 3760 664 4102
rect 604 3694 664 3700
rect 692 3760 752 4102
rect 692 3260 752 3700
rect 946 3760 1006 4102
rect 946 3694 1006 3700
rect 1034 3760 1094 4102
rect 1034 3260 1094 3700
rect 1288 3760 1348 4102
rect 1288 3694 1348 3700
rect 1376 3760 1436 4102
rect 1376 3260 1436 3700
use decoder_2to4  decoder_2to4_0
timestamp 1750825354
transform 1 0 -624 0 1 1790
box 602 -1812 2158 1470
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1704896540
transform -1 0 1119 0 -1 4079
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_1
timestamp 1704896540
transform -1 0 1468 0 -1 4079
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_2
timestamp 1704896540
transform -1 0 777 0 -1 4079
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_3
timestamp 1704896540
transform -1 0 435 0 -1 4079
box -66 -43 354 897
<< end >>
