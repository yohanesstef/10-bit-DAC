* PEX produced on Sat Jun 28 05:13:49 WIB 2025 using ./iic-pex.sh with m=2 and s=1
* NGSPICE file created from DAC_10b_top.ext - technology: sky130A

.subckt DAC_10b_posim_top DIN0 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 DIN9 ROUT1 ROUT2
+ VDD VDDH GND VOUT
X0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_45343_4538# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[1] a_6778_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X3 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_30056_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X5 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=33.8968 ps=329.23999 w=0.6 l=1
X6 a_44062_19517# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_14331_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X8 a_21927_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_23629_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1 GND sky130_fd_pr__res_xhigh_po_1p41 l=10.24
X10 a_44234_9966# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X11 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X12 a_44234_17252# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X13 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X14 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_45023_21964# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X17 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X18 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] a_43167_4358# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X20 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X22 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X23 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X24 a_14615_13536# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.VH2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X25 a_20656_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_19946_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X26 a_43698_8776# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A a_43724_9372# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X27 a_23307_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_22193_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X28 a_14948_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] a_14790_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X29 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] a_43167_3162# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB DIN2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X36 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_43240_20580# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X37 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_23307_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X38 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=11.57
X39 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X40 a_6923_9707# VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X41 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_8936# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X42 a_18284_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] a_15618_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X43 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X44 a_31042_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X45 a_36888_19550# a_36888_19786# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X46 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X47 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X48 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_24963_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X49 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[0] a_5050_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X50 a_43698_14716# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP a_43724_15312# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.99
X52 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X53 a_6923_9707# top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X54 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X55 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_21927_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X56 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_29780_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X58 a_31870_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X59 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.VL3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X60 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X61 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X62 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X63 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A a_44255_4614# GND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X64 a_23629_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.VL2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X65 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.37
X66 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X67 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT a_5050_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X68 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.087 pd=0.89 as=0.174 ps=1.78 w=0.6 l=20
X69 a_14615_14034# top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_final_switch_0.VOUT[3] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X70 a_20932_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_18724_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X71 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN a_45023_18840# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X72 a_24135_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_23629_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X73 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] a_15618_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X74 a_43167_4358# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X75 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.81
X76 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=124.854 ps=1.00292k w=1.8 l=1
X77 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] a_43391_3326# GND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X78 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X79 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X80 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X81 a_42982_21320# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_42724_21320# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X82 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X83 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_24135_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X84 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X85 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X86 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X87 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X88 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X89 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X90 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X91 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X92 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X93 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X94 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X95 a_15224_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X96 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB DIN1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X97 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 a_44234_11946# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X99 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 GND DIN2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X101 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X102 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_15629_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X103 a_31594_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X104 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 GND sky130_fd_pr__res_xhigh_po_1p41 l=6.09
X105 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] a_44255_3438# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X106 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] a_44479_3254# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X107 a_43698_9766# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_10322# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X108 a_14514_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] a_17148_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X109 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X110 GND DIN5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X111 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X112 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_14615_14034# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X113 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X114 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.45
X115 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X116 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_38672_20477# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X117 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X118 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_21375_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X119 GND DIN8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X120 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X121 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 a_16615_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X123 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_15866# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X124 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X125 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X126 a_45023_21136# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X127 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X129 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 a_33634_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_27620_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X131 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X132 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] GND GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X133 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_23629_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X134 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X135 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X136 a_43391_3878# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN a_43391_3794# GND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X137 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X139 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X140 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X141 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X142 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X143 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT a_8506_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X144 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_34304_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X145 a_5111_10963# a_5111_10963# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.464 ps=3.78 w=1.6 l=1
X146 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X147 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X148 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X149 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X151 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X152 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X153 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.58
X154 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X155 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X156 a_42724_21320# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X157 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X158 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X159 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_23859_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X160 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[2] a_8506_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X161 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X162 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_35132_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X163 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=6.65
X164 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X165 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X166 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X167 a_43240_22004# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_42982_22004# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X168 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN a_44255_3714# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X169 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X170 a_35453_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_34856_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X171 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X172 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X173 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X174 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_30608_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X175 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X176 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 a_44062_18449# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X178 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X179 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X180 GND DIN1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X181 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X182 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y a_44062_18093# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X183 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB DIN5 GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X184 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X185 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X186 VDDH top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A VOUT VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X187 a_15066_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] a_16596_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X188 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X189 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] DIN8 GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X190 a_14615_14283# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.VH2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X191 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X193 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X194 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_20823_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X195 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X196 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X198 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_14055_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X199 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X200 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.24
X201 GND top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X202 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X203 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X204 a_43240_18130# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_42982_18130# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X205 a_43240_19896# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_42982_19896# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X206 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X207 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X208 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X209 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X210 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X211 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.58
X212 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X213 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X214 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_24687_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X215 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.32
X216 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X218 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X219 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X220 a_8506_12595# top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X221 a_14672_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X222 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X223 a_35757_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_33634_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X224 a_43724_12342# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X225 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X226 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X227 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[1] a_6778_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X228 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X229 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X230 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X231 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X232 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X233 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.5
X234 a_8506_12595# VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X235 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X236 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X237 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X238 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X239 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X240 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X241 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X242 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_43240_18814# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X243 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT a_6778_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X244 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_21651_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X245 a_42847_4906# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X246 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X247 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X248 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_30332_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X249 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X250 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB a_44234_14916# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X251 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X252 a_45023_18840# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X253 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.087 ps=0.89 w=0.6 l=20
X254 a_44234_15906# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X255 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X256 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X257 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y a_44062_21653# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X258 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.88
X259 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_39936_22083# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=1
X260 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X261 a_8051_10107# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X262 a_43698_13726# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_14282# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X263 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X264 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X265 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X266 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X267 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X268 a_19468_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 top_DAC_0/top_rseg_n_dcell_0.VS4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X269 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 a_15863_13287# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 top_DAC_0/top_rseg_n_dcell_0.VH3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X271 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X272 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_final_switch_0.VOUT[0] VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X274 a_16872_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X275 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X276 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X277 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X278 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_30332_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X279 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=3.94
X280 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X281 VDD DIN9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X282 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X283 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X284 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.VS1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X285 a_39306_20477# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=5.3
X286 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X287 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X288 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X289 a_19946_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_16891_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X290 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X291 a_43724_12896# a_43698_12736# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X292 a_17732_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] a_14514_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X293 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 GND sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X294 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X295 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X296 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_15353_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X297 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X298 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_22203_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X299 GND top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X300 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.32
X301 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X302 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X303 GND a_5111_10963# a_5111_10963# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.232 ps=1.89 w=1.6 l=1
X304 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X305 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X306 a_33358_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_27344_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X307 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X308 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_20823_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X309 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X310 GND top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X311 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X312 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X313 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X314 a_8473_23194# ROUT1 ROUT1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X315 a_20076_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_19552_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X316 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_8051_10107# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X317 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X318 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.68
X319 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X320 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X321 a_44234_6996# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X322 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X323 a_8051_10107# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X324 a_44234_14282# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X325 a_34186_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_28172_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X326 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X327 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X329 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X331 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X332 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_23583_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X333 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.73
X334 a_45343_4622# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] a_45343_4538# GND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X335 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_43240_20238# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X336 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X337 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X338 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X339 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X340 a_45023_20264# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X341 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.73
X342 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X343 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X344 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X346 a_43724_9926# a_43698_9766# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X347 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_30332_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X348 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X349 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X352 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X353 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_22203_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X354 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X355 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.VL2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X356 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_21651_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X357 a_43724_16302# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X358 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 GND sky130_fd_pr__res_xhigh_po_1p41 l=6.14
X359 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X360 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X361 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X362 a_14615_13536# top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_final_switch_0.VOUT[1] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X363 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X364 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X365 a_20656_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_19468_10031# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X366 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN a_45343_3530# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X367 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X368 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X369 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_18284_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X370 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[3] a_8051_10107# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X371 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X373 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_24411_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X374 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[2] a_8506_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X375 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X376 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X377 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X378 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X379 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB a_45343_4622# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X380 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT a_8051_10107# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X381 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X382 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X383 a_43240_21320# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_42982_21320# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X384 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X385 a_38672_20477# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X386 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT a_8506_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X389 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X390 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_23031_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X391 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X392 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X393 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X396 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_final_switch_0.VOUT[3] VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X397 a_34569_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.VS1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X398 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X399 a_45023_19712# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X400 a_39306_20477# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X401 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X402 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X403 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X405 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_12896# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X406 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X407 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X408 a_6778_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X409 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.09
X411 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X412 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X413 a_44234_9332# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X414 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X415 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 a_4415_23194# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X416 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X417 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X418 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X419 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X420 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X421 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X422 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.VL2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X423 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X424 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X425 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X426 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_20547_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X427 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X428 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_45023_21136# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X429 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X430 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 GND sky130_fd_pr__res_xhigh_po_1p41 l=6.65
X431 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X432 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X433 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X434 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_30056_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X435 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X436 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X437 a_36033_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_34304_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X438 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 GND GND sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X440 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X441 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X442 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X443 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] a_43167_4634# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X444 a_43698_8776# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_9332# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X445 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X446 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X447 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_28172_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X448 a_14615_13785# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.VH2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X449 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.96
X450 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X451 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X452 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X453 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_27344_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X454 a_45023_19988# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X455 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 a_14615_13536# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X456 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_20498_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X457 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.68
X460 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X461 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X462 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X463 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_6956# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X464 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X465 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.73
X466 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.86
X467 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X468 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_5111_10963# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.232 ps=1.89 w=1.6 l=1
X469 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X470 a_16615_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X471 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X472 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_28172_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X473 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_9926# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X474 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_24963_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X475 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X476 a_36888_19550# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X477 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X478 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X479 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X480 VDD DIN6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X481 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_24411_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X482 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X483 a_36033_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_34873_10031# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X484 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB DIN4 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X485 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X486 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X487 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_21375_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X488 a_43698_15706# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP a_43724_16302# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X489 a_17443_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X490 a_44062_20941# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X491 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X492 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_43240_22004# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X493 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X494 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] DIN7 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X495 a_35177_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_35132_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X496 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X497 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] a_45023_21412# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X498 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X499 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X500 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] DIN9 GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X501 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X502 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X503 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X504 a_20222_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_17167_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X505 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_23031_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X506 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X507 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X508 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_22469_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X509 a_15224_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] a_15066_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X510 a_45343_3530# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X511 a_17732_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] a_15066_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X512 a_23629_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.VH2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X513 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_15863_13785# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X514 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X515 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[4] a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X516 a_42982_19156# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_42724_19156# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X517 GND a_36888_19786# a_36888_19550# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X518 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X519 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X520 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X521 GND top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X522 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_43240_18130# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X523 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X524 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X525 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_43240_19896# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X526 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X527 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB a_44234_11946# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X528 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X529 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X530 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X531 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X532 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X533 a_44234_12936# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X534 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X535 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_22203_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X536 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X537 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X538 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X539 a_17148_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X540 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=2.35
X541 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X542 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X543 a_43698_10756# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_11312# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X544 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.VS1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X545 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X546 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X547 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X548 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X549 a_5050_12595# top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X550 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X551 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_29780_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X553 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X554 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X555 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X556 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.94
X557 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X558 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X560 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_16856# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X561 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X562 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_20823_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X563 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X564 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X565 a_43724_10362# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X566 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X567 GND DIN4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X568 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X569 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X570 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X571 a_14948_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X572 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X573 VDD DIN0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X574 GND DIN7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X575 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X576 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X577 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X578 a_16891_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X579 a_5050_12595# VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X580 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X581 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X582 VDD DIN3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X583 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X584 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X585 a_17443_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X586 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X587 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X588 a_43167_3162# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X589 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_8051_10107# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X590 a_14672_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] a_14514_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X591 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X592 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X593 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X594 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X595 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X596 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X597 a_35453_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_34873_10031# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X598 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X599 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X600 a_42724_19156# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X601 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X602 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X603 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X604 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X605 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X606 a_44479_4254# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B a_44479_4170# GND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X607 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y a_44062_18805# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X608 VOUT top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X609 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X610 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X611 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X612 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.SH[3] a_15863_13785# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X613 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X614 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y a_44062_20229# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X615 a_16596_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X616 a_43167_4634# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X617 a_15618_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] a_14672_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X618 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X619 a_44234_11312# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X620 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X621 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT a_8051_10107# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X622 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X623 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.VH2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X624 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X625 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X626 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X627 a_21651_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_22469_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X628 a_8506_12595# VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X629 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 a_43724_7392# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X631 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X632 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_29780_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X633 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X634 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X635 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X636 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_14615_14283# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X637 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X638 a_43167_3438# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X639 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[3] a_8051_10107# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X640 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB DIN0 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X641 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X642 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_27896_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X643 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X644 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.81
X645 a_8506_12595# top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X646 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X647 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB DIN3 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X648 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 a_43724_6956# a_43698_6796# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X650 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_19670_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X651 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_30608_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X652 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X653 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X654 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 GND top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X656 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_27896_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X658 a_8473_23194# ROUT1 a_4415_23194# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X659 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB DIN6 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X660 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X661 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X662 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB DIN2 GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X663 a_43724_13332# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X664 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X665 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X666 a_44479_3254# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X667 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X668 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB a_44234_6996# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X669 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X670 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X671 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_22755_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X672 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_16181_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X673 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_27896_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X674 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X675 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X676 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X677 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.087 pd=0.89 as=0.174 ps=1.78 w=0.6 l=20
X678 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X679 a_42982_19554# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_42724_19554# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X680 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X681 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X682 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] a_43391_3878# GND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X683 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X684 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X685 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 a_17167_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X687 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X688 a_43391_3794# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] a_43391_3710# GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X689 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB a_44234_15906# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X690 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X691 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X692 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.94
X693 a_42982_20978# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_42724_20978# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X694 a_34580_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_31318_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X695 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_4415_23194# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X696 a_8051_10107# top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X697 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_24963_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X698 a_16615_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X699 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X700 a_35132_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_31870_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X701 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_8051_10107# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X702 a_43698_14716# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_15272# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X703 VOUT top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X704 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X705 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X706 a_15863_13536# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.VH3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X707 a_44062_18449# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X708 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X709 a_20352_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_20222_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X710 a_16320_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X711 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_final_switch_0.VOUT[1] VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X712 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X713 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN a_45023_19116# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X714 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X715 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X716 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X717 a_8051_10107# VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X718 a_17443_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X719 a_31594_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X720 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_15905_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X721 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X722 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=5.22
X723 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A a_42847_4906# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X724 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_23583_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X725 a_19772_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.VS4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X726 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X728 a_44255_3714# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X729 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X730 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN a_45023_20540# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X731 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X732 a_43698_9766# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A a_43724_10362# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X733 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X734 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X735 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB DIN1 GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X736 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X737 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X738 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X739 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X740 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X741 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X742 a_16891_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X743 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X744 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X745 a_43724_13886# a_43698_13726# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X746 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X747 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X748 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X749 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB a_45023_18288# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X750 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] a_43240_21320# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X751 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.63
X752 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X753 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X754 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X755 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X756 a_42847_3710# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X757 a_42724_19554# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X758 a_35453_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_33910_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X759 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 a_13779_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X760 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X761 a_20656_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_19000_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X762 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X763 a_23859_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_24209_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X764 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X765 a_16615_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X766 a_24963_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_22469_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X767 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X768 a_42724_20978# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X769 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.84
X770 a_42982_18472# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_42724_18472# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X771 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X772 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X773 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X774 a_44234_7986# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X775 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X776 a_44234_15272# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X777 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 a_14607_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X778 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X779 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X780 a_45023_19116# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X781 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X782 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 a_14948_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X784 a_44062_22009# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X785 VDDH top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X786 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X787 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X788 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X789 a_43698_6796# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A a_43724_7392# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X790 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X791 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X792 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN a_45023_18564# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X793 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X794 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X795 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 GND sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X796 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X797 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X798 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X799 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X800 a_17443_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X801 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X802 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X803 a_45023_18288# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X804 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X805 a_43724_17292# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X806 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X807 a_23307_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_24209_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X808 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X809 a_22203_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_22469_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X810 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X811 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X812 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X813 a_43698_12736# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP a_43724_13332# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X814 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X815 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X816 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_22479_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X817 a_43724_16856# a_43698_16696# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X818 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] a_44255_3162# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X819 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_18008_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X820 a_43698_6796# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_7352# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X821 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.12
X822 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X823 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X824 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] DIN9 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X825 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X826 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] GND GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X827 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_27896_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X828 a_42724_18472# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X829 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X830 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X831 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_27620_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X832 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X833 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X834 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_27620_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X835 a_37410_19098# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X836 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X837 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X838 a_43240_19156# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_42982_19156# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X839 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_21099_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X840 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A a_43391_4174# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X841 a_8506_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X842 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_22479_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X843 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X844 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X845 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X846 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.087 ps=0.89 w=0.6 l=20
X847 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X848 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X849 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_19946_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X850 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.09
X851 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X852 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X853 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X854 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X855 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X856 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X857 a_22755_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_24209_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X858 a_14790_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] a_16872_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X859 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_15353_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X860 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_27620_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X861 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X862 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X863 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X864 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X865 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X866 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_21099_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X867 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X868 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X869 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X870 a_39306_20477# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X871 a_15629_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_19000_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X872 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_27620_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X873 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X874 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_16181_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X875 a_36888_19786# a_36888_19786# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X876 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X877 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X878 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_13886# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X879 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X880 a_45023_20540# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X881 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X882 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X883 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X884 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.04
X885 a_34873_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 top_DAC_0/top_rseg_n_dcell_0.VS1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X886 a_19670_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_16615_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X887 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X888 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X889 a_39936_22083# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=1
X890 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X891 a_17167_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X892 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X893 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_15629_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X894 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X895 VDDH top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X896 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X897 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X898 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X899 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X900 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X901 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 a_15863_13287# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X902 a_20498_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_17443_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X903 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X904 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB a_44234_9966# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X905 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.SH[3] a_15863_13287# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X906 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X907 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X908 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X909 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X910 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.VH2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X911 VDDH top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A VOUT VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X912 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X913 a_14615_14283# top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_final_switch_0.VOUT[4] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X914 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X915 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X916 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X917 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X918 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_17732_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X919 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X920 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=2.5
X921 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X922 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_14615_13785# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X923 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.01
X924 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.VS1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X925 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X926 a_20547_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_23049_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X927 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.68
X928 a_34856_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_31594_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X929 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X930 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X931 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_7946# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X932 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X933 a_31042_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X934 a_17148_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X935 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X936 a_44062_21653# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X937 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X938 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X939 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X940 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.91
X941 a_45343_3978# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y a_45343_3894# GND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X942 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X943 a_31870_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X944 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X945 a_43698_16696# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP a_43724_17292# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X946 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X947 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X948 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X949 a_4415_23194# ROUT1 a_8473_23194# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X950 a_42982_21662# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_42724_21662# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X951 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X952 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y a_44062_19517# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X953 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.66
X954 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X955 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_8506_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X956 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.42
X957 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.19
X958 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.58
X959 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X960 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X961 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X962 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X963 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X964 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X965 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X966 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN a_43167_3438# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X967 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X968 a_21099_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_23049_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X969 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X970 a_43240_19554# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_42982_19554# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X971 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X972 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_23859_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X973 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X974 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X975 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X976 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X977 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_14607_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X978 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X979 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X980 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X981 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X982 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X983 a_17167_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X984 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X985 a_8506_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X986 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB a_44234_12936# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X987 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X988 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X989 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X990 a_43240_20978# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_42982_20978# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X991 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X992 a_44234_13926# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X993 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X994 a_20932_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_19670_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X995 VDDH a_5111_8388# a_5111_8388# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=0.696 ps=5.09 w=4.8 l=1
X996 GND top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B VOUT GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X997 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X998 a_43698_11746# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_12302# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X999 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_23859_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1000 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X1001 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_34856_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1002 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.VH2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1003 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_27344_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1004 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_23031_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1005 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.22
X1006 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1007 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1008 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1009 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 a_36888_19786# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1010 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0 ps=0 w=1.6 l=1
X1011 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1012 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1013 GND top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_27344_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1014 a_42724_21662# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1015 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1016 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_24687_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1017 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X1018 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1019 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1020 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1021 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1022 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1023 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1024 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_28172_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1025 a_43724_10916# a_43698_10756# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1026 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1027 a_20932_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_19772_10031# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1028 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6778_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1029 a_42982_20580# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_42724_20580# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1030 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1031 a_6923_9707# top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1032 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1033 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1034 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1035 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.01
X1036 a_15353_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_18724_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1037 a_20076_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_20498_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1038 a_5111_8388# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.696 pd=5.09 as=1.392 ps=10.18 w=4.8 l=1
X1039 a_36888_19786# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1040 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_27344_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1041 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN a_44479_3530# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1042 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1043 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_45023_21688# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1044 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1045 a_6923_9707# VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1046 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X1047 a_31318_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1048 a_16181_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_19552_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1049 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] a_44479_3898# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1050 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1051 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 GND sky130_fd_pr__res_xhigh_po_1p41 l=7.01
X1052 a_19000_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_14055_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1053 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1054 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1055 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_28172_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1056 a_16891_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1057 a_43240_18472# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_42982_18472# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1058 a_14672_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1059 a_45023_21412# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1060 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1061 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0 ps=0 w=1.6 l=1
X1062 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1063 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1064 a_44234_12302# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1065 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] a_45343_3254# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1066 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1067 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1068 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1069 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1070 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1071 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_15353_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1072 a_43724_8382# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1073 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_20222_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1074 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1075 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.VS1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1076 a_44234_16896# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1077 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1078 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.06
X1079 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1080 a_30332_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_33910_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1081 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X1082 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.89
X1083 a_44062_19161# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1084 a_20823_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_24209_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1085 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_15629_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1086 a_43724_7946# a_43698_7786# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1087 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1088 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1089 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X1090 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1091 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X1092 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1093 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=3.83
X1094 a_31042_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1095 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1096 a_15905_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_19276_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1097 a_42724_20580# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1098 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1099 a_44062_20585# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1100 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1101 a_43724_14322# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1102 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1103 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1104 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB a_44234_7986# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1105 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1106 a_8051_10107# VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1107 a_31870_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1108 a_45023_21688# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1109 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X1110 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1111 GND DIN6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1112 a_44479_3898# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1113 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1114 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1116 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1117 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB DIN4 GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1118 VDD DIN2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1119 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1120 VOUT top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1121 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1122 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1123 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1124 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0 ps=0 w=1.6 l=1
X1125 a_8051_10107# top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1126 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB a_44234_16896# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1127 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1128 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1129 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1130 a_44062_19161# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X1131 a_15224_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1132 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] DIN7 GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1133 VDD DIN5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1134 a_35757_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_34580_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1135 a_20352_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_19772_10031# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1136 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1137 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1138 a_38672_20477# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1769 pd=1.8 as=0.1769 ps=1.8 w=0.61 l=9.7
X1139 a_6778_12595# top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1140 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.6
X1141 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.17
X1142 VDD DIN8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1143 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1144 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1145 a_43698_15706# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_16262# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1146 a_43994_22522# ROUT2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X1147 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1148 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_5111_8388# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=0.696 ps=5.09 w=4.8 l=1
X1149 a_44062_20585# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X1150 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1151 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.19
X1152 GND top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1153 a_15342_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] a_16320_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1154 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1155 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A a_44479_4254# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1156 a_6778_12595# VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1157 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X1158 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_20547_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1159 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X1160 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1161 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.4
X1162 a_44479_4170# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1163 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1164 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1165 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1166 a_16891_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1167 a_44255_4614# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B a_44255_4530# GND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1168 a_43698_10756# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP a_43724_11352# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X1169 GND top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1170 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 a_15629_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1171 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_14331_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1172 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X1173 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1174 a_43724_14876# a_43698_14716# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1175 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_24411_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1176 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1177 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0 ps=0 w=1.6 l=1
X1178 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1179 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X1180 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1181 a_43391_3326# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] a_43391_3242# GND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1182 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1183 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_43240_19156# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1184 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X1185 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_10916# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1186 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1187 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1188 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_34580_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1189 a_36033_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_33358_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1190 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] a_45023_21964# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1191 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1192 a_17167_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1193 a_44234_7352# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1194 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1195 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1196 VDD DIN1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1197 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X1198 a_5111_8388# a_5111_8388# VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.696 pd=5.09 as=1.392 ps=10.18 w=4.8 l=1
X1199 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.78
X1200 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X1201 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_23049_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1202 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] a_15342_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1203 a_14615_13785# top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_final_switch_0.VOUT[2] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X1204 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB DIN5 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1205 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1206 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1207 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1208 GND DIN0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1209 a_18008_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] a_15342_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1210 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] DIN8 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1211 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1212 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X1213 a_8051_10107# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1214 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.47
X1215 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1216 a_44479_3530# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1217 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1218 a_44234_8976# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1219 GND DIN3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1220 a_44234_16262# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1221 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X1222 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1223 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1224 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_39936_22083# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9.2
X1225 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1226 a_5050_12595# VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1227 a_44062_18805# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1228 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_8506_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1229 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.37
X1230 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A a_42847_3710# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1231 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1232 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1233 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1234 a_31870_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1235 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1236 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1237 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1238 a_43698_7786# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A a_43724_8382# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X1239 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X1240 a_5050_12595# top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1241 a_42982_18814# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_42724_18814# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1242 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1243 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X1244 a_16596_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1245 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1246 a_35177_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_34186_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1247 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1248 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1249 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1250 a_18724_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_13779_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1251 a_43391_3710# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1252 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1253 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1254 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1255 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1256 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_14055_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1257 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X1258 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X1259 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1260 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.14
X1261 a_19552_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_14607_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1262 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1263 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1264 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1265 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=5.42
X1266 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1267 a_43240_21662# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_42982_21662# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1268 a_43698_13726# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP a_43724_14322# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X1269 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_final_switch_0.VOUT[4] VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X1270 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1271 a_44062_18093# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1272 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1273 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1274 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1275 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1276 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1277 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1278 a_43994_22522# ROUT2 ROUT2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X1279 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1280 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB DIN0 GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1281 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.VL3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1282 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1283 a_43698_7786# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_8342# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1284 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1285 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1286 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB DIN3 GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1287 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1288 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_20547_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1289 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1290 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_30608_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1291 a_30056_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_33634_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1292 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB DIN6 GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1293 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X1294 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X1295 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1296 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT a_5050_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1297 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1298 a_20352_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_19276_8950# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1299 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1300 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1301 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1302 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1303 a_31594_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1304 a_34304_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_31042_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1305 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1306 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1307 a_16872_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1308 ROUT1 ROUT1 a_8473_23194# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X1309 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[0] a_5050_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1310 a_42724_18814# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1311 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1312 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3 GND sky130_fd_pr__res_xhigh_po_1p41 l=8.5
X1313 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_23307_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1314 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_30332_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1315 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1316 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1317 a_44234_10956# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1318 a_18284_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] a_15066_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1319 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1320 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X1321 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1322 a_14615_14034# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.VH2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1323 a_37410_19098# a_37410_19098# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1856 pd=1.86 as=0.1856 ps=1.86 w=0.64 l=12
X1324 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.32
X1325 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1326 a_44062_20229# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1327 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1328 a_44255_4162# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] a_44255_4078# GND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1329 a_31318_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1330 a_22755_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_22193_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1331 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1332 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC a_37410_19098# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1333 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_21927_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1334 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.464 pd=3.78 as=0.464 ps=3.78 w=1.6 l=1
X1335 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.94
X1336 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1337 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_43240_19554# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1338 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1339 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1340 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_14876# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1341 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_21375_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1342 a_44255_4530# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C a_44255_4446# GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1343 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1344 a_42982_20238# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_42724_20238# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1345 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X1346 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1347 a_4415_23194# a_4415_23194# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=20
X1348 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.27
X1349 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1350 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] a_43240_20978# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1351 a_43391_3242# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB a_43391_3158# GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1352 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_15863_13536# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X1353 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1354 a_45023_18564# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1355 a_43240_20580# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_42982_20580# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1356 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1357 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1358 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 a_15353_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1359 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X1360 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_14055_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1361 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB a_44234_10956# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1362 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1363 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1364 GND a_36888_19786# a_36888_19786# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1365 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1366 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1367 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[4] a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1368 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1369 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 a_16181_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1370 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1371 GND top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X1372 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1373 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1374 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.VS1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1375 a_43994_22522# ROUT2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X1376 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 a_14331_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1377 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_22755_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1378 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1379 a_18008_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] a_14790_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1380 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB a_44255_4162# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1381 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1382 a_44255_3162# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1383 a_6778_12595# VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1384 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN a_45023_19988# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1385 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1386 a_44255_4078# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1388 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1389 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X1390 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1391 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1392 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1393 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_16181_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1394 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1395 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1396 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1397 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1 GND sky130_fd_pr__res_xhigh_po_1p41 l=11.57
X1398 a_44255_4446# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1399 a_6778_12595# top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1400 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1401 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1402 a_43391_4174# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1403 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X1404 a_42724_20238# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1405 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1406 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X1407 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1408 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 GND sky130_fd_pr__res_xhigh_po_1p41 l=7.88
X1409 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.83
X1410 a_31594_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1411 a_43391_3158# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1412 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_43240_18472# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1413 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1414 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1415 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 GND sky130_fd_pr__res_xhigh_po_1p41 l=5.47
X1416 a_43724_11352# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1417 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X1418 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1419 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1420 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X1421 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1422 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_23307_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1423 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1424 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1425 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1426 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_13779_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1427 a_44255_3438# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1428 top_DAC_0/top_final_switch_0.VOUT[3] top_DAC_0/top_rseg_n_dcell_0.SH[3] a_15863_13536# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1429 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] a_45023_20264# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1430 a_44234_10322# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1431 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1432 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1433 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.63
X1434 a_19276_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_14331_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1435 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1436 GND top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B VOUT GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1437 a_24209_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.VL2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1438 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1439 a_23031_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_23049_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1440 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1441 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1442 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1443 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=3.17
X1444 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1445 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB a_44234_13926# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1446 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_14607_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1447 a_44234_14916# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1448 a_44062_19873# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1449 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_21927_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1450 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_4415_23194# a_4415_23194# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=20
X1451 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1452 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1453 a_31318_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1454 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1455 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1456 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] a_29780_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1457 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1458 a_43698_12736# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_13292# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1459 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1460 a_29780_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_33358_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1463 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_13779_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1464 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1465 GND top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1466 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X1467 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X1468 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_24687_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1469 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1470 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1471 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1472 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1473 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X1474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1475 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_24135_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1476 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X1477 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1478 a_30608_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_34186_8950# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1479 a_35757_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_34569_10031# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1480 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_14607_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1481 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1482 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_21099_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1483 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_15905_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1484 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 GND sky130_fd_pr__res_xhigh_po_1p41 l=3.53
X1485 GND top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X1486 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_30056_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1487 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_8051_10107# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1488 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1489 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1490 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1491 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1492 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1493 a_44062_19873# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X1494 a_43724_11906# a_43698_11746# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1495 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1496 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1497 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_14331_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1498 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1499 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1500 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1501 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1502 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_22755_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1503 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X1504 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1505 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1506 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1507 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X1508 a_45343_3894# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1509 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X1510 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1511 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1512 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1513 a_42982_22004# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_42724_22004# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1514 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.35
X1515 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1516 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1517 a_8051_10107# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1518 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1519 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.232 ps=1.89 w=1.6 l=1
X1520 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1521 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1522 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] a_45023_19712# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1523 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X1524 a_44234_13292# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1525 a_31318_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1526 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1527 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X1528 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1529 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1530 VOUT top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X1531 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1532 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1533 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_13779_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1534 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1535 a_43724_9372# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1536 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1537 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1538 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=1.392 pd=10.18 as=1.392 ps=10.18 w=4.8 l=1
X1539 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3 GND sky130_fd_pr__res_xhigh_po_1p41 l=9.22
X1540 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1541 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_24135_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1542 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X1543 a_43240_18814# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_42982_18814# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1544 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1545 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 a_15905_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1546 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_23583_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1547 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_30608_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1548 a_15863_13785# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.VH3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.0609 pd=0.71 as=0.1218 ps=1.42 w=0.42 l=0.5
X1549 a_44062_21297# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1550 a_42982_18130# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_42724_18130# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1551 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1552 a_42982_19896# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_42724_19896# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1553 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_final_switch_0.VOUT[2] VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X1554 a_43724_8936# a_43698_8776# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1555 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X1556 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y a_44062_20941# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X1557 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 a_14055_6250# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1558 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 GND sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X1559 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1560 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1561 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1562 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1563 a_20823_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_22193_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1564 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1565 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1566 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1567 a_43724_15312# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1568 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_5050_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1569 GND top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB a_44234_8976# GND sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1570 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X1571 a_5050_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1572 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1573 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_final_switch_0.VOUT[0] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.0609 ps=0.71 w=0.42 l=0.5
X1574 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1575 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_15905_7686# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1576 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1577 a_35177_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_34569_10031# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1578 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1579 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1580 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1581 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 a_36888_19550# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1582 a_42724_22004# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1583 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y a_45343_3978# GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1584 a_44062_22009# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1585 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1586 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1587 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1588 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1589 a_44062_21297# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X1590 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1591 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X1592 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1593 a_20076_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_19468_10031# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1594 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1595 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1596 a_43698_16696# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_17252# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1597 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_21651_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1598 a_16320_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1599 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1600 VDD DIN4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1601 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_18008_18696# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1602 a_5111_10963# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.232 pd=1.89 as=0.464 ps=3.78 w=1.6 l=1
X1603 a_33910_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_27896_6250# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1604 a_22479_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_23629_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1605 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1606 VDD DIN7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1607 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] a_43240_21662# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1608 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1609 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X1610 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1611 a_21375_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_22193_18133# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1612 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X1613 GND DIN9 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] GND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1614 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1615 GND GND GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0 ps=0 w=0.6 l=1
X1616 a_42724_18130# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1617 GND GND sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1618 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_30056_7686# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1619 a_42724_19896# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1620 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 GND sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X1621 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X1622 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1623 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1624 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1625 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1626 a_43698_11746# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP a_43724_12342# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X1627 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1628 a_43994_22522# ROUT2 ROUT2 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X1629 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 GND sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1630 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1631 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1632 a_43724_15866# a_43698_15706# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1633 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1634 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1635 a_31042_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1636 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1637 a_45343_3254# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] GND GND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1638 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT a_6778_12595# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1639 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1640 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 GND sky130_fd_pr__res_xhigh_po_1p41 l=7.42
X1641 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1642 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_11906# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X1643 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6923_9707# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1644 a_43240_20238# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_42982_20238# VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1645 GND GND GND sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X1646 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1647 VDDH VDDH VDDH VDDH sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1648 a_44234_8342# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN GND GND sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1649 GND top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1650 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X1651 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_22479_20174# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1652 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
C0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.08365f
C1 top_DAC_0/top_rseg_n_dcell_0.VH2 a_23629_18133# 0.26291f
C2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_17443_7686# 0.18047f
C3 a_19276_8950# a_20352_10031# 0.03999f
C4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 1.15809f
C5 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.03925f
C6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.10923f
C7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_31318_7686# 0.11573f
C8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15224_18696# 0.11194f
C9 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.02784f
C10 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.16417f
C11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 a_21375_20174# 0.0516f
C12 a_23629_18133# a_22479_20174# 0.04085f
C13 a_24209_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.42807f
C14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 1.26125f
C15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 0.04506f
C16 a_17148_18696# a_14514_18696# 0.04589f
C17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 0.05522f
C18 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_6923_9707# 0.05319f
C19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 a_28172_6250# 0.03309f
C20 a_15353_7686# a_18724_8950# 0.03934f
C21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.06177f
C22 VDDH a_16596_18696# 0.28004f
C23 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 a_29158_6250# 0.05085f
C24 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 8.67322f
C25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.30645f
C26 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_13332# 0.03597f
C27 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 a_28882_6250# 0.0856f
C28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 a_28606_6250# 0.03285f
C29 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 a_21099_20174# 0.05515f
C30 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.13554f
C31 a_34186_8950# a_35132_8950# 0.1022f
C32 a_34304_8950# a_34856_8950# 0.09199f
C33 VOUT a_8506_12595# 0.46012f
C34 a_31042_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.03929f
C35 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.05693f
C36 a_30332_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.07404f
C37 DIN5 VDD 0.67364f
C38 VDDH a_43724_17292# 0.09226f
C39 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.04419f
C40 a_15353_7686# a_14607_6250# 0.05354f
C41 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 a_15224_18696# 0.05173f
C42 a_15629_7686# a_14331_6250# 0.02789f
C43 a_15905_7686# a_14055_6250# 0.02786f
C44 a_15869_6250# a_15041_6250# 0.18522f
C45 a_39883_19479# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.02736f
C46 a_16181_7686# a_13779_6250# 0.03169f
C47 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_14916# 0.03855f
C48 a_31318_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.02708f
C49 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.28651f
C50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 1.33058f
C51 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.92839f
C52 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_final_switch_0.VOUT[1] 0.01859f
C53 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.0394f
C54 a_14615_14283# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.1083f
C55 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 0.53808f
C56 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 0.02066f
C57 a_39768_20665# a_39768_20389# 0.02286f
C58 a_14615_13785# a_14615_13536# 0.1195f
C59 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_2678_22970# 0.07653f
C60 a_14790_18696# a_15342_18696# 0.08353f
C61 a_14514_18696# a_15618_18696# 0.10675f
C62 a_24135_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 0.06476f
C63 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB a_44234_15906# 0.08412f
C64 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] VDDH 2.21503f
C65 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] VDDH 0.88599f
C66 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 0.07805f
C67 a_33358_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.02254f
C68 a_35177_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.15755f
C69 top_DAC_0/top_final_switch_0.VOUT[0] a_14615_13536# 0.09871f
C70 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.04328f
C71 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.06351f
C72 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.15973f
C73 a_24687_20174# a_21651_20174# 0.13223f
C74 a_24963_20174# a_21375_20174# 0.14448f
C75 a_29780_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.11538f
C76 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.07764f
C77 a_16181_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.0776f
C78 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 0.06384f
C79 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 a_13779_6250# 0.04915f
C80 a_22193_18133# a_23049_18133# 0.19287f
C81 top_DAC_0/top_rseg_n_dcell_0.VL2 a_22469_18133# 0.5366f
C82 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.03029f
C83 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.03617f
C84 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 a_13779_6250# 0.04304f
C85 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.VS4 0.03086f
C86 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.14571f
C87 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_28882_6250# 0.34979f
C88 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 1.79255f
C89 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_15629_7686# 0.08674f
C90 VDDH a_19552_8950# 0.27813f
C91 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 1.33533f
C92 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 a_21927_20174# 0.04145f
C93 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_20547_20174# 0.15594f
C94 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.04269f
C95 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.02791f
C96 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.11852f
C97 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 VDDH 0.24469f
C98 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 3.28115f
C99 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.15933f
C100 a_22469_18133# a_23629_18133# 0.1849f
C101 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15041_6250# 0.14352f
C102 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.23291f
C103 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] VDDH 0.01029f
C104 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.0686f
C105 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.06598f
C106 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 a_27896_6250# 0.02786f
C107 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 a_27344_6250# 0.13824f
C108 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.18677f
C109 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 1.09015f
C110 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 0.12088f
C111 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 0.25126f
C112 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.29164f
C113 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.21785f
C114 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.57519f
C115 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.3441f
C116 a_1636_13708# VOUT 0.0165f
C117 a_43698_9766# a_43724_10362# 0.06762f
C118 a_29158_6250# a_31318_7686# 0.02794f
C119 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 a_22479_20174# 0.0849f
C120 a_30056_7686# a_30332_7686# 6.43201f
C121 a_28606_6250# a_31870_7686# 0.23705f
C122 a_28882_6250# a_31594_7686# 0.02807f
C123 a_29434_6250# a_31042_7686# 0.03864f
C124 a_29780_7686# a_30608_7686# 0.20841f
C125 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.02665f
C126 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.09657f
C127 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 1.48f
C128 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_9901_14150# 0.04994f
C129 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.0759f
C130 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 0.04946f
C131 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 1.96915f
C132 a_24687_20174# a_23031_20174# 4.95717f
C133 a_24963_20174# a_22755_20174# 4.63841f
C134 a_24411_20174# a_23307_20174# 5.3026f
C135 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.08345f
C136 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 9.03926f
C137 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 0.0119f
C138 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_20222_8950# 0.19554f
C139 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 1.68518f
C140 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP a_44234_12936# 0.06668f
C141 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.09979f
C142 a_24135_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1 0.04143f
C143 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 0.02159f
C144 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C145 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 0.06186f
C146 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.33336f
C147 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 0.06502f
C148 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 1.68908f
C149 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 0.02084f
C150 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_27896_6250# 0.21279f
C151 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_21927_20174# 0.17166f
C152 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_44062_19161# 0.02354f
C153 a_35132_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.11604f
C154 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_15593_6250# 0.14732f
C155 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04402f
C156 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.28898f
C157 top_DAC_0/top_final_switch_0.VOUT[2] a_9353_12507# 0.01061f
C158 a_16891_7686# a_17167_7686# 6.30798f
C159 a_16615_7686# a_17443_7686# 0.17805f
C160 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.01105f
C161 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 1.40678f
C162 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 0.10118f
C163 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.22711f
C164 VDDH top_DAC_0/top_final_switch_0.VOUT[4] 2.1005f
C165 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] a_16320_18696# 0.11863f
C166 a_17148_18696# a_16596_18696# 0.10042f
C167 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.55413f
C168 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_28172_6250# 0.16633f
C169 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 VDDH 0.14565f
C170 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 a_14948_18696# 0.05505f
C171 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 0.20475f
C172 a_35453_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.04964f
C173 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.03943f
C174 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB VDD 0.63982f
C175 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 a_15869_6250# 0.04387f
C176 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.16758f
C177 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.30168f
C178 a_19468_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.26189f
C179 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.11561f
C180 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C VDD 0.26024f
C181 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09914f
C182 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.08642f
C183 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 1.01892f
C184 top_DAC_0/top_rseg_n_dcell_0.VH2 a_14615_14283# 0.15488f
C185 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_20547_20174# 0.24099f
C186 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 0.16142f
C187 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.26598f
C188 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.02242f
C189 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_14615_14034# 0.09164f
C190 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.05169f
C191 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.27586f
C192 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.09063f
C193 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_17148_18696# 0.22491f
C194 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 1.54537f
C195 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.05346f
C196 a_5897_15057# VOUT 0.04644f
C197 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.12876f
C198 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 a_27344_6250# 0.05089f
C199 a_23583_20174# a_24687_20174# 0.29545f
C200 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[2] 0.59509f
C201 a_23859_20174# a_24411_20174# 0.15434f
C202 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.0127f
C203 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.04506f
C204 a_23049_18133# a_24963_20174# 0.06769f
C205 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 a_28882_6250# 0.02795f
C206 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.13628f
C207 a_15629_7686# a_15905_7686# 6.27398f
C208 a_15353_7686# a_16181_7686# 0.20823f
C209 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.27678f
C210 a_43698_13726# a_43724_13886# 0.02395f
C211 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 a_22203_20174# 0.04143f
C212 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.VS1 0.07652f
C213 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.1278f
C214 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP a_44234_13926# 0.06668f
C215 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.25101f
C216 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 0.08832f
C217 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y VDD 0.49613f
C218 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.40887f
C219 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 a_27620_6250# 0.07802f
C220 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.02797f
C221 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_17732_18696# 0.14577f
C222 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.11776f
C223 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.18541f
C224 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 0.04506f
C225 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02493f
C226 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 0.0126f
C227 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 1.21429f
C228 a_31318_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.06185f
C229 a_24135_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 0.04172f
C230 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.04541f
C231 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.05696f
C232 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_15618_18696# 0.05915f
C233 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 0.05431f
C234 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP a_44234_15906# 0.06668f
C235 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.06862f
C236 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 a_15353_7686# 0.04539f
C237 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_21927_20174# 0.17476f
C238 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.08705f
C239 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.11848f
C240 a_14055_6250# a_17443_7686# 0.04961f
C241 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_14916# 0.14379f
C242 a_14331_6250# a_17167_7686# 0.02801f
C243 a_15041_6250# a_16615_7686# 0.04051f
C244 a_14607_6250# a_16891_7686# 0.04273f
C245 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_27896_6250# 0.15674f
C246 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 1.94958f
C247 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 0.08427f
C248 a_11081_12507# top_DAC_0/top_final_switch_0.VOUT[3] 0.01061f
C249 a_8173_15057# top_DAC_0/top_final_switch_0.VOUT[2] 0.03029f
C250 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 0.3076f
C251 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.02785f
C252 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.05433f
C253 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.11409f
C254 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.02595f
C255 a_43698_12736# a_44234_13292# 0.07082f
C256 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_34873_10031# 0.15163f
C257 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 a_17167_7686# 0.03929f
C258 a_28172_6250# a_29158_6250# 0.1647f
C259 a_28606_6250# a_28882_6250# 8.21854f
C260 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.02791f
C261 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 a_8051_10107# 0.5084f
C262 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.02873f
C263 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.85005f
C264 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04883f
C265 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 a_13779_6250# 0.04328f
C266 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.18998f
C267 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 1.96543f
C268 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 0.1298f
C269 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.1111f
C270 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 0.61284f
C271 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04929f
C272 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_17167_7686# 0.07921f
C273 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.08564f
C274 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.82224f
C275 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 0.09131f
C276 a_31042_7686# a_27620_6250# 0.02789f
C277 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.02015f
C278 a_30608_7686# a_27896_6250# 0.02792f
C279 a_31318_7686# a_27344_6250# 0.03762f
C280 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 a_15593_6250# 0.04474f
C281 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 23.5069f
C282 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.03749f
C283 a_20932_10031# a_18724_8950# 0.0898f
C284 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_15863_13536# 0.04948f
C285 a_36813_19462# a_36888_19786# 0.03172f
C286 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 0.03971f
C287 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.15048f
C288 a_20656_10031# a_19000_8950# 0.03997f
C289 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_44062_19161# 0.06327f
C290 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.23412f
C291 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_9901_12507# 0.02171f
C292 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.03925f
C293 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 0.12176f
C294 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_20656_10031# 0.27487f
C295 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.50346f
C296 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.09135f
C297 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.15123f
C298 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_21375_20174# 0.20734f
C299 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.04382f
C300 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.56698f
C301 a_14055_6250# a_19000_8950# 0.03929f
C302 a_31870_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.03966f
C303 a_44234_11312# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.02704f
C304 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN VDD 0.3628f
C305 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 0.14746f
C306 VDDH a_2678_16243# 0.72648f
C307 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 1.8611f
C308 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.1591f
C309 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 0.52808f
C310 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 0.05143f
C311 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.15088f
C312 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.48636f
C313 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 a_16891_7686# 0.07402f
C314 a_15374_19866# a_16596_18696# 0.0884f
C315 a_15098_19866# a_16872_18696# 0.10119f
C316 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.03934f
C317 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.09294f
C318 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_final_switch_0.VOUT[4] 0.06373f
C319 a_2678_19053# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 0.05235f
C320 a_44234_7352# a_44234_6996# 0.08026f
C321 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_38584_20665# 0.01092f
C322 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.4374f
C323 a_14331_6250# a_14607_6250# 7.49126f
C324 a_14055_6250# a_15041_6250# 0.17838f
C325 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05451f
C326 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.02163f
C327 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.11848f
C328 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.27905f
C329 a_15066_18696# VDDH 0.31303f
C330 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A VDD 0.35622f
C331 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04788f
C332 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.17902f
C333 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.15992f
C334 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 a_37804_20713# 0.03421f
C335 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] a_14672_18696# 0.03073f
C336 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 a_29434_6250# 0.03934f
C337 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.0184f
C338 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 a_14607_6250# 0.02789f
C339 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_18724_8950# 0.0657f
C340 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.0494f
C341 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 a_15593_6250# 0.02795f
C342 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.04365f
C343 a_37595_19462# a_37737_19479# 0.04234f
C344 a_4978_9535# a_5642_9535# 0.02543f
C345 a_19468_10031# VDDH 0.17518f
C346 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 4.7892f
C347 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_15374_19866# 0.17301f
C348 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_19946_8950# 0.03391f
C349 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_6956# 0.03597f
C350 a_43698_10756# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.24498f
C351 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.07852f
C352 VDDH a_43724_16302# 0.09227f
C353 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.07479f
C354 VDDH ROUT1 29.7603f
C355 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.VL3 0.1844f
C356 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.10293f
C357 a_34186_8950# a_30608_7686# 0.03938f
C358 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 0.04812f
C359 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.05872f
C360 a_43724_11352# a_43698_10756# 0.06762f
C361 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_22755_20174# 0.02888f
C362 a_15618_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.22383f
C363 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC ROUT2 0.01108f
C364 a_43698_15706# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.7858f
C365 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_14607_6250# 0.15518f
C366 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 2.73645f
C367 a_44234_9332# a_44234_9966# 0.02262f
C368 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 1.97694f
C369 VDDH top_DAC_0/top_rseg_n_dcell_0.SH[3] 1.2895f
C370 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.08366f
C371 a_43724_11352# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.03597f
C372 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 0.01178f
C373 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 0.03841f
C374 a_1896_17510# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 0.03145f
C375 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 2.01068f
C376 a_43698_8776# a_43724_9372# 0.06762f
C377 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B VDD 0.36582f
C378 a_44234_12302# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.08412f
C379 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.01814f
C380 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 0.2138f
C381 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 2.48553f
C382 a_44062_21297# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.09819f
C383 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.08425f
C384 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.13405f
C385 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_15869_6250# 0.30978f
C386 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.36581f
C387 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_final_switch_0.VOUT[0] 0.0151f
C388 a_16181_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 0.0808f
C389 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 2.35144f
C390 a_16891_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.07419f
C391 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.19658f
C392 a_17443_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.0394f
C393 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_20823_20174# 0.11552f
C394 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.14199f
C395 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.25378f
C396 a_15905_7686# a_17167_7686# 0.16165f
C397 a_16181_7686# a_16891_7686# 0.16678f
C398 a_15629_7686# a_17443_7686# 0.17897f
C399 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.15057f
C400 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 0.86006f
C401 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 a_28606_6250# 0.03927f
C402 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 a_14607_6250# 0.02784f
C403 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.01174f
C404 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.02352f
C405 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.0935f
C406 DIN4 VDDH 0.42749f
C407 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_23629_18133# 0.25057f
C408 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 VDDH 0.11991f
C409 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B VDD 0.25878f
C410 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6778_12595# 0.8028f
C411 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.04187f
C412 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.11031f
C413 a_5111_8388# a_5642_9535# 0.03284f
C414 VDDH a_11629_14150# 0.49013f
C415 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.14066f
C416 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_13779_6250# 1.293f
C417 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.11523f
C418 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04362f
C419 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 0.16406f
C420 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.10029f
C421 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_37022_20295# 0.01181f
C422 a_28172_6250# a_27344_6250# 0.33712f
C423 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 1.40088f
C424 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_12936# 0.03152f
C425 a_44062_20941# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.06327f
C426 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 0.04508f
C427 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.37208f
C428 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 1.32603f
C429 a_43698_13726# a_43698_14716# 0.01563f
C430 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 0.02497f
C431 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.36573f
C432 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.06309f
C433 a_44062_19873# a_44062_19517# 0.04238f
C434 a_22193_18133# a_23307_20174# 0.09185f
C435 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.01069f
C436 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.02757f
C437 a_35177_10031# a_35453_10031# 1.72453f
C438 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.11733f
C439 a_34873_10031# a_35757_10031# 0.35722f
C440 a_19670_8950# a_20222_8950# 0.09199f
C441 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.09312f
C442 VDDH a_7625_14150# 0.49013f
C443 a_1896_22970# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.06357f
C444 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.0938f
C445 a_19552_8950# a_20498_8950# 0.10162f
C446 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN a_44234_16262# 0.08412f
C447 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04799f
C448 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 a_5050_12595# 0.20391f
C449 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_22203_20174# 0.12118f
C450 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.33091f
C451 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 16.8068f
C452 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.11409f
C453 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09099f
C454 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y a_44062_19517# 0.07788f
C455 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 a_14055_6250# 0.02787f
C456 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.16197f
C457 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.08427f
C458 a_8051_10107# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.55166f
C459 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 2.0142f
C460 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.12637f
C461 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_31870_7686# 0.20287f
C462 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.02784f
C463 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_14672_18696# 0.12567f
C464 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 1.85343f
C465 a_44062_21297# a_44062_20941# 0.04238f
C466 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.19471f
C467 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 0.56552f
C468 a_23629_18133# a_23031_20174# 0.06781f
C469 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.09623f
C470 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 4.12073f
C471 a_15629_7686# a_19000_8950# 0.03932f
C472 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.11409f
C473 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 0.64103f
C474 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 a_28882_6250# 0.02796f
C475 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.14065f
C476 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_2678_19053# 0.06357f
C477 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.01854f
C478 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 a_29780_7686# 0.04526f
C479 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.02794f
C480 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.05594f
C481 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 0.05832f
C482 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 a_29158_6250# 0.02797f
C483 top_DAC_0/top_final_switch_0.VOUT[0] a_5050_12595# 0.47498f
C484 a_34580_8950# a_35132_8950# 0.10459f
C485 a_14331_6250# a_19276_8950# 0.03929f
C486 VOUT a_8173_12507# 0.03463f
C487 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.158f
C488 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.02788f
C489 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 0.0543f
C490 DIN4 DIN5 0.34355f
C491 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.11771f
C492 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.0973f
C493 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_8506_12595# 0.51626f
C494 a_1636_15118# a_1636_14353# 0.02286f
C495 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.04069f
C496 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.61579f
C497 top_DAC_0/top_rseg_n_dcell_0.VS1 a_20076_10031# 0.09814f
C498 a_15905_7686# a_14607_6250# 0.0413f
C499 a_15629_7686# a_15041_6250# 0.0383f
C500 a_16181_7686# a_14331_6250# 0.02791f
C501 a_31870_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.02521f
C502 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.05719f
C503 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.0119f
C504 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09272f
C505 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_17510# 0.06384f
C506 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 1.97317f
C507 a_43698_12736# a_43698_13726# 0.01563f
C508 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN a_44234_8976# 0.06923f
C509 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 4.37057f
C510 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 1.52401f
C511 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_2678_21703# 0.01199f
C512 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.0517f
C513 a_15066_18696# a_15618_18696# 0.09456f
C514 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.02523f
C515 a_35757_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.27766f
C516 top_DAC_0/top_final_switch_0.VOUT[2] a_9353_15057# 0.03805f
C517 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 a_30332_7686# 0.07456f
C518 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.02786f
C519 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.63882f
C520 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 0.77088f
C521 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_final_switch_0.VOUT[1] 0.01878f
C522 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 a_6923_9707# 0.02693f
C523 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN VDD 6.73678f
C524 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_19276_8950# 0.0735f
C525 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 0.1237f
C526 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] a_45015_4828# 0.02963f
C527 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.65418f
C528 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.04529f
C529 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 a_14331_6250# 0.02786f
C530 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 1.41253f
C531 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 a_14331_6250# 0.03524f
C532 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.0436f
C533 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.02165f
C534 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 1.7882f
C535 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 0.17104f
C536 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 0.04735f
C537 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_29434_6250# 0.52669f
C538 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 0.02201f
C539 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_16181_7686# 0.08174f
C540 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 1.55513f
C541 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP 0.10923f
C542 VDDH a_19946_8950# 0.2909f
C543 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.11127f
C544 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_36888_19786# 0.03571f
C545 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 a_21651_20174# 0.04143f
C546 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 3.83937f
C547 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.04211f
C548 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_21099_20174# 0.16779f
C549 a_6923_9707# a_6778_12595# 0.02789f
C550 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.04267f
C551 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.11006f
C552 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.13075f
C553 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.16722f
C554 a_4415_23194# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 6.32681f
C555 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04799f
C556 a_23583_20174# a_23629_18133# 0.06767f
C557 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.1484f
C558 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y a_45023_18288# 0.01032f
C559 VDDH a_2300_15118# 0.54014f
C560 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 a_27896_6250# 0.04376f
C561 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.24146f
C562 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 a_17148_18696# 0.04033f
C563 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_1896_16243# 0.08441f
C564 a_43698_9766# a_44234_9966# 0.0139f
C565 a_24963_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 0.04143f
C566 a_29780_7686# a_31318_7686# 0.20433f
C567 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.01138f
C568 a_29434_6250# a_31594_7686# 0.03867f
C569 a_30056_7686# a_31042_7686# 0.16668f
C570 a_29158_6250# a_31870_7686# 0.05007f
C571 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 0.1048f
C572 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.04684f
C573 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.09942f
C574 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.VL3 0.06485f
C575 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 0.98571f
C576 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_8506_12595# 0.55664f
C577 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 0.01848f
C578 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 a_28172_6250# 0.04365f
C579 a_24963_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 0.08491f
C580 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.VH3 0.13103f
C581 a_30332_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.03985f
C582 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 a_13779_6250# 0.22304f
C583 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 a_23307_20174# 0.06393f
C584 a_24963_20174# a_23307_20174# 0.17068f
C585 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C586 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 1.15763f
C587 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_38617_19854# 0.02826f
C588 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.19276f
C589 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.71703f
C590 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.32264f
C591 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 0.33228f
C592 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.06127f
C593 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 0.24606f
C594 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.07915f
C595 a_31594_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 0.03976f
C596 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 1.34308f
C597 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_2678_21703# 0.13435f
C598 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 1.05222f
C599 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_16615_7686# 0.12435f
C600 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.14205f
C601 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_6996# 0.01131f
C602 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.12585f
C603 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_22479_20174# 0.17903f
C604 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_15353_7686# 0.49839f
C605 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_11629_14150# 0.04994f
C606 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.11775f
C607 a_43698_12736# a_43724_12896# 0.02395f
C608 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.01045f
C609 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 2.20196f
C610 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 0.05218f
C611 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 0.0549f
C612 a_23859_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 0.05527f
C613 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.02213f
C614 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.0142f
C615 a_17167_7686# a_17443_7686# 6.41047f
C616 a_35177_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.23822f
C617 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 3.4847f
C618 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] a_16872_18696# 0.13882f
C619 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.18829f
C620 a_43698_10756# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.02387f
C621 a_31870_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.0394f
C622 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 a_20823_20174# 0.06393f
C623 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.01032f
C624 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_28882_6250# 0.24414f
C625 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_7625_14150# 0.04959f
C626 a_36033_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.07439f
C627 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.29779f
C628 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 0.02179f
C629 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 a_15629_7686# 0.04025f
C630 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 a_14615_13785# 0.07377f
C631 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.0839f
C632 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.04736f
C633 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_5642_9535# 0.01613f
C634 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 0.14118f
C635 top_DAC_0/top_rseg_n_dcell_0.VH2 a_14615_13785# 0.11752f
C636 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.02784f
C637 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 0.0174f
C638 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.0596f
C639 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_21099_20174# 0.17158f
C640 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.05371f
C641 a_15098_19866# a_15342_18696# 0.01348f
C642 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.0923f
C643 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 a_21651_20174# 0.04143f
C644 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 a_13779_6250# 0.08114f
C645 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_final_switch_0.VOUT[0] 0.01053f
C646 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.01196f
C647 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.01074f
C648 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.14539f
C649 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.20862f
C650 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.04885f
C651 a_15905_7686# a_19276_8950# 0.03932f
C652 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 0.0518f
C653 a_5897_14150# VOUT 0.06743f
C654 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 0.04791f
C655 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.11097f
C656 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.1675f
C657 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 a_27896_6250# 0.03699f
C658 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 2.40428f
C659 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.09596f
C660 a_2678_20320# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.01554f
C661 a_24135_20174# a_24687_20174# 0.22999f
C662 a_23859_20174# a_24963_20174# 0.32655f
C663 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 a_27344_6250# 0.08425f
C664 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 1.18645f
C665 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 1.77943f
C666 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 a_29434_6250# 0.04713f
C667 a_15905_7686# a_16181_7686# 6.22879f
C668 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.09312f
C669 a_5050_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.02955f
C670 a_14514_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.53077f
C671 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05095f
C672 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.17777f
C673 a_20547_20174# a_20823_20174# 1.13177f
C674 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.10008f
C675 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 0.12879f
C676 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.21439f
C677 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.03135f
C678 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 14.0478f
C679 a_14615_14034# top_DAC_0/top_final_switch_0.VOUT[3] 0.10128f
C680 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_5642_10963# 0.0541f
C681 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_8051_10107# 3.25971f
C682 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.01392f
C683 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_18284_18696# 0.12145f
C684 a_33634_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.02723f
C685 a_17443_7686# a_18724_8950# 0.17302f
C686 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.10421f
C687 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.06993f
C688 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 0.32254f
C689 a_6778_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 0.12565f
C690 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.01392f
C691 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.3835f
C692 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 1.85532f
C693 a_15629_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.04025f
C694 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_14055_6250# 0.17048f
C695 a_31870_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.26664f
C696 a_44234_8976# a_44234_8342# 0.02262f
C697 a_43698_15706# a_43724_16302# 0.06762f
C698 a_44234_7352# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.06548f
C699 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.07957f
C700 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.96812f
C701 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.07627f
C702 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.35307f
C703 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP 0.01782f
C704 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.18597f
C705 DIN5 VDDH 0.42749f
C706 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 0.02199f
C707 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_22479_20174# 0.19488f
C708 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 a_15905_7686# 0.03985f
C709 a_14607_6250# a_17443_7686# 0.12868f
C710 a_15041_6250# a_17167_7686# 0.05985f
C711 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 1.14685f
C712 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_27620_6250# 0.15597f
C713 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.44826f
C714 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.29614f
C715 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.46012f
C716 a_43724_17292# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.03147f
C717 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_35453_10031# 0.12639f
C718 a_44234_17252# a_43698_16696# 0.07082f
C719 a_39768_20665# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.03153f
C720 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.08366f
C721 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_final_switch_0.VOUT[2] 0.01031f
C722 a_28606_6250# a_29434_6250# 0.19193f
C723 a_28172_6250# a_29780_7686# 0.05609f
C724 a_28882_6250# a_29158_6250# 7.83144f
C725 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.05128f
C726 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 0.08969f
C727 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.02803f
C728 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.44079f
C729 a_20823_20174# a_21927_20174# 5.19083f
C730 a_20547_20174# a_22203_20174# 4.80072f
C731 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_13292# 0.03855f
C732 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.05175f
C733 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 a_23031_20174# 0.06425f
C734 top_DAC_0/top_final_switch_0.VOUT[0] VOUT 6.7893f
C735 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 1.21986f
C736 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.0119f
C737 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 1.28355f
C738 a_19468_10031# a_20498_8950# 0.01896f
C739 a_19468_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.22126f
C740 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.21864f
C741 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 6.03974f
C742 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.06296f
C743 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.65108f
C744 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 1.49083f
C745 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_21375_20174# 0.08102f
C746 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.VS1 0.1802f
C747 a_2678_20320# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.05719f
C748 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP 0.3001f
C749 a_19552_8950# a_20076_10031# 0.04005f
C750 a_31870_7686# a_27344_6250# 0.1294f
C751 a_31318_7686# a_27896_6250# 0.02796f
C752 a_31594_7686# a_27620_6250# 0.02794f
C753 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 1.95068f
C754 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 0.01485f
C755 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_23629_18133# 0.26434f
C756 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] a_38672_20477# 0.01006f
C757 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 0.8735f
C758 VOUT a_12809_13005# 0.02119f
C759 a_18724_8950# a_19000_8950# 2.70394f
C760 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.12764f
C761 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_14615_14283# 0.02376f
C762 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.11563f
C763 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.09505f
C764 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.0288f
C765 a_17148_18696# VDDH 0.53265f
C766 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 a_20547_20174# 0.08784f
C767 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.4235f
C768 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.06152f
C769 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.09437f
C770 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_18724_8950# 0.02425f
C771 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 0.04867f
C772 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.0421f
C773 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.15407f
C774 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.02784f
C775 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.09079f
C776 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y a_44062_18449# 0.09819f
C777 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 0.14051f
C778 a_34580_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.08719f
C779 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.07852f
C780 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.03535f
C781 a_21927_20174# a_22203_20174# 1.03985f
C782 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.53884f
C783 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.14089f
C784 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.05833f
C785 a_44234_7352# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.13862f
C786 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.VH3 0.34015f
C787 a_33910_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05127f
C788 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 0.02575f
C789 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.04824f
C790 a_14607_6250# a_15041_6250# 5.50282f
C791 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_39306_20477# 0.22975f
C792 a_44234_10956# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.03152f
C793 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP a_43724_12342# 0.03147f
C794 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 1.85588f
C795 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.01121f
C796 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_6996# 0.13393f
C797 a_15618_18696# VDDH 0.25878f
C798 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A VDD 0.33616f
C799 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 0.84983f
C800 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_16891_7686# 0.06399f
C801 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB a_44234_14916# 0.08412f
C802 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 0.05743f
C803 DIN8 VDD 0.72319f
C804 DIN3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.03505f
C805 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 0.39192f
C806 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 0.05585f
C807 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] a_16596_18696# 0.03124f
C808 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.17986f
C809 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.01808f
C810 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.05995f
C811 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB a_44234_7986# 0.06683f
C812 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.05183f
C813 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44062_19161# 0.02575f
C814 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1896_12504# 0.06294f
C815 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.17402f
C816 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 a_30056_7686# 0.03929f
C817 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.01068f
C818 a_44234_12302# a_43698_11746# 0.07082f
C819 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.14301f
C820 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 17.4806f
C821 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 0.02537f
C822 a_34304_8950# a_31042_7686# 0.03954f
C823 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.08389f
C824 a_17443_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.03016f
C825 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.01646f
C826 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 1.27914f
C827 a_44234_10956# a_43698_10756# 0.0139f
C828 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.01132f
C829 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.05427f
C830 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_11629_13005# 0.0208f
C831 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 a_27620_6250# 0.02787f
C832 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.20712f
C833 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] VDD 1.04528f
C834 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04075f
C835 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.46871f
C836 a_43698_8776# a_44234_8976# 0.0139f
C837 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 a_31318_7686# 0.03989f
C838 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.16693f
C839 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 a_30608_7686# 0.08075f
C840 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.04017f
C841 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.02791f
C842 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_15629_7686# 0.1228f
C843 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_final_switch_0.VOUT[3] 0.06917f
C844 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.08478f
C845 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.08961f
C846 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.05752f
C847 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 0.01906f
C848 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.13705f
C849 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_21375_20174# 0.11545f
C850 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 a_15593_6250# 0.02794f
C851 a_16181_7686# a_17443_7686# 0.17595f
C852 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 2.17542f
C853 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 7.26391f
C854 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.01835f
C855 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.04313f
C856 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.04824f
C857 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.0239f
C858 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.25263f
C859 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.17254f
C860 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_5050_12595# 0.64856f
C861 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.1906f
C862 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 10.7528f
C863 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 12.2409f
C864 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.08701f
C865 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.11409f
C866 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.90412f
C867 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 2.89603f
C868 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.09198f
C869 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.21776f
C870 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 a_31870_7686# 0.0394f
C871 a_24209_18133# a_21927_20174# 0.06876f
C872 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.08611f
C873 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.01992f
C874 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_14331_6250# 0.16519f
C875 a_15629_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 0.07446f
C876 a_28172_6250# a_27896_6250# 8.19109f
C877 a_28882_6250# a_27344_6250# 0.18989f
C878 a_28606_6250# a_27620_6250# 0.1783f
C879 ROUT2 VDD 0.6068f
C880 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 a_16320_18696# 0.05633f
C881 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.13686f
C882 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.17799f
C883 VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.75441f
C884 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04942f
C885 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP 0.08366f
C886 a_35453_10031# a_35757_10031# 1.3412f
C887 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.15976f
C888 a_35177_10031# a_36033_10031# 0.08853f
C889 a_19946_8950# a_20498_8950# 0.10402f
C890 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C VDD 0.33516f
C891 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.05594f
C892 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.12623f
C893 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04845f
C894 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.02794f
C895 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 7.84438f
C896 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_22755_20174# 0.12485f
C897 VDDH a_43698_6796# 0.23384f
C898 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 a_14607_6250# 0.02789f
C899 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.09644f
C900 a_19276_8950# a_19000_8950# 2.74482f
C901 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.04405f
C902 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 2.23765f
C903 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.06658f
C904 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_13292# 0.14379f
C905 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.03931f
C906 a_15374_19866# VDDH 0.3323f
C907 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_16596_18696# 0.11864f
C908 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 1.25806f
C909 a_34856_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.01646f
C910 a_15317_6250# a_19946_8950# 0.03942f
C911 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.0981f
C912 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.06511f
C913 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.10418f
C914 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 0.69233f
C915 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.02784f
C916 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 a_29434_6250# 0.04772f
C917 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] DIN8 0.01582f
C918 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_19276_8950# 0.02609f
C919 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y a_44062_19161# 0.07788f
C920 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 2.15145f
C921 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 1.4939f
C922 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.04264f
C923 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.11522f
C924 a_14615_13536# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.01931f
C925 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.01675f
C926 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.98465f
C927 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.0331f
C928 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44062_20941# 0.02575f
C929 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_8173_12507# 0.02171f
C930 VDDH a_43698_15706# 0.24088f
C931 a_44062_20585# a_44062_20941# 0.12219f
C932 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 1.57718f
C933 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.23003f
C934 a_2300_15118# a_2300_14353# 0.02286f
C935 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[3] 0.59534f
C936 VDDH a_1896_21703# 0.73997f
C937 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.05677f
C938 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 1.21016f
C939 a_16181_7686# a_15041_6250# 0.03938f
C940 a_15863_13785# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.1596f
C941 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.61942f
C942 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.11733f
C943 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_final_switch_0.VOUT[2] 0.01423f
C944 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] a_18008_18696# 0.24061f
C945 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 1.58334f
C946 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.14082f
C947 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_16243# 0.07145f
C948 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.03533f
C949 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.03944f
C950 a_34186_8950# a_28172_6250# 0.0393f
C951 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.01788f
C952 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 3.33267f
C953 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.03366f
C954 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.01752f
C955 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.90443f
C956 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 a_15317_6250# 0.03792f
C957 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.041f
C958 a_33358_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.02566f
C959 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.0497f
C960 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.09244f
C961 top_DAC_0/top_final_switch_0.VOUT[2] a_9353_14150# 0.01867f
C962 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.02789f
C963 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 0.1236f
C964 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.04718f
C965 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_2678_11886# 0.04314f
C966 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.02599f
C967 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 0.01963f
C968 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 a_15041_6250# 0.03611f
C969 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 a_15041_6250# 0.02789f
C970 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 1.63811f
C971 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.05244f
C972 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 0.07667f
C973 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.18669f
C974 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_30056_7686# 0.08126f
C975 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] a_15224_18696# 0.03517f
C976 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.02122f
C977 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_final_switch_0.VOUT[3] 0.01676f
C978 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 0.02654f
C979 VDDH a_20498_8950# 0.51929f
C980 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.02784f
C981 top_DAC_0/top_final_switch_0.VOUT[2] a_9901_15057# 0.01175f
C982 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 1.23475f
C983 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_21651_20174# 0.16896f
C984 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_6445_15057# 0.04959f
C985 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 1.25889f
C986 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 1.60406f
C987 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.33598f
C988 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 3.55677f
C989 a_17443_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.21674f
C990 a_24135_20174# a_23629_18133# 0.04025f
C991 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 0.80785f
C992 a_24209_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.10167f
C993 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 a_16891_7686# 0.03929f
C994 VDDH a_15317_6250# 0.91727f
C995 VDDH a_2300_14353# 0.53441f
C996 a_19468_10031# a_20076_10031# 0.17553f
C997 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 1.63629f
C998 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_44062_20229# 0.02123f
C999 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 6.21616f
C1000 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09116f
C1001 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.13514f
C1002 a_30056_7686# a_31594_7686# 0.1611f
C1003 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.07012f
C1004 a_29780_7686# a_31870_7686# 0.38908f
C1005 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 10.1642f
C1006 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.28513f
C1007 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 a_28606_6250# 0.02787f
C1008 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 0.3156f
C1009 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.1105f
C1010 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 0.07818f
C1011 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_8976# 0.01697f
C1012 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 a_28882_6250# 0.04192f
C1013 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 a_14331_6250# 0.04485f
C1014 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 a_28606_6250# 0.11044f
C1015 a_44234_13292# a_44234_12936# 0.08026f
C1016 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 a_28172_6250# 0.02784f
C1017 DIN6 VDD 0.70858f
C1018 VOUT top_DAC_0/top_final_switch_0.VOUT[2] 6.36553f
C1019 a_30608_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.03955f
C1020 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.07772f
C1021 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_9332# 0.02028f
C1022 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_17167_7686# 0.12865f
C1023 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN a_44234_17252# 0.08412f
C1024 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.14159f
C1025 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.06101f
C1026 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 1.49134f
C1027 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_15905_7686# 0.06629f
C1028 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_23031_20174# 0.20325f
C1029 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_15353_7686# 0.0464f
C1030 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.07765f
C1031 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.06145f
C1032 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.13661f
C1033 a_31870_7686# top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.05514f
C1034 a_15374_19866# a_17148_18696# 0.09833f
C1035 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 0.01965f
C1036 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.11344f
C1037 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD 0.23151f
C1038 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_44062_18805# 0.02123f
C1039 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 a_21099_20174# 0.05514f
C1040 a_2678_10356# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.02366f
C1041 a_35757_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.34967f
C1042 a_44234_11312# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.03855f
C1043 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 0.16205f
C1044 DIN9 VDD 0.75623f
C1045 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_29434_6250# 0.29804f
C1046 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.09248f
C1047 a_15224_18696# a_14948_18696# 2.12656f
C1048 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.0151f
C1049 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_19000_8950# 0.25159f
C1050 VDDH a_43698_11746# 0.24088f
C1051 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.15447f
C1052 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_28172_6250# 0.05171f
C1053 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB a_42847_4906# 0.0113f
C1054 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.30067f
C1055 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 0.0119f
C1056 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_5642_8388# 0.10623f
C1057 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.2656f
C1058 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 0.87032f
C1059 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.10072f
C1060 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.02785f
C1061 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_21651_20174# 0.17378f
C1062 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.48284f
C1063 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04995f
C1064 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.01807f
C1065 a_15374_19866# a_15618_18696# 0.07217f
C1066 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.02793f
C1067 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.77003f
C1068 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.06435f
C1069 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 a_14331_6250# 0.02788f
C1070 a_43994_22522# VDDH 0.78839f
C1071 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.94034f
C1072 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.37332f
C1073 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_20076_10031# 0.32677f
C1074 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.03617f
C1075 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 VOUT 0.13389f
C1076 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 a_27620_6250# 0.02789f
C1077 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 8.33205f
C1078 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 0.57622f
C1079 a_2678_19053# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.01343f
C1080 a_24411_20174# a_24963_20174# 0.12523f
C1081 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 a_27896_6250# 0.02791f
C1082 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 0.02715f
C1083 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 4.14551f
C1084 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 1.2479f
C1085 a_33358_8950# a_31870_7686# 0.19113f
C1086 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 0.1146f
C1087 a_15066_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.30999f
C1088 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.2177f
C1089 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 0.57986f
C1090 a_20823_20174# a_21099_20174# 1.23587f
C1091 a_20547_20174# a_21375_20174# 0.1678f
C1092 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD 0.23023f
C1093 a_34186_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.02764f
C1094 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 0.0216f
C1095 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01428f
C1096 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 0.10409f
C1097 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.17638f
C1098 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.09063f
C1099 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 a_22479_20174# 0.08495f
C1100 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.16804f
C1101 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_14607_6250# 0.23958f
C1102 VOUT a_4717_13005# 0.0131f
C1103 a_43698_14716# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.40164f
C1104 a_16615_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.07989f
C1105 a_43698_15706# a_44234_15906# 0.0139f
C1106 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_final_switch_0.VOUT[1] 0.05518f
C1107 a_1896_22970# a_2678_22970# 0.02127f
C1108 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.01826f
C1109 top_DAC_0/top_rseg_n_dcell_0.VS4 a_19772_10031# 0.06291f
C1110 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 0.02097f
C1111 a_8473_23194# ROUT1 1.17669f
C1112 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_23031_20174# 0.19294f
C1113 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 a_13779_6250# 0.04304f
C1114 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.91327f
C1115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.42123f
C1116 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 3.59569f
C1117 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 VDDH 0.11236f
C1118 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.04843f
C1119 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_36033_10031# 0.02887f
C1120 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 0.05308f
C1121 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 a_14948_18696# 0.06345f
C1122 a_43724_16856# a_43698_16696# 0.02395f
C1123 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 a_15317_6250# 0.0856f
C1124 a_44234_16896# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.06668f
C1125 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.05423f
C1126 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 0.02734f
C1127 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.12894f
C1128 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.10061f
C1129 a_28882_6250# a_29780_7686# 0.0423f
C1130 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.12809f
C1131 a_28606_6250# a_30056_7686# 0.03909f
C1132 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.1304f
C1133 a_29158_6250# a_29434_6250# 8.10664f
C1134 top_DAC_0/top_final_switch_0.VOUT[1] a_14615_13785# 0.07338f
C1135 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 a_8051_10107# 0.03683f
C1136 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_43698_13726# 0.24498f
C1137 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.05166f
C1138 a_21375_20174# a_21927_20174# 0.15512f
C1139 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.01375f
C1140 a_20823_20174# a_22479_20174# 0.13852f
C1141 a_21099_20174# a_22203_20174# 0.14267f
C1142 a_20547_20174# a_22755_20174# 0.17927f
C1143 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 a_37022_20713# 0.04385f
C1144 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.01142f
C1145 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.1019f
C1146 a_6923_9707# top_DAC_0/top_final_switch_0.VOUT[4] 0.43838f
C1147 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_final_switch_0.VOUT[1] 5.80043f
C1148 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.20436f
C1149 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 1.24994f
C1150 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 0.02015f
C1151 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.21475f
C1152 a_44234_8976# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.06335f
C1153 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.05032f
C1154 a_2678_19053# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.0593f
C1155 a_31870_7686# a_27896_6250# 0.06285f
C1156 a_20222_8950# a_19772_10031# 0.0125f
C1157 a_7625_12507# a_8173_12507# 0.0103f
C1158 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.07143f
C1159 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 a_22479_20174# 0.04149f
C1160 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 0.08515f
C1161 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_final_switch_0.VOUT[2] 0.01655f
C1162 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.09106f
C1163 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.09702f
C1164 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.15627f
C1165 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04935f
C1166 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05891f
C1167 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.01642f
C1168 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.08561f
C1169 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 a_27344_6250# 0.04335f
C1170 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09062f
C1171 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.04304f
C1172 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] DIN9 0.17935f
C1173 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.0203f
C1174 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.11246f
C1175 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.06886f
C1176 a_17732_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.1136f
C1177 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.11034f
C1178 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.09869f
C1179 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 a_27896_6250# 0.03927f
C1180 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.0864f
C1181 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.41311f
C1182 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 0.16157f
C1183 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.02784f
C1184 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.08546f
C1185 DIN6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.03492f
C1186 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.02791f
C1187 a_44234_12302# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.02704f
C1188 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.15569f
C1189 a_35132_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.0684f
C1190 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 0.11409f
C1191 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.VL3 0.0398f
C1192 a_19276_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.01953f
C1193 a_21927_20174# a_22755_20174# 0.17759f
C1194 a_22203_20174# a_22479_20174# 1.1942f
C1195 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.04039f
C1196 a_34304_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.04818f
C1197 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15066_18696# 0.12138f
C1198 a_15863_13785# top_DAC_0/top_final_switch_0.VOUT[2] 0.0759f
C1199 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.0249f
C1200 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.03419f
C1201 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 1.789f
C1202 a_43698_9766# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.01234f
C1203 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.16951f
C1204 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.04329f
C1205 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_27620_6250# 0.12436f
C1206 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.10472f
C1207 a_1896_17510# a_2678_17510# 0.02127f
C1208 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_17443_7686# 0.28489f
C1209 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.06038f
C1210 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 0.05551f
C1211 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_16891_7686# 0.05967f
C1212 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.14262f
C1213 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.04843f
C1214 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 1.19056f
C1215 a_23049_18133# a_20547_20174# 0.04087f
C1216 a_22469_18133# a_20823_20174# 0.06841f
C1217 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 1.2419f
C1218 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 0.0944f
C1219 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 15.7968f
C1220 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.05594f
C1221 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.VL3 0.03007f
C1222 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 0.0847f
C1223 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.04651f
C1224 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 1.33973f
C1225 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.40016f
C1226 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.04219f
C1227 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.31321f
C1228 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 1.48649f
C1229 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A VDDH 0.90804f
C1230 VDDH top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 4.75556f
C1231 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.82681f
C1232 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_7625_15057# 0.04959f
C1233 a_44234_11312# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.14379f
C1234 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] VDD 1.73139f
C1235 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.15349f
C1236 a_34580_8950# a_31318_7686# 0.03944f
C1237 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.16534f
C1238 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.11848f
C1239 a_43698_9766# a_43698_10756# 0.01563f
C1240 a_43724_10916# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP 0.08245f
C1241 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.17853f
C1242 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_2678_12504# 0.04249f
C1243 VDDH a_20076_10031# 0.2709f
C1244 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_12809_13005# 0.01625f
C1245 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.02948f
C1246 VDDH a_43724_9926# 0.09227f
C1247 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.47771f
C1248 a_43698_9766# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.06167f
C1249 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 0.22168f
C1250 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.88317f
C1251 VDDH a_43698_8776# 0.23565f
C1252 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.05823f
C1253 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_16181_7686# 0.11336f
C1254 a_21375_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.08147f
C1255 DIN7 VDD 0.71581f
C1256 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.02121f
C1257 VOUT a_8173_14150# 0.0409f
C1258 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.13217f
C1259 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.02615f
C1260 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 1.47977f
C1261 a_7625_15057# a_8173_15057# 0.0237f
C1262 a_22469_18133# a_22203_20174# 0.04096f
C1263 DIN3 DIN2 0.33146f
C1264 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.04651f
C1265 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.02147f
C1266 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_33910_8950# 0.11409f
C1267 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 0.58367f
C1268 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.03532f
C1269 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 0.05687f
C1270 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.8597f
C1271 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.85676f
C1272 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 0.13531f
C1273 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.06701f
C1274 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.13022f
C1275 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.10358f
C1276 a_43698_7786# a_43724_8382# 0.06762f
C1277 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.09591f
C1278 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.04804f
C1279 a_24209_18133# a_22479_20174# 0.06806f
C1280 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A a_43724_9372# 0.03253f
C1281 a_4978_8388# a_5642_8388# 0.02543f
C1282 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.98177f
C1283 a_44062_19517# a_44062_19161# 0.12219f
C1284 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_15041_6250# 0.24058f
C1285 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 10.5451f
C1286 a_29434_6250# a_27344_6250# 0.21524f
C1287 a_28882_6250# a_27896_6250# 0.15498f
C1288 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 0.0245f
C1289 a_29158_6250# a_27620_6250# 0.15325f
C1290 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.12365f
C1291 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 a_29158_6250# 0.03953f
C1292 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.26862f
C1293 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 1.16389f
C1294 a_8051_10107# top_DAC_0/top_final_switch_0.VOUT[3] 0.43675f
C1295 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.30956f
C1296 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y a_44062_18093# 0.07788f
C1297 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 a_29158_6250# 0.01211f
C1298 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 0.03198f
C1299 a_35757_10031# a_36033_10031# 0.93291f
C1300 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.01283f
C1301 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 1.73225f
C1302 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_16896# 0.02704f
C1303 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_20498_8950# 0.10233f
C1304 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 1.13576f
C1305 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 0.7035f
C1306 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 a_5050_12595# 0.17196f
C1307 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_23307_20174# 0.13941f
C1308 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.01611f
C1309 a_15593_6250# a_20222_8950# 0.0394f
C1310 a_15863_13287# top_DAC_0/top_final_switch_0.VOUT[0] 0.07961f
C1311 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.09354f
C1312 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_17252# 0.03345f
C1313 a_8051_10107# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.2514f
C1314 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 1.3506f
C1315 a_5897_14150# a_6445_14150# 0.0237f
C1316 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.10472f
C1317 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP 0.01045f
C1318 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_31870_7686# 0.21933f
C1319 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.19135f
C1320 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.21387f
C1321 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 a_30056_7686# 0.04025f
C1322 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 0.16861f
C1323 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.04086f
C1324 a_6445_13005# a_5897_13005# 0.0103f
C1325 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 0.12736f
C1326 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.84452f
C1327 a_6778_12595# a_5050_12595# 2.85565f
C1328 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 0.16476f
C1329 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.05164f
C1330 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.20364f
C1331 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 a_17443_7686# 0.03929f
C1332 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 1.54852f
C1333 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.01649f
C1334 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.05322f
C1335 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.10646f
C1336 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD 0.21864f
C1337 VDDH a_8473_23194# 0.06477f
C1338 a_44062_22009# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.06327f
C1339 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 a_14055_6250# 0.03971f
C1340 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.09372f
C1341 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.01088f
C1342 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.08827f
C1343 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 a_28882_6250# 0.08556f
C1344 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44737_4828# 0.04364f
C1345 VDDH a_41907_22057# 0.31401f
C1346 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.VL3 0.05812f
C1347 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.06052f
C1348 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.09474f
C1349 a_22469_18133# a_24209_18133# 0.22368f
C1350 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.03879f
C1351 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 a_28172_6250# 0.03927f
C1352 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.56233f
C1353 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 1.81035f
C1354 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.05253f
C1355 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.10242f
C1356 a_34304_8950# a_28606_6250# 0.03945f
C1357 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.09577f
C1358 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 a_30608_7686# 0.07998f
C1359 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 a_15869_6250# 0.29269f
C1360 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[4] 0.47259f
C1361 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.10422f
C1362 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] VDD 1.60464f
C1363 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 0.06597f
C1364 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.05607f
C1365 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 0.01023f
C1366 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 0.60342f
C1367 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.VH3 0.01446f
C1368 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.21911f
C1369 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] a_14672_18696# 0.0525f
C1370 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 0.13233f
C1371 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.06718f
C1372 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.6218f
C1373 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.09992f
C1374 DIN8 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.17935f
C1375 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.02785f
C1376 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 0.01927f
C1377 a_23859_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.88724f
C1378 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.17921f
C1379 top_DAC_0/top_final_switch_0.VOUT[0] a_6445_14150# 0.01199f
C1380 VDDH DIN8 0.4277f
C1381 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.04138f
C1382 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 2.97868f
C1383 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.12599f
C1384 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04845f
C1385 a_24687_20174# a_23629_18133# 0.04272f
C1386 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_final_switch_0.VOUT[3] 0.01093f
C1387 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_30608_7686# 0.08023f
C1388 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.05622f
C1389 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05297f
C1390 VDDH a_15869_6250# 1.05868f
C1391 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 1.92248f
C1392 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.70128f
C1393 a_22755_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 0.11072f
C1394 a_19468_10031# a_20656_10031# 0.06376f
C1395 a_4415_23194# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.01802f
C1396 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.60156f
C1397 a_43391_3326# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.01036f
C1398 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.VH3 0.09189f
C1399 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_final_switch_0.VOUT[4] 0.5995f
C1400 a_22755_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 0.08577f
C1401 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] a_45343_3978# 0.01187f
C1402 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.16773f
C1403 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.05244f
C1404 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 a_29158_6250# 0.02787f
C1405 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.15598f
C1406 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.11989f
C1407 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 0.07638f
C1408 VDDH a_43724_13886# 0.09227f
C1409 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 a_28606_6250# 0.039f
C1410 a_17732_18696# a_18008_18696# 0.85268f
C1411 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 2.1111f
C1412 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_9901_13005# 0.0208f
C1413 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 a_29434_6250# 0.08622f
C1414 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 a_15041_6250# 0.04056f
C1415 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 0.24855f
C1416 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 a_28882_6250# 0.02784f
C1417 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.01273f
C1418 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN a_44234_8342# 0.06685f
C1419 a_37022_20295# a_36888_19550# 0.01701f
C1420 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_final_switch_0.VOUT[2] 5.5062f
C1421 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.35945f
C1422 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_final_switch_0.VOUT[2] 0.20339f
C1423 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.39803f
C1424 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 a_27896_6250# 0.08519f
C1425 a_15863_13785# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.03829f
C1426 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.63397f
C1427 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.09111f
C1428 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.57187f
C1429 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_15905_7686# 0.05946f
C1430 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 9.82456f
C1431 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.13355f
C1432 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 a_16615_7686# 0.03998f
C1433 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.02029f
C1434 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 18.2729f
C1435 a_35757_10031# a_33910_8950# 0.0648f
C1436 a_35453_10031# a_34186_8950# 0.06482f
C1437 a_35177_10031# a_34304_8950# 0.05067f
C1438 a_27344_6250# a_27620_6250# 8.06436f
C1439 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.04736f
C1440 a_36033_10031# a_33634_8950# 0.06493f
C1441 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 1.18085f
C1442 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 VDDH 1.27454f
C1443 a_14790_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.25324f
C1444 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_30056_7686# 0.11409f
C1445 a_15224_18696# a_16320_18696# 0.08897f
C1446 a_14948_18696# a_14672_18696# 2.57618f
C1447 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 a_37804_20295# 0.0477f
C1448 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 ROUT2 0.01358f
C1449 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.1547f
C1450 a_17148_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.0309f
C1451 VOUT a_12809_12507# 0.04641f
C1452 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 0.69152f
C1453 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_28882_6250# 0.05568f
C1454 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.0582f
C1455 a_33910_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.36318f
C1456 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.12688f
C1457 a_17167_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.07166f
C1458 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 a_15317_6250# 0.02785f
C1459 a_43698_13726# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP 0.7858f
C1460 a_44062_20229# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.1286f
C1461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 0.48023f
C1462 a_43724_11906# VDDH 0.09227f
C1463 VDDH ROUT2 9.92565f
C1464 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.SH[2] 16.9983f
C1465 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_final_switch_0.VOUT[2] 0.01082f
C1466 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.07771f
C1467 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 0.10826f
C1468 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_8936# 0.03597f
C1469 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.02803f
C1470 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.02015f
C1471 VDDH a_4717_14150# 0.48125f
C1472 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 a_15041_6250# 0.0279f
C1473 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.06058f
C1474 VDDH a_1896_19053# 0.722f
C1475 a_39861_22057# VDDH 0.2924f
C1476 a_30056_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.03087f
C1477 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 0.01326f
C1478 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A a_43698_6796# 0.40011f
C1479 a_23629_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.08418f
C1480 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.0433f
C1481 a_43698_7786# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.02387f
C1482 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 11.5953f
C1483 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_30608_7686# 0.11721f
C1484 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 1.39454f
C1485 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 1.68068f
C1486 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.57553f
C1487 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_19670_8950# 0.02521f
C1488 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VDDH 3.43289f
C1489 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_final_switch_0.VOUT[3] 0.05206f
C1490 a_15618_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.51672f
C1491 a_5050_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.19638f
C1492 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.06721f
C1493 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.05182f
C1494 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 a_23307_20174# 0.06406f
C1495 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 0.06117f
C1496 a_21099_20174# a_21375_20174# 0.95595f
C1497 a_20823_20174# a_21651_20174# 0.18401f
C1498 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 a_28606_6250# 0.02791f
C1499 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.91043f
C1500 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 0.01784f
C1501 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 0.04147f
C1502 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.0888f
C1503 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[2] 0.39626f
C1504 a_16891_7686# a_19670_8950# 0.1105f
C1505 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05983f
C1506 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.15602f
C1507 a_24135_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.17801f
C1508 a_16615_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.03947f
C1509 VOUT a_5897_13005# 0.02204f
C1510 a_6778_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 0.10076f
C1511 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_1896_21703# 0.0991f
C1512 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] VDD 1.57937f
C1513 a_36888_19786# a_36888_19550# 2.53242f
C1514 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.02784f
C1515 a_33634_8950# a_27620_6250# 0.03929f
C1516 VDDH a_43724_7946# 0.09227f
C1517 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 a_14331_6250# 0.02786f
C1518 a_44234_11946# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP 0.06668f
C1519 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.3935f
C1520 a_30332_7686# a_31042_7686# 0.17054f
C1521 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB VDD 0.67205f
C1522 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 0.06133f
C1523 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.09502f
C1524 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 1.04282f
C1525 a_44234_15272# a_44234_15906# 0.02262f
C1526 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 0.01392f
C1527 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.31886f
C1528 a_31594_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.03944f
C1529 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02801f
C1530 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.19767f
C1531 a_43698_15706# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.40164f
C1532 VDDH a_4717_15057# 0.49013f
C1533 top_DAC_0/top_rseg_n_dcell_0.VH2 a_21375_20174# 0.01296f
C1534 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.VH3 0.05427f
C1535 a_29158_6250# a_30056_7686# 0.02791f
C1536 a_29434_6250# a_29780_7686# 0.28232f
C1537 VOUT a_6778_12595# 0.46013f
C1538 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 0.05163f
C1539 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 1.73155f
C1540 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.04379f
C1541 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.1193f
C1542 a_21651_20174# a_22203_20174# 0.26801f
C1543 a_21375_20174# a_22479_20174# 0.15298f
C1544 a_20547_20174# a_23307_20174# 0.17801f
C1545 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 a_36888_19550# 0.58096f
C1546 a_21099_20174# a_22755_20174# 0.17726f
C1547 a_20823_20174# a_23031_20174# 0.13276f
C1548 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.12539f
C1549 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.0478f
C1550 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.02789f
C1551 a_8051_10107# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.03682f
C1552 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.09312f
C1553 DIN3 VDD 0.67007f
C1554 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB a_44234_6996# 0.07436f
C1555 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.56064f
C1556 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_21927_20174# 0.0314f
C1557 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.02787f
C1558 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01425f
C1559 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 1.40144f
C1560 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.69015f
C1561 a_20498_8950# a_20076_10031# 0.05271f
C1562 a_20222_8950# a_20352_10031# 0.04441f
C1563 a_19552_8950# a_18724_8950# 0.09125f
C1564 a_19946_8950# a_20656_10031# 0.04106f
C1565 a_19670_8950# a_20932_10031# 0.04084f
C1566 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_20076_10031# 0.07139f
C1567 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.06276f
C1568 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 a_27344_6250# 0.04702f
C1569 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_17148_18696# 0.15001f
C1570 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.02786f
C1571 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 a_27620_6250# 0.05097f
C1572 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_12342# 0.03597f
C1573 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 0.5522f
C1574 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB DIN1 0.01607f
C1575 VDDH a_16615_7686# 0.46016f
C1576 a_14607_6250# a_19552_8950# 0.0393f
C1577 a_18284_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.07188f
C1578 a_43698_16696# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.01799f
C1579 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y VDD 0.33964f
C1580 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 VOUT 0.17766f
C1581 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.12411f
C1582 a_33634_8950# a_33910_8950# 2.89482f
C1583 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_4717_13005# 0.02092f
C1584 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.04091f
C1585 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.61305f
C1586 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.02784f
C1587 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.31049f
C1588 a_44234_16896# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.08412f
C1589 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.02791f
C1590 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.19658f
C1591 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_15906# 0.02704f
C1592 a_24135_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.11869f
C1593 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 a_15041_6250# 0.11045f
C1594 a_22203_20174# a_23031_20174# 0.13292f
C1595 a_22479_20174# a_22755_20174# 6.25438f
C1596 a_21927_20174# a_23307_20174# 0.17704f
C1597 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 2.07729f
C1598 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 0.08427f
C1599 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.96636f
C1600 VDDH DIN6 0.42765f
C1601 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.02032f
C1602 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.05716f
C1603 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.01028f
C1604 a_34856_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.04765f
C1605 a_15863_13287# top_DAC_0/top_final_switch_0.VOUT[2] 0.02598f
C1606 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15618_18696# 0.19271f
C1607 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.18751f
C1608 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 3.7974f
C1609 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_10322# 0.01697f
C1610 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 1.39623f
C1611 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.05213f
C1612 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_16262# 0.03152f
C1613 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.02116f
C1614 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_1896_16243# 0.0335f
C1615 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 0.05125f
C1616 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_final_switch_0.VOUT[3] 0.01337f
C1617 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_19670_8950# 0.05389f
C1618 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_38672_20477# 0.12954f
C1619 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_17443_7686# 0.26279f
C1620 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 0.0658f
C1621 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.04022f
C1622 a_23859_20174# a_20547_20174# 0.33451f
C1623 a_22469_18133# a_21375_20174# 0.08772f
C1624 a_23049_18133# a_21099_20174# 0.04207f
C1625 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.08366f
C1626 a_23583_20174# a_20823_20174# 0.13239f
C1627 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.17262f
C1628 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 8.31336f
C1629 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.33162f
C1630 a_1636_13708# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.02725f
C1631 a_42847_3710# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.01316f
C1632 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 a_14055_6250# 0.0358f
C1633 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.11045f
C1634 VDDH a_43698_14716# 0.24088f
C1635 a_45015_4828# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.01008f
C1636 a_33358_8950# a_29434_6250# 0.02007f
C1637 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.02784f
C1638 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.04526f
C1639 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_4717_14150# 0.05017f
C1640 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.04623f
C1641 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 0.09468f
C1642 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.01904f
C1643 VDDH DIN9 0.40422f
C1644 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.17257f
C1645 a_34856_8950# a_31594_7686# 0.03939f
C1646 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.02523f
C1647 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.10475f
C1648 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.06092f
C1649 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] VDD 2.59466f
C1650 a_44234_11312# a_44234_10956# 0.08026f
C1651 VDDH a_20656_10031# 0.2252f
C1652 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.08257f
C1653 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 0.11409f
C1654 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.11848f
C1655 a_9901_15057# top_DAC_0/top_final_switch_0.VOUT[3] 0.03029f
C1656 a_30056_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.05396f
C1657 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.11469f
C1658 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 0.20097f
C1659 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_24209_18133# 0.42807f
C1660 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.05244f
C1661 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 1.64648f
C1662 VDDH a_14055_6250# 0.64476f
C1663 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 2.84584f
C1664 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.18515f
C1665 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.62163f
C1666 a_14514_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.53315f
C1667 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.12088f
C1668 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_44062_18449# 0.02123f
C1669 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_final_switch_0.VOUT[2] 0.01823f
C1670 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.04326f
C1671 DIN5 DIN6 0.36448f
C1672 top_DAC_0/top_rseg_n_dcell_0.VH2 a_23049_18133# 0.4769f
C1673 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 1.30585f
C1674 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 1.26639f
C1675 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.03957f
C1676 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_10362# 0.03597f
C1677 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 0.10213f
C1678 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 0.71512f
C1679 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 a_15905_7686# 0.03985f
C1680 a_23583_20174# a_22203_20174# 0.13241f
C1681 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 0.12957f
C1682 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09013f
C1683 a_23859_20174# a_21927_20174# 0.15658f
C1684 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.03606f
C1685 a_22469_18133# a_22755_20174# 0.07062f
C1686 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.02791f
C1687 top_DAC_0/top_final_switch_0.VOUT[1] a_8173_14150# 0.01201f
C1688 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.15968f
C1689 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 0.2711f
C1690 a_1896_10974# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.03761f
C1691 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 8.23983f
C1692 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.61039f
C1693 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_34304_8950# 0.11454f
C1694 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_19000_8950# 0.1703f
C1695 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.02113f
C1696 a_43698_12736# VDDH 0.24088f
C1697 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_37410_19098# 0.37572f
C1698 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.18941f
C1699 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 3.26761f
C1700 VOUT top_DAC_0/top_final_switch_0.VOUT[3] 6.36704f
C1701 top_DAC_0/top_rseg_n_dcell_0.VL2 a_23629_18133# 0.72984f
C1702 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_8976# 0.01693f
C1703 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 1.45438f
C1704 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC a_38584_20665# 0.02697f
C1705 a_43698_7786# a_44234_7986# 0.0139f
C1706 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 14.96f
C1707 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04863f
C1708 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.98976f
C1709 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A a_44234_8976# 0.05897f
C1710 VDDH top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.63542f
C1711 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 2.14311f
C1712 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.0852f
C1713 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.03375f
C1714 a_29780_7686# a_27620_6250# 0.04204f
C1715 a_30056_7686# a_27344_6250# 0.03758f
C1716 a_29434_6250# a_27896_6250# 0.17891f
C1717 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 a_14055_6250# 0.03971f
C1718 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.6099f
C1719 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.05843f
C1720 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 0.05254f
C1721 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.29277f
C1722 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.04293f
C1723 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.05844f
C1724 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.0166f
C1725 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.17721f
C1726 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.VL3 0.11021f
C1727 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 a_29780_7686# 0.03929f
C1728 VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.02946f
C1729 a_36033_10031# a_33358_8950# 0.0898f
C1730 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 1.87285f
C1731 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.06101f
C1732 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.02567f
C1733 a_19276_8950# a_19552_8950# 2.75909f
C1734 a_15905_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.03985f
C1735 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.06171f
C1736 a_5050_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.0665f
C1737 a_4415_23194# ROUT1 6.87753f
C1738 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 4.1684f
C1739 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.22509f
C1740 a_6445_15057# VOUT 0.01454f
C1741 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.09125f
C1742 a_16181_7686# a_19552_8950# 0.03938f
C1743 a_15869_6250# a_20498_8950# 0.03965f
C1744 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.05327f
C1745 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD a_8173_15057# 0.01033f
C1746 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 0.14136f
C1747 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 0.9064f
C1748 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 a_31042_7686# 0.03996f
C1749 a_22469_18133# a_23049_18133# 3.93715f
C1750 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 0.06364f
C1751 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 a_30332_7686# 0.0757f
C1752 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.02784f
C1753 a_15317_6250# a_15869_6250# 0.17854f
C1754 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 0.02106f
C1755 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.07378f
C1756 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 2.81584f
C1757 a_35177_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.07138f
C1758 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.02308f
C1759 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.VS1 1.245f
C1760 a_44062_21297# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.06327f
C1761 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_23859_20174# 0.04967f
C1762 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.22976f
C1763 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.10924f
C1764 a_2300_13352# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.03772f
C1765 VDDH a_40525_21457# 0.35437f
C1766 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.11409f
C1767 a_44234_9332# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.06554f
C1768 a_33634_8950# a_30056_7686# 0.03932f
C1769 a_34580_8950# a_28882_6250# 0.03942f
C1770 DIN5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.01586f
C1771 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_16856# 0.03597f
C1772 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 a_15629_7686# 0.07245f
C1773 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.14577f
C1774 VDDH a_43724_14876# 0.09227f
C1775 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.01642f
C1776 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 0.01397f
C1777 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.01617f
C1778 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 a_31594_7686# 0.03944f
C1779 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] VDDH 1.07221f
C1780 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.30111f
C1781 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.11842f
C1782 a_33358_8950# a_27620_6250# 0.11111f
C1783 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.08498f
C1784 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 ROUT2 0.23312f
C1785 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_14282# 0.02704f
C1786 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 1.86798f
C1787 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 a_14672_18696# 0.07029f
C1788 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 0.18787f
C1789 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 1.94253f
C1790 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09789f
C1791 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.VS4 0.74491f
C1792 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.22275f
C1793 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.58792f
C1794 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.13753f
C1795 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15317_6250# 0.17027f
C1796 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.06117f
C1797 a_24963_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 0.04148f
C1798 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.17276f
C1799 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.25749f
C1800 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.10201f
C1801 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 11.8244f
C1802 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_31318_7686# 0.07527f
C1803 VDDH a_15629_7686# 0.60256f
C1804 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 11.41f
C1805 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_16596_18696# 0.01716f
C1806 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 1.25122f
C1807 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.25693f
C1808 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.04843f
C1809 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.08451f
C1810 a_5111_10963# a_4978_10963# 0.02841f
C1811 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 a_16596_18696# 0.06355f
C1812 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB DIN2 0.17961f
C1813 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 0.06043f
C1814 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.19835f
C1815 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.01056f
C1816 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04368f
C1817 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.14077f
C1818 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.22837f
C1819 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 a_29158_6250# 0.04275f
C1820 a_39883_19479# a_38672_20477# 0.01392f
C1821 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 2.43082f
C1822 a_19772_10031# a_20352_10031# 0.17109f
C1823 a_18008_18696# a_18284_18696# 0.53191f
C1824 a_17732_18696# top_DAC_0/top_rseg_n_dcell_0.VL3 0.07318f
C1825 VDDH a_8173_15057# 0.49886f
C1826 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.VS4 0.01859f
C1827 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 a_29434_6250# 0.04091f
C1828 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_final_switch_0.VOUT[3] 0.07232f
C1829 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A a_43698_8776# 0.02387f
C1830 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_final_switch_0.VOUT[3] 0.5979f
C1831 a_15863_13536# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.1455f
C1832 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 0.09855f
C1833 a_37410_19098# a_36888_19786# 0.01634f
C1834 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.05244f
C1835 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.09083f
C1836 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 a_20547_20174# 0.01747f
C1837 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 a_27896_6250# 0.08519f
C1838 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.05769f
C1839 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04809f
C1840 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 a_16596_18696# 0.06085f
C1841 DIN7 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.01582f
C1842 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 0.01634f
C1843 top_DAC_0/top_rseg_n_dcell_0.VL2 a_14615_14283# 0.04364f
C1844 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_14322# 0.03597f
C1845 VDDH DIN7 0.42767f
C1846 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 0.0562f
C1847 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.03132f
C1848 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.05001f
C1849 a_33358_8950# a_33910_8950# 0.10275f
C1850 a_34873_10031# a_35132_8950# 0.01422f
C1851 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 2.28703f
C1852 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 0.04143f
C1853 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.VS4 0.03139f
C1854 a_27620_6250# a_27896_6250# 8.11706f
C1855 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.2455f
C1856 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_19552_8950# 0.09559f
C1857 a_15342_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.05485f
C1858 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.5508f
C1859 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.26321f
C1860 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.VS1 0.06165f
C1861 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.04809f
C1862 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 2.91357f
C1863 a_15224_18696# a_16872_18696# 0.08844f
C1864 a_14672_18696# a_16320_18696# 1.87591f
C1865 a_14948_18696# a_16596_18696# 0.089f
C1866 a_44234_12302# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.03855f
C1867 a_15863_13785# top_DAC_0/top_final_switch_0.VOUT[3] 0.01312f
C1868 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_8976# 0.1344f
C1869 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_14615_14034# 0.07377f
C1870 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 0.06039f
C1871 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 0.66055f
C1872 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_29434_6250# 0.02393f
C1873 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.04946f
C1874 a_9353_14150# a_9901_14150# 0.0237f
C1875 a_34304_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.22273f
C1876 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_12809_12507# 0.01625f
C1877 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 a_23307_20174# 0.05516f
C1878 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 a_15869_6250# 0.04181f
C1879 a_43724_11906# a_43698_11746# 0.02395f
C1880 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 2.40873f
C1881 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP VDDH 0.92594f
C1882 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 0.04159f
C1883 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 0.05286f
C1884 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.05329f
C1885 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.1675f
C1886 VDDH a_1896_17510# 0.722f
C1887 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_8342# 0.01727f
C1888 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.08344f
C1889 top_DAC_0/top_final_switch_0.VOUT[3] a_11081_15057# 0.03805f
C1890 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 1.3376f
C1891 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_44062_18449# 0.06327f
C1892 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_14948_18696# 0.17366f
C1893 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.04593f
C1894 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_31318_7686# 0.12561f
C1895 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.VH3 0.0514f
C1896 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.27327f
C1897 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.02537f
C1898 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP 0.01782f
C1899 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx a_2678_16243# 0.08404f
C1900 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_20222_8950# 0.02761f
C1901 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 0.54711f
C1902 a_43994_22522# ROUT2 0.41323f
C1903 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 0.04809f
C1904 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 0.0191f
C1905 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.04282f
C1906 a_15905_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 0.07575f
C1907 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 a_28172_6250# 0.03205f
C1908 a_21375_20174# a_21651_20174# 6.3301f
C1909 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 1.97444f
C1910 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_30332_7686# 0.07894f
C1911 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 a_29158_6250# 0.02801f
C1912 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 7.06738f
C1913 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.07698f
C1914 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 1.08835f
C1915 a_17167_7686# a_19946_8950# 0.08495f
C1916 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 a_28606_6250# 0.0331f
C1917 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 1.36225f
C1918 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 a_20823_20174# 0.06241f
C1919 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_21375_20174# 0.20237f
C1920 a_31042_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.07987f
C1921 a_35132_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.20946f
C1922 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_21099_20174# 0.03179f
C1923 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 a_21099_20174# 0.05513f
C1924 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.17762f
C1925 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.09478f
C1926 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.0232f
C1927 a_30332_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.03985f
C1928 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.06435f
C1929 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02537f
C1930 a_43698_15706# a_43698_14716# 0.01563f
C1931 VOUT a_5897_12507# 0.04473f
C1932 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.09057f
C1933 a_14790_18696# a_17732_18696# 0.35769f
C1934 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.04531f
C1935 a_33910_8950# a_27896_6250# 0.03929f
C1936 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.19335f
C1937 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.08559f
C1938 a_15317_6250# a_16615_7686# 0.028f
C1939 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.05786f
C1940 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.4978f
C1941 VOUT a_9901_14150# 0.0409f
C1942 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.11409f
C1943 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.26099f
C1944 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 a_15041_6250# 0.02789f
C1945 a_43698_10756# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP 0.40164f
C1946 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.03927f
C1947 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.04984f
C1948 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.09259f
C1949 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09485f
C1950 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 0.06393f
C1951 a_30608_7686# a_31318_7686# 0.16678f
C1952 a_30332_7686# a_31594_7686# 0.16165f
C1953 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 11.1111f
C1954 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.05167f
C1955 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_24209_18133# 0.38802f
C1956 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_28172_6250# 0.52753f
C1957 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP 0.3001f
C1958 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.02796f
C1959 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.01045f
C1960 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_8382# 0.03597f
C1961 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.01392f
C1962 a_29780_7686# a_30056_7686# 6.53418f
C1963 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 10.4407f
C1964 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.02015f
C1965 VOUT a_6445_12507# 0.03463f
C1966 a_21099_20174# a_23307_20174# 0.17696f
C1967 a_21375_20174# a_23031_20174# 0.14456f
C1968 a_21651_20174# a_22755_20174# 0.17716f
C1969 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 0.02715f
C1970 top_DAC_0/top_final_switch_0.VOUT[1] a_6778_12595# 0.43692f
C1971 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] VDDH 0.01064f
C1972 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.21492f
C1973 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 1.36638f
C1974 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04929f
C1975 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.02794f
C1976 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 14.4869f
C1977 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_6778_12595# 0.51626f
C1978 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 0.05786f
C1979 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.1264f
C1980 VDDH a_4415_23194# 31.1956f
C1981 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.09823f
C1982 DIN3 DIN4 0.3362f
C1983 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 a_22203_20174# 0.07766f
C1984 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_22755_20174# 0.03178f
C1985 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.02115f
C1986 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.02787f
C1987 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.6219f
C1988 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.03934f
C1989 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.03985f
C1990 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.03852f
C1991 a_19670_8950# a_19000_8950# 0.0814f
C1992 a_19946_8950# a_18724_8950# 0.09865f
C1993 a_20498_8950# a_20656_10031# 0.01885f
C1994 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 0.01524f
C1995 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.06214f
C1996 a_7625_15057# VOUT 0.04641f
C1997 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.SH[1] 2.74289f
C1998 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_20656_10031# 0.25734f
C1999 VDDH a_43724_13332# 0.09227f
C2000 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.96629f
C2001 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 a_27896_6250# 0.02788f
C2002 VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.21011f
C2003 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.05138f
C2004 DIN0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.01622f
C2005 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD a_9353_15057# 0.01034f
C2006 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.05384f
C2007 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 a_15593_6250# 0.02801f
C2008 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 a_27344_6250# 0.05187f
C2009 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.09202f
C2010 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.02789f
C2011 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.04066f
C2012 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 0.02715f
C2013 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 0.51123f
C2014 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.29337f
C2015 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 a_27620_6250# 0.02784f
C2016 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_16896# 0.03855f
C2017 a_34304_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.01715f
C2018 VDDH a_17167_7686# 0.58575f
C2019 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.61294f
C2020 a_15041_6250# a_19670_8950# 0.03945f
C2021 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.10302f
C2022 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.08269f
C2023 a_33910_8950# a_34186_8950# 2.84824f
C2024 a_33634_8950# a_34304_8950# 0.0814f
C2025 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.02207f
C2026 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.02784f
C2027 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.0386f
C2028 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.15473f
C2029 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_5897_13005# 0.0208f
C2030 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 0.02501f
C2031 a_34580_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.02838f
C2032 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.04747f
C2033 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 1.81252f
C2034 a_24135_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 0.04172f
C2035 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.06161f
C2036 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.11586f
C2037 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 1.25389f
C2038 a_15593_6250# a_13779_6250# 0.18773f
C2039 a_22479_20174# a_23307_20174# 0.17763f
C2040 a_15317_6250# a_14055_6250# 0.15453f
C2041 a_22755_20174# a_23031_20174# 1.10111f
C2042 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.1506f
C2043 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 2.63875f
C2044 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.07088f
C2045 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.0483f
C2046 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 0.05349f
C2047 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 ROUT1 0.01978f
C2048 VDDH a_20547_20174# 0.04145f
C2049 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.08468f
C2050 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.24317f
C2051 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 0.01966f
C2052 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 a_23307_20174# 0.05525f
C2053 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.09845f
C2054 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] a_14948_18696# 0.02569f
C2055 a_43698_7786# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.01234f
C2056 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04937f
C2057 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.07928f
C2058 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.05179f
C2059 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.04851f
C2060 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_20222_8950# 0.05287f
C2061 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.24087f
C2062 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.10002f
C2063 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_27620_6250# 0.06546f
C2064 a_24135_20174# a_20823_20174# 0.1324f
C2065 a_23583_20174# a_21375_20174# 0.14452f
C2066 a_24411_20174# a_20547_20174# 0.13321f
C2067 a_23859_20174# a_21099_20174# 0.16643f
C2068 a_23049_18133# a_21651_20174# 0.0732f
C2069 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.15073f
C2070 a_39768_20665# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.01079f
C2071 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 a_14607_6250# 0.04142f
C2072 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 a_14948_18696# 0.06348f
C2073 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 0.80029f
C2074 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_6778_12595# 0.55664f
C2075 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_9966# 0.01931f
C2076 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.40324f
C2077 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.10246f
C2078 a_44234_8342# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.06328f
C2079 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 0.01929f
C2080 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.36573f
C2081 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 0.05302f
C2082 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.0279f
C2083 VDDH a_1896_20320# 0.72706f
C2084 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.17474f
C2085 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.10771f
C2086 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.03876f
C2087 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_43698_16696# 0.01234f
C2088 a_44234_12302# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.14379f
C2089 a_35132_8950# a_31870_7686# 0.04133f
C2090 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 0.3226f
C2091 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_final_switch_0.VOUT[4] 0.02498f
C2092 VDDH a_18724_8950# 0.5549f
C2093 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 a_20823_20174# 0.06243f
C2094 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 1.3467f
C2095 a_1896_19053# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 0.13749f
C2096 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.70899f
C2097 a_43698_7786# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.06167f
C2098 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_final_switch_0.VOUT[2] 0.01317f
C2099 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 15.9041f
C2100 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 a_27344_6250# 0.04213f
C2101 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.26041f
C2102 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.28795f
C2103 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.04811f
C2104 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_2678_10974# 0.04394f
C2105 VDDH a_14607_6250# 0.75085f
C2106 VDDH a_9353_15057# 0.49783f
C2107 a_15066_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.15182f
C2108 a_28172_6250# a_30608_7686# 0.03909f
C2109 a_28606_6250# a_30332_7686# 0.0396f
C2110 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.20199f
C2111 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 a_20823_20174# 0.06398f
C2112 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN a_5642_11461# 0.01003f
C2113 a_11629_15057# top_DAC_0/top_final_switch_0.VOUT[3] 0.01175f
C2114 a_23859_20174# a_22479_20174# 0.1541f
C2115 a_24411_20174# a_21927_20174# 0.1323f
C2116 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 a_27620_6250# 0.03927f
C2117 a_22469_18133# a_23307_20174# 0.06766f
C2118 a_23049_18133# a_23031_20174# 0.04294f
C2119 a_24135_20174# a_22203_20174# 0.13238f
C2120 a_23583_20174# a_22755_20174# 0.13293f
C2121 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.02801f
C2122 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.05944f
C2123 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.01222f
C2124 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.02785f
C2125 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.18261f
C2126 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.04864f
C2127 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 0.25806f
C2128 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.0486f
C2129 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43698_16696# 0.07243f
C2130 a_44062_19161# a_44062_18805# 0.04238f
C2131 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.77656f
C2132 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.02136f
C2133 a_15863_13785# a_15863_13536# 0.23441f
C2134 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_34856_8950# 0.11524f
C2135 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.47318f
C2136 a_43698_12736# a_43698_11746# 0.01563f
C2137 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.11733f
C2138 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 0.06082f
C2139 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.03939f
C2140 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.01844f
C2141 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.10148f
C2142 a_33910_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.12694f
C2143 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC a_39306_20477# 0.26172f
C2144 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_final_switch_0.VOUT[3] 0.10582f
C2145 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A a_43724_7946# 0.08029f
C2146 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_final_switch_0.VOUT[3] 0.20319f
C2147 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.0505f
C2148 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.9653f
C2149 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.02839f
C2150 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.20918f
C2151 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.03446f
C2152 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.13975f
C2153 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 0.03662f
C2154 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.0954f
C2155 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 1.31906f
C2156 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.18203f
C2157 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.90751f
C2158 a_30056_7686# a_27896_6250# 0.02791f
C2159 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB VDD 0.64193f
C2160 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.04788f
C2161 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.02254f
C2162 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.05177f
C2163 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 1.38015f
C2164 a_15863_13287# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.16718f
C2165 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.10707f
C2166 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C2167 VDDH a_5642_9535# 0.79462f
C2168 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_final_switch_0.VOUT[2] 0.01859f
C2169 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.05362f
C2170 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.05175f
C2171 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.04304f
C2172 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y a_44255_4078# 0.01129f
C2173 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.0163f
C2174 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.01836f
C2175 VOUT top_DAC_0/top_final_switch_0.VOUT[4] 8.15099f
C2176 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.23878f
C2177 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 1.46307f
C2178 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.12879f
C2179 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_final_switch_0.VOUT[3] 0.17157f
C2180 a_43698_6796# a_44234_7352# 0.07082f
C2181 a_16891_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.07419f
C2182 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A a_43724_7392# 0.03253f
C2183 a_19276_8950# a_19946_8950# 0.0895f
C2184 a_17148_18696# a_20547_20174# 0.02881f
C2185 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 2.13767f
C2186 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 a_14055_6250# 0.02784f
C2187 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 8.29955f
C2188 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.08386f
C2189 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 0.17836f
C2190 DIN3 VDDH 0.42749f
C2191 a_6445_15057# top_DAC_0/top_final_switch_0.VOUT[1] 0.03029f
C2192 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 1.27523f
C2193 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_final_switch_0.VOUT[3] 0.01686f
C2194 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 1.91899f
C2195 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_15272# 0.02704f
C2196 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.02047f
C2197 a_44234_12302# a_44234_12936# 0.02262f
C2198 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 1.3027f
C2199 a_15066_18696# a_14948_18696# 0.07321f
C2200 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.18999f
C2201 a_15342_18696# a_15224_18696# 0.07133f
C2202 a_14790_18696# a_14672_18696# 0.07191f
C2203 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.14544f
C2204 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.10119f
C2205 a_38584_20665# a_37410_19098# 0.01967f
C2206 a_23049_18133# a_23583_20174# 0.04025f
C2207 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 VDDH 0.0402f
C2208 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.04198f
C2209 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 a_15593_6250# 0.07771f
C2210 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.29339f
C2211 a_15593_6250# a_15353_7686# 0.04241f
C2212 a_15317_6250# a_15629_7686# 0.02803f
C2213 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.5492f
C2214 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.03397f
C2215 a_35757_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.26012f
C2216 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.06095f
C2217 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.5188f
C2218 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_16896# 0.14503f
C2219 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.08425f
C2220 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[3] 0.39596f
C2221 VDDH top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.39611f
C2222 a_24135_20174# a_24209_18133# 0.06779f
C2223 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN a_44234_7352# 0.06676f
C2224 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.08427f
C2225 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.05183f
C2226 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 2.09546f
C2227 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 1.29039f
C2228 a_34856_8950# a_29158_6250# 0.0394f
C2229 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN a_44234_13292# 0.08828f
C2230 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.11049f
C2231 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.09497f
C2232 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD 0.21618f
C2233 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.07123f
C2234 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.11032f
C2235 a_44062_20585# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.06327f
C2236 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.02784f
C2237 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.06812f
C2238 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.13214f
C2239 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_39936_22083# 0.5803f
C2240 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB VDD 1.19559f
C2241 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] VDD 1.24016f
C2242 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.15175f
C2243 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 a_28882_6250# 0.03939f
C2244 a_18008_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.26678f
C2245 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.16543f
C2246 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_21375_20174# 0.20237f
C2247 a_24963_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.21466f
C2248 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.08314f
C2249 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15869_6250# 0.18546f
C2250 VDDH a_19276_8950# 0.31885f
C2251 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 a_8506_12595# 1.6476f
C2252 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.24261f
C2253 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.25253f
C2254 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02788f
C2255 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.5557f
C2256 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_13926# 0.03152f
C2257 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.21415f
C2258 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.20842f
C2259 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.26895f
C2260 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.54094f
C2261 VDDH a_16181_7686# 0.45072f
C2262 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_18284_18696# 0.27182f
C2263 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_31870_7686# 0.11685f
C2264 a_19468_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.13822f
C2265 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 0.31595f
C2266 a_4415_23194# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.0184f
C2267 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.10492f
C2268 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.17603f
C2269 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.62948f
C2270 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 3.15778f
C2271 a_5642_11461# a_5642_10963# 0.015f
C2272 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09271f
C2273 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 a_16872_18696# 0.03988f
C2274 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.48595f
C2275 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.11132f
C2276 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] VDDH 0.01046f
C2277 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_23629_18133# 0.05861f
C2278 a_20076_10031# a_20656_10031# 0.05093f
C2279 a_19772_10031# a_20932_10031# 0.10606f
C2280 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 a_29780_7686# 0.04526f
C2281 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.0245f
C2282 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.18775f
C2283 a_18284_18696# top_DAC_0/top_rseg_n_dcell_0.VL3 0.40158f
C2284 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.05635f
C2285 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.05996f
C2286 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.12671f
C2287 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 a_13779_6250# 0.04213f
C2288 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.15469f
C2289 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 0.01575f
C2290 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.15972f
C2291 a_44234_11946# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.08412f
C2292 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.VS1 0.04547f
C2293 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 VDDH 0.36689f
C2294 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] ROUT2 0.06337f
C2295 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.69667f
C2296 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.15152f
C2297 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 0.13263f
C2298 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 25.2932f
C2299 a_34873_10031# a_34569_10031# 0.71565f
C2300 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.02015f
C2301 top_DAC_0/top_rseg_n_dcell_0.VL2 a_14615_13785# 0.04346f
C2302 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.08682f
C2303 a_35177_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.33041f
C2304 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_44062_20229# 0.06327f
C2305 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 a_28606_6250# 0.11045f
C2306 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_final_switch_0.VOUT[0] 0.05663f
C2307 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.07353f
C2308 a_35757_10031# a_34856_8950# 0.06662f
C2309 a_35453_10031# a_35132_8950# 0.08323f
C2310 a_33358_8950# a_34304_8950# 0.09145f
C2311 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_final_switch_0.VOUT[4] 0.01346f
C2312 a_36033_10031# a_34580_8950# 0.06546f
C2313 a_15098_19866# a_15224_18696# 0.26978f
C2314 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 1.98281f
C2315 a_44234_11946# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.03152f
C2316 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 a_30332_7686# 0.07456f
C2317 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.16949f
C2318 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.0921f
C2319 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_19946_8950# 0.11896f
C2320 a_34580_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.01661f
C2321 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_44062_21297# 0.02123f
C2322 VDDH a_43724_6956# 0.09226f
C2323 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB a_44234_6996# 0.13692f
C2324 a_16320_18696# a_16596_18696# 1.86139f
C2325 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.VS1 0.27984f
C2326 a_14672_18696# a_16872_18696# 0.08905f
C2327 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.1676f
C2328 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_15906# 0.03855f
C2329 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.09158f
C2330 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.0481f
C2331 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 a_15224_18696# 0.06354f
C2332 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV VDDH 1.06415f
C2333 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 0.32173f
C2334 a_34856_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.19575f
C2335 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.08272f
C2336 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP a_43698_11746# 0.02263f
C2337 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A VDD 0.32055f
C2338 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.17446f
C2339 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 0.84969f
C2340 a_43724_11352# VDDH 0.09227f
C2341 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_10322# 0.0248f
C2342 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.08478f
C2343 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.88718f
C2344 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.09426f
C2345 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.01131f
C2346 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.07181f
C2347 top_DAC_0/top_final_switch_0.VOUT[3] a_11081_14150# 0.01871f
C2348 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 15.6649f
C2349 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.84443f
C2350 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.09128f
C2351 a_15863_13785# top_DAC_0/top_final_switch_0.VOUT[4] 0.03215f
C2352 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.05383f
C2353 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y a_45023_19988# 0.01005f
C2354 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.09535f
C2355 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_16320_18696# 0.20514f
C2356 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 1.2875f
C2357 a_22755_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 0.04143f
C2358 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.06351f
C2359 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_31870_7686# 0.14673f
C2360 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 1.78008f
C2361 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_19670_8950# 0.01313f
C2362 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 a_21375_20174# 0.0516f
C2363 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 a_21099_20174# 0.06393f
C2364 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.09946f
C2365 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01021f
C2366 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.09461f
C2367 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.14522f
C2368 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 0.9083f
C2369 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 a_28882_6250# 0.02791f
C2370 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_7986# 0.01484f
C2371 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.33687f
C2372 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 0.21449f
C2373 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.09513f
C2374 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_31042_7686# 0.07726f
C2375 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.01745f
C2376 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.05838f
C2377 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 a_28172_6250# 0.04331f
C2378 a_17443_7686# a_20222_8950# 0.07934f
C2379 a_15863_13536# top_DAC_0/top_final_switch_0.VOUT[1] 0.07667f
C2380 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 a_29158_6250# 0.02801f
C2381 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 a_29434_6250# 0.03927f
C2382 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 0.05194f
C2383 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_2300_15118# 0.04824f
C2384 VDDH a_5050_12595# 0.01047f
C2385 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.2707f
C2386 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 2.01688f
C2387 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.16626f
C2388 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.06054f
C2389 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB DIN3 0.17953f
C2390 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.33138f
C2391 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_21651_20174# 0.03231f
C2392 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 1.23034f
C2393 a_15342_18696# a_17732_18696# 0.2541f
C2394 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 0.13356f
C2395 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 0.15193f
C2396 a_15066_18696# a_18008_18696# 0.62343f
C2397 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.03539f
C2398 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 1.27501f
C2399 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 a_27620_6250# 0.07808f
C2400 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_final_switch_0.VOUT[3] 0.02123f
C2401 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.68733f
C2402 a_15593_6250# a_16891_7686# 0.02794f
C2403 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_5897_12507# 0.0208f
C2404 a_15317_6250# a_17167_7686# 0.02809f
C2405 a_15869_6250# a_16615_7686# 0.03863f
C2406 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 0.05959f
C2407 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 2.7521f
C2408 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.05506f
C2409 a_31042_7686# a_31594_7686# 0.16691f
C2410 a_30608_7686# a_31870_7686# 0.17976f
C2411 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.46005f
C2412 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.0483f
C2413 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_15863_13536# 0.01107f
C2414 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.VS4 0.0322f
C2415 a_4717_15057# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.01033f
C2416 a_43698_14716# a_44234_15272# 0.07082f
C2417 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_28882_6250# 0.40634f
C2418 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44062_18449# 0.02511f
C2419 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 0.11411f
C2420 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.19037f
C2421 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3 0.04143f
C2422 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.12629f
C2423 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.01782f
C2424 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.13341f
C2425 VOUT a_11629_14150# 0.0409f
C2426 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.02715f
C2427 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.21426f
C2428 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 0.02026f
C2429 a_15863_13536# top_DAC_0/top_rseg_n_dcell_0.VL3 0.17548f
C2430 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.08824f
C2431 a_21651_20174# a_23307_20174# 0.1769f
C2432 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 a_16320_18696# 0.09568f
C2433 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 0.73274f
C2434 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 0.55355f
C2435 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_6445_12507# 0.02171f
C2436 a_8051_10107# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.78597f
C2437 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.77409f
C2438 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_23307_20174# 0.02886f
C2439 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.04093f
C2440 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 0.40134f
C2441 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_6923_9707# 2.13138f
C2442 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.04186f
C2443 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.26869f
C2444 top_DAC_0/top_final_switch_0.VOUT[0] a_5897_15057# 0.03805f
C2445 DIN8 DIN9 0.33674f
C2446 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 1.58886f
C2447 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 0.05546f
C2448 VDDH top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A 3.88898f
C2449 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 4.55333f
C2450 a_20498_8950# a_18724_8950# 0.16175f
C2451 a_7625_14150# VOUT 0.06741f
C2452 a_20222_8950# a_19000_8950# 0.08868f
C2453 top_DAC_0/top_final_switch_0.VOUT[1] a_7625_15057# 0.03805f
C2454 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 a_21927_20174# 0.04145f
C2455 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_16615_7686# 0.11949f
C2456 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 a_27896_6250# 0.038f
C2457 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.20513f
C2458 a_8506_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.17245f
C2459 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD 0.21631f
C2460 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_30332_7686# 0.11409f
C2461 a_44234_7986# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.06901f
C2462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_2678_10974# 0.02444f
C2463 VDDH a_27344_6250# 0.01731f
C2464 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.05973f
C2465 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 a_28172_6250# 0.03732f
C2466 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_1896_12504# 0.01649f
C2467 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.02163f
C2468 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.58839f
C2469 VDDH a_14948_18696# 0.30303f
C2470 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB a_44234_7986# 0.21463f
C2471 a_34186_8950# a_34304_8950# 3.2779f
C2472 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.3001f
C2473 a_33910_8950# a_34580_8950# 0.0895f
C2474 a_33634_8950# a_34856_8950# 0.08868f
C2475 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 0.06041f
C2476 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.04795f
C2477 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 1.16723f
C2478 a_35132_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.23586f
C2479 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.08189f
C2480 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 0.15608f
C2481 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.07862f
C2482 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 1.916f
C2483 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.18208f
C2484 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.02737f
C2485 a_38617_19854# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.01035f
C2486 a_15353_7686# a_13779_6250# 0.04585f
C2487 a_15593_6250# a_14331_6250# 0.15321f
C2488 a_30332_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.02941f
C2489 a_15869_6250# a_14055_6250# 0.17253f
C2490 a_15317_6250# a_14607_6250# 0.17893f
C2491 a_23031_20174# a_23307_20174# 0.89932f
C2492 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 0.1166f
C2493 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.14754f
C2494 top_DAC_0/top_rseg_n_dcell_0.VH3 a_18284_18696# 0.17595f
C2495 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 16.1091f
C2496 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.05628f
C2497 a_38672_20477# a_39768_20665# 0.01967f
C2498 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] a_16320_18696# 0.02168f
C2499 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 a_15593_6250# 0.02801f
C2500 a_14514_18696# a_14790_18696# 1.81369f
C2501 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN DIN1 0.03521f
C2502 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.01753f
C2503 a_24135_20174# a_21375_20174# 0.14456f
C2504 a_24411_20174# a_21099_20174# 0.13227f
C2505 a_24963_20174# a_20547_20174# 0.25578f
C2506 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.07096f
C2507 a_24687_20174# a_20823_20174# 0.13259f
C2508 a_23859_20174# a_21651_20174# 0.15679f
C2509 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.35811f
C2510 a_31318_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.03948f
C2511 a_39768_20389# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.02668f
C2512 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.06295f
C2513 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.14826f
C2514 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD VOUT 0.67332f
C2515 a_15353_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.5644f
C2516 a_15098_19866# a_17732_18696# 0.01367f
C2517 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.23555f
C2518 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_15593_6250# 0.44165f
C2519 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.22293f
C2520 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 1.73509f
C2521 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.48789f
C2522 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_5642_10963# 0.01106f
C2523 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04845f
C2524 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.05552f
C2525 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_15906# 0.14379f
C2526 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB VDD 0.32717f
C2527 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.10073f
C2528 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 0.06569f
C2529 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.02792f
C2530 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.0921f
C2531 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 0.0953f
C2532 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.01165f
C2533 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 1.28515f
C2534 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.04626f
C2535 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 1.06014f
C2536 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 0.27414f
C2537 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_15866# 0.03597f
C2538 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.1143f
C2539 top_DAC_0/top_rseg_n_dcell_0.VH2 VDDH 0.20437f
C2540 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_14282# 0.03855f
C2541 a_1896_17510# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 0.01034f
C2542 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 a_16891_7686# 0.03991f
C2543 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 a_23031_20174# 0.064f
C2544 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_14055_6250# 0.26602f
C2545 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44062_21653# 0.0205f
C2546 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.05544f
C2547 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_10322# 0.14048f
C2548 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.04852f
C2549 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 a_27896_6250# 0.02788f
C2550 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 0.05177f
C2551 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_5111_10963# 0.0135f
C2552 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.11733f
C2553 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 0.21283f
C2554 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04064f
C2555 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 a_27344_6250# 0.05951f
C2556 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.03198f
C2557 a_15618_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.48017f
C2558 VDDH a_9353_14150# 0.49013f
C2559 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 0.08663f
C2560 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 0.16825f
C2561 a_28172_6250# a_31318_7686# 0.04373f
C2562 a_28882_6250# a_30608_7686# 0.02798f
C2563 a_28606_6250# a_31042_7686# 0.04804f
C2564 a_29158_6250# a_30332_7686# 0.02791f
C2565 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.2482f
C2566 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.08341f
C2567 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.17102f
C2568 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 a_23031_20174# 0.06393f
C2569 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.03142f
C2570 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.31212f
C2571 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.VL3 0.06558f
C2572 a_24135_20174# a_22755_20174# 0.13273f
C2573 a_24687_20174# a_22203_20174# 0.13261f
C2574 a_24411_20174# a_22479_20174# 0.13264f
C2575 a_23859_20174# a_23031_20174# 0.1525f
C2576 a_24963_20174# a_21927_20174# 0.13259f
C2577 a_23583_20174# a_23307_20174# 0.60366f
C2578 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_19552_8950# 0.20678f
C2579 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.17254f
C2580 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 a_15593_6250# 0.02785f
C2581 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.02786f
C2582 a_38672_20477# a_39306_20477# 0.20495f
C2583 a_38584_20389# a_38584_20665# 0.02286f
C2584 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 0.90195f
C2585 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 0.01777f
C2586 VDDH a_9901_15057# 0.49792f
C2587 a_15863_13536# a_15863_13287# 0.21795f
C2588 a_15863_13785# top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.07888f
C2589 a_15618_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.01189f
C2590 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 6.01491f
C2591 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.11848f
C2592 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_15312# 0.03597f
C2593 a_34304_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.09341f
C2594 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 10.5012f
C2595 a_11629_15057# top_DAC_0/top_final_switch_0.VOUT[4] 0.03029f
C2596 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.90617f
C2597 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04939f
C2598 top_DAC_0/top_final_switch_0.VOUT[2] a_8506_12595# 0.43678f
C2599 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 4.16288f
C2600 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.38211f
C2601 a_44234_9332# a_44234_8976# 0.08026f
C2602 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 1.34685f
C2603 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.12314f
C2604 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 0.05271f
C2605 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] a_15224_18696# 0.11401f
C2606 a_17148_18696# a_14948_18696# 0.09851f
C2607 VDDH a_5642_8388# 0.72861f
C2608 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_37804_20713# 0.0211f
C2609 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.12689f
C2610 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.02786f
C2611 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.19452f
C2612 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 0.80848f
C2613 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.02788f
C2614 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_final_switch_0.VOUT[4] 0.11625f
C2615 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_final_switch_0.VOUT[4] 0.07919f
C2616 a_16891_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.03948f
C2617 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 1.15703f
C2618 VDDH VOUT 8.72574f
C2619 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A a_44234_6996# 0.05897f
C2620 a_19276_8950# a_20498_8950# 0.10102f
C2621 a_43698_6796# a_43724_6956# 0.02395f
C2622 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.02785f
C2623 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.68535f
C2624 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_final_switch_0.VOUT[2] 0.01788f
C2625 a_5050_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.09303f
C2626 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 a_14607_6250# 0.02784f
C2627 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_43698_6796# 0.24498f
C2628 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04834f
C2629 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.93455f
C2630 a_15863_13536# top_DAC_0/top_rseg_n_dcell_0.VH3 0.04213f
C2631 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 0.3191f
C2632 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.02795f
C2633 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.03935f
C2634 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_final_switch_0.VOUT[4] 0.04554f
C2635 a_37410_19098# a_39306_20477# 0.21877f
C2636 a_22469_18133# a_24411_20174# 0.04028f
C2637 a_23583_20174# a_23859_20174# 0.33401f
C2638 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.08622f
C2639 a_15869_6250# a_15629_7686# 0.04338f
C2640 a_15317_6250# a_16181_7686# 0.028f
C2641 a_15593_6250# a_15905_7686# 0.02792f
C2642 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 3.65825f
C2643 a_43698_13726# a_43724_14322# 0.06762f
C2644 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_20352_10031# 0.21608f
C2645 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_8342# 0.01743f
C2646 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_14916# 0.03152f
C2647 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_43698_15706# 0.24618f
C2648 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.02209f
C2649 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.02791f
C2650 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_8506_12595# 0.26324f
C2651 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_24963_20174# 0.01066f
C2652 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_final_switch_0.VOUT[4] 0.02878f
C2653 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 0.30567f
C2654 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.04862f
C2655 a_24687_20174# a_24209_18133# 0.06784f
C2656 a_30332_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.06223f
C2657 a_36813_19760# a_36888_19786# 0.04493f
C2658 VDDH a_18008_18696# 0.24564f
C2659 a_14615_14034# top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.05501f
C2660 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_14790_18696# 0.0594f
C2661 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.11733f
C2662 a_35132_8950# a_29434_6250# 0.03993f
C2663 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.44293f
C2664 a_7625_13005# a_8173_13005# 0.0103f
C2665 DIN8 DIN7 0.33719f
C2666 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.17417f
C2667 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 a_15317_6250# 0.02791f
C2668 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 a_31870_7686# 0.03929f
C2669 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 a_15317_6250# 0.03878f
C2670 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.0126f
C2671 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.04506f
C2672 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 0.50237f
C2673 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.03837f
C2674 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.98671f
C2675 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 0.47118f
C2676 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 1.34913f
C2677 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.02784f
C2678 a_13779_6250# a_16891_7686# 0.03171f
C2679 a_14055_6250# a_16615_7686# 0.02789f
C2680 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.02427f
C2681 DIN4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.17948f
C2682 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 1.24832f
C2683 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_39861_21457# 0.06598f
C2684 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 1.42737f
C2685 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 1.9603f
C2686 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.09964f
C2687 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 0.11559f
C2688 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 0.25566f
C2689 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 0.05773f
C2690 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[4] 0.31502f
C2691 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 0.05286f
C2692 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.06329f
C2693 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] ROUT2 0.01445f
C2694 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 1.34056f
C2695 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP 0.92832f
C2696 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04794f
C2697 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.0279f
C2698 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 8.86068f
C2699 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15629_7686# 0.13166f
C2700 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02791f
C2701 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 1.57251f
C2702 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 1.17367f
C2703 a_1896_20320# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 0.06418f
C2704 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.03545f
C2705 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 17.3149f
C2706 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.01643f
C2707 a_16891_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.07264f
C2708 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB a_44234_8976# 0.28536f
C2709 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.10107f
C2710 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.20881f
C2711 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.19454f
C2712 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.05042f
C2713 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_9353_14150# 0.04959f
C2714 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.048f
C2715 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.09704f
C2716 a_30332_7686# a_27344_6250# 0.03759f
C2717 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.08134f
C2718 VOUT a_11081_13005# 0.02203f
C2719 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.02024f
C2720 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.03641f
C2721 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 0.04287f
C2722 a_20352_10031# a_20932_10031# 0.05788f
C2723 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 0.08581f
C2724 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_7352# 0.01481f
C2725 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.1884f
C2726 a_44062_20585# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.02575f
C2727 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.02788f
C2728 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 a_30608_7686# 0.03929f
C2729 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_14282# 0.14379f
C2730 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.04456f
C2731 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 a_14331_6250# 0.02788f
C2732 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP a_43724_15312# 0.03147f
C2733 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 0.13284f
C2734 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 a_21651_20174# 0.06393f
C2735 a_35453_10031# a_34569_10031# 0.38399f
C2736 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_20547_20174# 0.03043f
C2737 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_44062_19517# 0.06327f
C2738 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_23307_20174# 0.03149f
C2739 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.11272f
C2740 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.06065f
C2741 a_4415_23194# a_8473_23194# 0.42742f
C2742 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 0.02582f
C2743 DIN6 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.17939f
C2744 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.0532f
C2745 a_15374_19866# a_14948_18696# 0.09179f
C2746 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.03344f
C2747 a_15098_19866# a_14672_18696# 0.2153f
C2748 a_33358_8950# a_34856_8950# 0.0996f
C2749 a_36033_10031# a_35132_8950# 0.02529f
C2750 a_43698_10756# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.01234f
C2751 a_13779_6250# a_14331_6250# 0.19435f
C2752 a_44737_4828# VDD 0.02571f
C2753 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_20498_8950# 0.11687f
C2754 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.VH3 0.05787f
C2755 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.10742f
C2756 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 a_31318_7686# 0.03948f
C2757 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.04637f
C2758 VDDH top_DAC_0/top_rseg_n_dcell_0.SH[1] 1.78593f
C2759 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 1.70953f
C2760 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 1.06161f
C2761 a_16596_18696# a_16872_18696# 1.8469f
C2762 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.10024f
C2763 a_4717_15057# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.04959f
C2764 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C2765 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 0.03971f
C2766 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_43698_11746# 0.24498f
C2767 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB VOUT 3.98706f
C2768 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 0.05997f
C2769 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.09836f
C2770 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 a_13779_6250# 0.055f
C2771 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.05371f
C2772 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.03944f
C2773 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 a_16181_7686# 0.03955f
C2774 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_20352_10031# 0.06447f
C2775 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 0.279f
C2776 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.96668f
C2777 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_7392# 0.03597f
C2778 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 0.01396f
C2779 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.21565f
C2780 a_37277_19098# a_37410_19098# 0.02707f
C2781 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] DIN8 0.0349f
C2782 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.0203f
C2783 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.02179f
C2784 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.02194f
C2785 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_13779_6250# 0.77109f
C2786 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44062_20229# 0.0242f
C2787 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_16872_18696# 0.2298f
C2788 a_44062_20585# a_44062_20229# 0.04238f
C2789 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_20222_8950# 0.08905f
C2790 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 1.78725f
C2791 a_43698_8776# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.78464f
C2792 a_43698_10756# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.06167f
C2793 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.17015f
C2794 VDDH a_15863_13785# 0.1926f
C2795 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.04736f
C2796 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.02181f
C2797 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.2275f
C2798 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 0.10095f
C2799 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 a_14331_6250# 0.03957f
C2800 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.0256f
C2801 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.13238f
C2802 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 a_29434_6250# 0.04267f
C2803 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_31594_7686# 0.07546f
C2804 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 a_28882_6250# 0.04196f
C2805 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.11466f
C2806 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 1.61573f
C2807 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 3.18174f
C2808 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_final_switch_0.VOUT[1] 0.06657f
C2809 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.22936f
C2810 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_2300_14353# 0.04784f
C2811 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 0.0616f
C2812 a_23859_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.02856f
C2813 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 1.17003f
C2814 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 1.71248f
C2815 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 15.5261f
C2816 a_15618_18696# a_18008_18696# 0.37273f
C2817 a_15342_18696# a_18284_18696# 0.03043f
C2818 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.02339f
C2819 VDDH a_11081_15057# 0.49886f
C2820 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04846f
C2821 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 0.14638f
C2822 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 0.01875f
C2823 a_16181_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.03955f
C2824 a_15353_7686# a_16891_7686# 0.20414f
C2825 a_15593_6250# a_17443_7686# 0.04806f
C2826 a_15629_7686# a_16615_7686# 0.16668f
C2827 a_15869_6250# a_17167_7686# 0.03867f
C2828 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 0.05755f
C2829 a_44234_13292# a_44234_13926# 0.02262f
C2830 a_20547_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 0.01567f
C2831 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_8342# 0.1344f
C2832 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 9.60185f
C2833 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 a_13779_6250# 0.04219f
C2834 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.17416f
C2835 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 4.05624f
C2836 a_31318_7686# a_31870_7686# 0.18799f
C2837 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.13425f
C2838 top_DAC_0/top_final_switch_0.VOUT[4] a_12809_15057# 0.03952f
C2839 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 VDDH 0.16077f
C2840 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_29434_6250# 0.41121f
C2841 a_43698_14716# a_43724_14876# 0.02395f
C2842 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP a_44234_14916# 0.06668f
C2843 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.04783f
C2844 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_12504# 0.05618f
C2845 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_final_switch_0.VOUT[4] 0.03086f
C2846 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.01335f
C2847 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 0.48841f
C2848 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.06115f
C2849 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 0.76371f
C2850 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD a_6445_15057# 0.01033f
C2851 top_DAC_0/top_rseg_n_dcell_0.VH2 a_22193_18133# 0.1537f
C2852 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.VL3 0.20205f
C2853 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.13152f
C2854 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.22605f
C2855 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.01649f
C2856 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.04978f
C2857 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.01121f
C2858 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.19295f
C2859 a_44234_9966# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.06749f
C2860 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.12567f
C2861 a_11081_12507# a_11629_12507# 0.0103f
C2862 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_final_switch_0.VOUT[3] 0.01859f
C2863 a_19552_8950# a_19670_8950# 3.08648f
C2864 a_2678_10974# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.02385f
C2865 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04695f
C2866 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 0.0556f
C2867 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.03653f
C2868 a_44234_7352# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.06328f
C2869 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.09546f
C2870 top_DAC_0/top_final_switch_0.VOUT[0] a_5897_14150# 0.01852f
C2871 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.12695f
C2872 DIN0 DIN1 0.32901f
C2873 a_15629_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.07245f
C2874 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 0.01814f
C2875 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_final_switch_0.VOUT[1] 0.16754f
C2876 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.26402f
C2877 top_DAC_0/top_final_switch_0.VOUT[1] a_7625_14150# 0.01864f
C2878 VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.03004f
C2879 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.11848f
C2880 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_17167_7686# 0.11901f
C2881 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 a_15905_7686# 0.07456f
C2882 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.05884f
C2883 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.04219f
C2884 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.05944f
C2885 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_31042_7686# 0.11496f
C2886 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.08546f
C2887 a_1896_16243# a_2678_16243# 0.02127f
C2888 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.04106f
C2889 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.17825f
C2890 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.08793f
C2891 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.05305f
C2892 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.26638f
C2893 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 0.02078f
C2894 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 1.58612f
C2895 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.049f
C2896 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.05356f
C2897 DIN6 DIN7 0.33364f
C2898 a_15869_6250# a_18724_8950# 0.02235f
C2899 VDDH a_16320_18696# 0.27916f
C2900 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 0.01852f
C2901 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_1896_11886# 0.02524f
C2902 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 a_28882_6250# 0.03894f
C2903 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 1.89276f
C2904 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 0.01836f
C2905 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 1.47954f
C2906 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.055f
C2907 a_34186_8950# a_34856_8950# 0.08994f
C2908 a_33910_8950# a_35132_8950# 0.10159f
C2909 a_34304_8950# a_34580_8950# 3.17836f
C2910 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 a_28172_6250# 0.02791f
C2911 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.01812f
C2912 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.09934f
C2913 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.43907f
C2914 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04903f
C2915 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 0.38473f
C2916 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.05053f
C2917 a_15869_6250# a_14607_6250# 0.18306f
C2918 a_15629_7686# a_14055_6250# 0.02786f
C2919 a_15353_7686# a_14331_6250# 0.0421f
C2920 a_15593_6250# a_15041_6250# 0.16898f
C2921 a_37737_19479# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.02737f
C2922 a_15905_7686# a_13779_6250# 0.03168f
C2923 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_15272# 0.03855f
C2924 a_31042_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.02804f
C2925 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.02388f
C2926 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 0.48684f
C2927 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.11045f
C2928 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.05514f
C2929 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP 0.01782f
C2930 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.96691f
C2931 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.VL3 0.03391f
C2932 a_38672_20477# a_39768_20389# 0.01857f
C2933 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 0.86278f
C2934 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.02493f
C2935 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.02615f
C2936 a_14790_18696# a_15066_18696# 1.82015f
C2937 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 a_31594_7686# 0.03929f
C2938 a_14514_18696# a_15342_18696# 0.09822f
C2939 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.1308f
C2940 a_23859_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 0.05531f
C2941 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] VDDH 0.88394f
C2942 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 18.3073f
C2943 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.01651f
C2944 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 0.04264f
C2945 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.89962f
C2946 a_24411_20174# a_21651_20174# 0.13222f
C2947 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 0.1321f
C2948 a_24963_20174# a_21099_20174# 0.13245f
C2949 a_24687_20174# a_21375_20174# 0.146f
C2950 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.04851f
C2951 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.2548f
C2952 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.11409f
C2953 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_8173_13005# 0.0208f
C2954 a_15905_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.07894f
C2955 a_22193_18133# a_22469_18133# 4.14664f
C2956 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 1.83395f
C2957 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.01647f
C2958 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_28606_6250# 0.15698f
C2959 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 2.32271f
C2960 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_18724_8950# 0.03789f
C2961 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.32075f
C2962 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.32371f
C2963 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_15353_7686# 0.49776f
C2964 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.10925f
C2965 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 0.07865f
C2966 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.02797f
C2967 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 0.15788f
C2968 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.02514f
C2969 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.28713f
C2970 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 1.07647f
C2971 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.02789f
C2972 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 0.0142f
C2973 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP 0.3001f
C2974 top_DAC_0/top_rseg_n_dcell_0.VL2 a_24209_18133# 0.12882f
C2975 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.07f
C2976 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.08957f
C2977 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 3.60244f
C2978 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09038f
C2979 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.03404f
C2980 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_14607_6250# 0.23478f
C2981 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.01392f
C2982 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 8.75672f
C2983 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 a_27620_6250# 0.02803f
C2984 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 0.09515f
C2985 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.37729f
C2986 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 2.8803f
C2987 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.05459f
C2988 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.02163f
C2989 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 a_27896_6250# 0.02788f
C2990 a_44234_10956# a_44234_10322# 0.02262f
C2991 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.17797f
C2992 a_29780_7686# a_30332_7686# 0.20828f
C2993 a_29158_6250# a_31042_7686# 0.02792f
C2994 a_28172_6250# a_31870_7686# 0.12966f
C2995 a_29434_6250# a_30608_7686# 0.04155f
C2996 a_28606_6250# a_31594_7686# 0.06225f
C2997 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.15063f
C2998 a_28882_6250# a_31318_7686# 0.02801f
C2999 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 a_22203_20174# 0.04147f
C3000 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_43698_8776# 0.24498f
C3001 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 0.06345f
C3002 a_23629_18133# a_24209_18133# 3.47409f
C3003 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.18654f
C3004 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.02445f
C3005 a_24135_20174# a_23307_20174# 0.12572f
C3006 a_24411_20174# a_23031_20174# 0.13437f
C3007 a_24963_20174# a_22479_20174# 0.13713f
C3008 a_24687_20174# a_22755_20174# 0.13502f
C3009 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.05431f
C3010 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.20774f
C3011 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_19946_8950# 0.20162f
C3012 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.04802f
C3013 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 0.02138f
C3014 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.06984f
C3015 a_15863_13287# top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.10915f
C3016 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.11049f
C3017 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09039f
C3018 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.14053f
C3019 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.10426f
C3020 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_27620_6250# 0.2146f
C3021 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.03915f
C3022 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_15317_6250# 0.14677f
C3023 a_34856_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.11689f
C3024 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 0.02568f
C3025 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.03397f
C3026 a_16615_7686# a_17167_7686# 0.16691f
C3027 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.18985f
C3028 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.01796f
C3029 VDDH a_11629_15057# 0.49751f
C3030 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.VS1 1.61787f
C3031 a_17148_18696# a_16320_18696# 0.09912f
C3032 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] a_14672_18696# 0.11614f
C3033 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02077f
C3034 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 a_15224_18696# 0.06345f
C3035 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.05175f
C3036 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 0.02063f
C3037 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_21375_20174# 0.08113f
C3038 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.02214f
C3039 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.22101f
C3040 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.03917f
C3041 a_35177_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05937f
C3042 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 a_15593_6250# 0.02933f
C3043 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.09522f
C3044 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 1.34563f
C3045 VDDH top_DAC_0/top_final_switch_0.VOUT[1] 1.66034f
C3046 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 2.32693f
C3047 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.02537f
C3048 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.06345f
C3049 a_15098_19866# a_14514_18696# 0.04604f
C3050 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.01148f
C3051 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_14615_14283# 0.07377f
C3052 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 4.38923f
C3053 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN a_5642_9535# 0.01975f
C3054 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.32243f
C3055 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.65489f
C3056 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.08636f
C3057 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.15936f
C3058 a_15342_18696# a_16596_18696# 0.0652f
C3059 a_15066_18696# a_16872_18696# 0.06533f
C3060 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_8051_10107# 1.05749f
C3061 a_45343_4622# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.01243f
C3062 a_15618_18696# a_16320_18696# 0.06563f
C3063 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.07676f
C3064 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_15863_13287# 0.03169f
C3065 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN VDD 0.4425f
C3066 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.98493f
C3067 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.05178f
C3068 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.0433f
C3069 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.04707f
C3070 a_23583_20174# a_24411_20174# 5.48788f
C3071 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04361f
C3072 a_23859_20174# a_24135_20174# 5.86941f
C3073 a_22469_18133# a_24963_20174# 0.04042f
C3074 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_8173_15057# 0.04959f
C3075 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 a_28606_6250# 0.02791f
C3076 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.14095f
C3077 a_15353_7686# a_15905_7686# 0.20809f
C3078 a_15869_6250# a_16181_7686# 0.04152f
C3079 a_11629_14150# a_11081_14150# 0.0237f
C3080 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_20932_10031# 0.24632f
C3081 a_43698_13726# a_44234_13926# 0.0139f
C3082 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 VDDH 2.92054f
C3083 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 a_27344_6250# 0.0426f
C3084 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_5111_10963# 0.7841f
C3085 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.02794f
C3086 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.87726f
C3087 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.11733f
C3088 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.25891f
C3089 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.31218f
C3090 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04805f
C3091 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.64599f
C3092 a_31042_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.03243f
C3093 a_37595_19760# a_36888_19550# 0.01891f
C3094 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.02801f
C3095 VDDH top_DAC_0/top_rseg_n_dcell_0.VL3 0.57817f
C3096 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_15342_18696# 0.05514f
C3097 a_14615_13536# top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.10671f
C3098 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 1.82529f
C3099 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 1.31057f
C3100 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.19456f
C3101 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 a_15869_6250# 0.30093f
C3102 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 a_15869_6250# 0.04262f
C3103 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_27620_6250# 0.16757f
C3104 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_15272# 0.14379f
C3105 a_14055_6250# a_17167_7686# 0.02794f
C3106 a_14607_6250# a_16615_7686# 0.0397f
C3107 a_13779_6250# a_17443_7686# 0.04934f
C3108 a_14331_6250# a_16891_7686# 0.02796f
C3109 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 0.10239f
C3110 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B VDD 0.25715f
C3111 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.11902f
C3112 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 0.03652f
C3113 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.09709f
C3114 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.12293f
C3115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.14083f
C3116 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.02785f
C3117 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.0483f
C3118 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 1.1572f
C3119 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.48603f
C3120 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.29715f
C3121 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] DIN7 0.0349f
C3122 a_43698_12736# a_43724_13332# 0.06762f
C3123 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 0.50407f
C3124 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 0.05667f
C3125 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 0.82312f
C3126 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD a_7625_15057# 0.01033f
C3127 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.16361f
C3128 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 a_16891_7686# 0.07419f
C3129 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 17.3348f
C3130 a_28172_6250# a_28882_6250# 0.17811f
C3131 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.08425f
C3132 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.03122f
C3133 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 2.24695f
C3134 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.VH3 0.08714f
C3135 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.61812f
C3136 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_16181_7686# 0.12058f
C3137 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.24589f
C3138 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.07455f
C3139 a_1636_13352# VOUT 0.01053f
C3140 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.07155f
C3141 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_21375_20174# 0.08101f
C3142 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 3.73465f
C3143 a_17443_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.11293f
C3144 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 0.09136f
C3145 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.02717f
C3146 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_16891_7686# 0.07974f
C3147 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.08855f
C3148 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 a_16872_18696# 0.08386f
C3149 a_30332_7686# a_27896_6250# 0.02791f
C3150 a_30608_7686# a_27620_6250# 0.02788f
C3151 a_31042_7686# a_27344_6250# 0.0376f
C3152 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.10225f
C3153 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.32504f
C3154 a_6778_12595# a_8506_12595# 0.11851f
C3155 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 a_15317_6250# 0.04185f
C3156 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.68258f
C3157 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.03694f
C3158 VOUT a_11081_12507# 0.04471f
C3159 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.11186f
C3160 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_15863_13785# 0.14514f
C3161 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.01029f
C3162 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.04324f
C3163 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.09522f
C3164 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.72782f
C3165 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.0259f
C3166 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.02785f
C3167 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 a_15041_6250# 0.02791f
C3168 a_44234_7986# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.06548f
C3169 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.01514f
C3170 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_20352_10031# 0.17361f
C3171 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.11583f
C3172 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.38436f
C3173 a_14055_6250# a_18724_8950# 0.11111f
C3174 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_6996# 0.01554f
C3175 a_6923_9707# a_8051_10107# 0.15848f
C3176 a_31594_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.07153f
C3177 a_34569_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.13734f
C3178 VDDH a_1896_16243# 0.72203f
C3179 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.4555f
C3180 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 0.02449f
C3181 a_15098_19866# a_16596_18696# 0.10122f
C3182 a_15374_19866# a_16320_18696# 0.08856f
C3183 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.07771f
C3184 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.05434f
C3185 a_1896_19053# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 0.03145f
C3186 a_13779_6250# a_15041_6250# 0.20977f
C3187 a_14055_6250# a_14607_6250# 0.16227f
C3188 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.10655f
C3189 a_44062_18093# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.02123f
C3190 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.03612f
C3191 a_14790_18696# VDDH 0.27361f
C3192 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.0405f
C3193 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 2.66628f
C3194 a_17148_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.01386f
C3195 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.05653f
C3196 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 a_29158_6250# 0.07764f
C3197 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_final_switch_0.VOUT[2] 0.05518f
C3198 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 0.05852f
C3199 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.02255f
C3200 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 a_28606_6250# 0.03939f
C3201 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_final_switch_0.VOUT[1] 0.20373f
C3202 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 a_14331_6250# 0.02788f
C3203 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_20932_10031# 0.06163f
C3204 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 1.31964f
C3205 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.14755f
C3206 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y a_45343_4828# 0.01335f
C3207 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 a_15317_6250# 0.02792f
C3208 a_43698_9766# VDDH 0.23565f
C3209 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04797f
C3210 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.04748f
C3211 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.14454f
C3212 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A a_43724_9926# 0.08029f
C3213 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_15098_19866# 0.18368f
C3214 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y a_45023_21136# 0.01031f
C3215 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.17508f
C3216 a_44234_17252# a_44234_16896# 0.08026f
C3217 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax VOUT 0.0675f
C3218 a_34186_8950# a_30332_7686# 0.11059f
C3219 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] a_18284_18696# 0.06994f
C3220 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_22479_20174# 0.03035f
C3221 a_44234_11312# a_44234_11946# 0.02262f
C3222 a_15342_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.30851f
C3223 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.06102f
C3224 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44062_19517# 0.02575f
C3225 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_14331_6250# 0.1553f
C3226 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.03996f
C3227 a_43698_8776# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.40011f
C3228 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_11081_13005# 0.0208f
C3229 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] VDDH 0.85743f
C3230 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05296f
C3231 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 3.76093f
C3232 VDDH a_15863_13287# 0.15166f
C3233 a_14615_13785# top_DAC_0/top_final_switch_0.VOUT[2] 0.09077f
C3234 a_43698_13726# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.02263f
C3235 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.90337f
C3236 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.22399f
C3237 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 0.07536f
C3238 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.13135f
C3239 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_final_switch_0.VOUT[2] 0.43345f
C3240 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 a_29434_6250# 0.08626f
C3241 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.09148f
C3242 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.17953f
C3243 top_DAC_0/top_rseg_n_dcell_0.VL2 a_21375_20174# 0.01482f
C3244 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_5050_12595# 4.21941f
C3245 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_15593_6250# 0.19959f
C3246 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.01417f
C3247 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.03021f
C3248 a_15905_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 0.03929f
C3249 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.19658f
C3250 a_44234_6996# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.0685f
C3251 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.20454f
C3252 a_15618_18696# top_DAC_0/top_rseg_n_dcell_0.VL3 0.03849f
C3253 VDDH a_11081_14150# 0.49013f
C3254 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_20547_20174# 0.0892f
C3255 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.43879f
C3256 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01451f
C3257 a_17167_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.07166f
C3258 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 0.10167f
C3259 a_16181_7686# a_16615_7686# 6.11601f
C3260 a_15905_7686# a_16891_7686# 0.16296f
C3261 a_15353_7686# a_17443_7686# 0.39018f
C3262 a_15629_7686# a_17167_7686# 0.1611f
C3263 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 0.01986f
C3264 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB a_44234_6996# 0.07929f
C3265 a_36888_19550# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.07596f
C3266 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.11835f
C3267 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 0.06168f
C3268 a_23629_18133# a_21375_20174# 0.01734f
C3269 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.VS1 0.07695f
C3270 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.01383f
C3271 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_final_switch_0.VOUT[2] 0.16603f
C3272 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 a_14331_6250# 0.02784f
C3273 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_12936# 0.02704f
C3274 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.05155f
C3275 top_DAC_0/top_final_switch_0.VOUT[4] a_12809_14150# 0.01964f
C3276 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 a_30608_7686# 0.03955f
C3277 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 0.58085f
C3278 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_30056_7686# 0.08497f
C3279 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.09522f
C3280 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB VDD 0.31603f
C3281 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.04742f
C3282 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN a_5050_12595# 1.39442f
C3283 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.23045f
C3284 VDDH a_12809_15057# 0.48955f
C3285 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.61765f
C3286 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 1.27264f
C3287 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.05972f
C3288 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 1.88678f
C3289 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_13292# 0.03152f
C3290 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 0.16844f
C3291 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 1.45197f
C3292 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.09009f
C3293 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 0.02172f
C3294 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 0.28555f
C3295 VDDH top_DAC_0/top_rseg_n_dcell_0.VH3 0.46642f
C3296 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.08933f
C3297 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 2.09225f
C3298 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.03331f
C3299 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] DIN6 0.01584f
C3300 a_8051_10107# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 0.43083f
C3301 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.17474f
C3302 a_34873_10031# a_35453_10031# 0.17152f
C3303 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.09386f
C3304 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 0.02052f
C3305 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 0.07766f
C3306 a_19552_8950# a_20222_8950# 0.08994f
C3307 a_19670_8950# a_19946_8950# 3.02842f
C3308 VDDH a_6445_14150# 0.49013f
C3309 a_30056_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.07155f
C3310 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44062_18093# 0.01914f
C3311 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_21927_20174# 0.11574f
C3312 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.11409f
C3313 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.73748f
C3314 a_19276_8950# a_20656_10031# 0.0648f
C3315 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 a_13779_6250# 0.04213f
C3316 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01401f
C3317 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_31594_7686# 0.11771f
C3318 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.02784f
C3319 a_8506_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.22623f
C3320 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_14948_18696# 0.18233f
C3321 a_43724_12896# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.08245f
C3322 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 VDDH 0.15179f
C3323 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 a_21651_20174# 0.06393f
C3324 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_final_switch_0.VOUT[3] 0.01843f
C3325 a_17148_18696# a_14790_18696# 0.06536f
C3326 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_9353_15057# 0.04959f
C3327 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.17828f
C3328 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1896_19053# 0.02486f
C3329 a_15353_7686# a_19000_8950# 0.07803f
C3330 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 a_28606_6250# 0.02793f
C3331 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_final_switch_0.VOUT[4] 0.01837f
C3332 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 1.47626f
C3333 VDDH a_16872_18696# 0.29355f
C3334 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 a_29434_6250# 0.2523f
C3335 top_DAC_0/top_final_switch_0.VOUT[0] a_4717_13005# 0.02832f
C3336 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 a_28882_6250# 0.02794f
C3337 a_34304_8950# a_35132_8950# 0.1029f
C3338 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 a_15317_6250# 0.03939f
C3339 a_34580_8950# a_34856_8950# 3.18941f
C3340 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 a_21375_20174# 0.06393f
C3341 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 a_29158_6250# 0.03986f
C3342 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 0.05675f
C3343 VOUT a_9353_13005# 0.02203f
C3344 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.02787f
C3345 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.09267f
C3346 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04929f
C3347 a_1636_15118# a_2300_15118# 0.01589f
C3348 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.04356f
C3349 a_15629_7686# a_14607_6250# 0.04155f
C3350 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 a_27896_6250# 0.03957f
C3351 a_16181_7686# a_14055_6250# 0.02787f
C3352 a_15353_7686# a_15041_6250# 0.05229f
C3353 a_15905_7686# a_14331_6250# 0.0279f
C3354 a_31594_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.02681f
C3355 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 1.85017f
C3356 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 0.05989f
C3357 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.02433f
C3358 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.02218f
C3359 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.02156f
C3360 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD 0.21631f
C3361 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN a_44234_9332# 0.27324f
C3362 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_1896_21703# 0.06357f
C3363 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.09271f
C3364 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.12526f
C3365 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 0.05104f
C3366 a_14790_18696# a_15618_18696# 0.09082f
C3367 a_15066_18696# a_15342_18696# 1.99649f
C3368 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.02015f
C3369 DIN4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.03501f
C3370 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.03939f
C3371 a_35453_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.17274f
C3372 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.04212f
C3373 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 0.01456f
C3374 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 0.35706f
C3375 a_24963_20174# a_21651_20174# 0.13435f
C3376 a_30056_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.12792f
C3377 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.15149f
C3378 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 a_14055_6250# 0.03503f
C3379 top_DAC_0/top_rseg_n_dcell_0.VL2 a_23049_18133# 0.57932f
C3380 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 a_14055_6250# 0.02804f
C3381 a_24963_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.0304f
C3382 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.19936f
C3383 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 0.0205f
C3384 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_29158_6250# 0.46027f
C3385 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 0.87542f
C3386 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_43698_14716# 0.24498f
C3387 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.14057f
C3388 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.12651f
C3389 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_15905_7686# 0.08296f
C3390 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 0.1869f
C3391 VDDH a_19670_8950# 0.26787f
C3392 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 a_22203_20174# 0.07763f
C3393 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.16354f
C3394 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_20823_20174# 0.17206f
C3395 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.02794f
C3396 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.09346f
C3397 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.07179f
C3398 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.18966f
C3399 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_final_switch_0.VOUT[1] 0.05883f
C3400 a_23049_18133# a_23629_18133# 3.42875f
C3401 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.2781f
C3402 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN a_43391_3794# 0.01004f
C3403 VDDH a_1636_15118# 0.554f
C3404 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.25426f
C3405 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.0765f
C3406 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 a_27620_6250# 0.04583f
C3407 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_4978_9535# 0.11619f
C3408 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 0.42912f
C3409 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B a_2678_17510# 0.06357f
C3410 a_43698_9766# a_44234_10322# 0.07082f
C3411 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 4.05461f
C3412 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 0.04501f
C3413 a_30056_7686# a_30608_7686# 0.17062f
C3414 a_29780_7686# a_31042_7686# 0.2076f
C3415 a_28882_6250# a_31870_7686# 0.05986f
C3416 a_29434_6250# a_31318_7686# 0.03865f
C3417 a_29158_6250# a_31594_7686# 0.02797f
C3418 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_11081_14150# 0.04959f
C3419 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 3.40713f
C3420 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.66352f
C3421 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 0.04154f
C3422 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 a_23031_20174# 0.06246f
C3423 a_24963_20174# a_23031_20174# 4.76539f
C3424 a_24687_20174# a_23307_20174# 5.15441f
C3425 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.03788f
C3426 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 0.02715f
C3427 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 0.21461f
C3428 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.04809f
C3429 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 3.9742f
C3430 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.04638f
C3431 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.1433f
C3432 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 0.15493f
C3433 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_20498_8950# 0.18566f
C3434 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.10584f
C3435 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1 0.07424f
C3436 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04891f
C3437 a_31318_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 0.07402f
C3438 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 1.73459f
C3439 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.15587f
C3440 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_7352# 0.0135f
C3441 DIN0 VDD 0.71624f
C3442 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 8.15945f
C3443 a_43698_12736# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.24498f
C3444 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_22203_20174# 0.17392f
C3445 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_15869_6250# 0.30043f
C3446 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.28825f
C3447 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.VL3 0.10185f
C3448 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.0583f
C3449 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.12577f
C3450 a_16891_7686# a_17443_7686# 0.18419f
C3451 a_17148_18696# a_16872_18696# 1.84244f
C3452 a_31594_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.07166f
C3453 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 a_20547_20174# 0.08782f
C3454 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] a_16596_18696# 0.12303f
C3455 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_28606_6250# 0.31084f
C3456 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.03011f
C3457 VDDH a_43724_8936# 0.09227f
C3458 a_31042_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.03947f
C3459 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.05396f
C3460 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD VOUT 0.61932f
C3461 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_6445_14150# 0.04994f
C3462 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 1.24381f
C3463 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.09114f
C3464 a_35757_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05279f
C3465 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 VOUT 0.13144f
C3466 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.22726f
C3467 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB 2.66992f
C3468 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_5111_8388# 1.28797f
C3469 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.07006f
C3470 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 0.02179f
C3471 top_DAC_0/top_rseg_n_dcell_0.VH2 a_14615_14034# 0.14285f
C3472 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 0.02197f
C3473 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09344f
C3474 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.7893f
C3475 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 0.06616f
C3476 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.05223f
C3477 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.02784f
C3478 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_20823_20174# 0.17184f
C3479 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 0.77514f
C3480 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.06292f
C3481 a_5050_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 0.12707f
C3482 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.23991f
C3483 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN a_5642_8388# 0.01976f
C3484 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.09997f
C3485 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 16.6023f
C3486 a_15629_7686# a_19276_8950# 0.08519f
C3487 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.05174f
C3488 a_4717_14150# VOUT 0.05095f
C3489 a_17148_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 0.0686f
C3490 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 0.19125f
C3491 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 2.32429f
C3492 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04798f
C3493 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 a_27620_6250# 0.03677f
C3494 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.21873f
C3495 a_5897_15057# a_6445_15057# 0.0237f
C3496 a_24135_20174# a_24411_20174# 0.47801f
C3497 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 a_27344_6250# 0.03333f
C3498 a_23859_20174# a_24687_20174# 0.15275f
C3499 a_23583_20174# a_24963_20174# 0.12463f
C3500 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.05928f
C3501 a_15629_7686# a_16181_7686# 0.17062f
C3502 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 a_29158_6250# 0.02801f
C3503 top_DAC_0/top_rseg_n_dcell_0.VS1 a_34569_10031# 0.38809f
C3504 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP a_43724_13886# 0.08245f
C3505 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 a_22479_20174# 0.08495f
C3506 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN VOUT 0.44339f
C3507 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.14904f
C3508 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.26447f
C3509 a_14615_14283# top_DAC_0/top_final_switch_0.VOUT[3] 0.05835f
C3510 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.05681f
C3511 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.04269f
C3512 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_18008_18696# 0.13999f
C3513 a_19468_10031# top_DAC_0/top_rseg_n_dcell_0.VS4 0.38967f
C3514 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 16.8926f
C3515 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.1019f
C3516 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 0.07411f
C3517 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 10.3939f
C3518 a_31594_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.05498f
C3519 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_13779_6250# 0.1074f
C3520 a_44234_16896# a_44234_16262# 0.02262f
C3521 DIN1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.17975f
C3522 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_43698_13726# 0.01234f
C3523 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 a_15629_7686# 0.07155f
C3524 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_22203_20174# 0.17684f
C3525 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.55643f
C3526 a_15041_6250# a_16891_7686# 0.05053f
C3527 a_14331_6250# a_17443_7686# 0.06275f
C3528 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 0.04881f
C3529 a_14607_6250# a_17167_7686# 0.04941f
C3530 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.VS4 0.06204f
C3531 a_1896_17510# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.06357f
C3532 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.01806f
C3533 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_24209_18133# 0.0628f
C3534 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 0.07007f
C3535 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.04417f
C3536 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.03135f
C3537 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 1.19314f
C3538 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_27344_6250# 0.74054f
C3539 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 VDDH 0.02285f
C3540 a_43698_12736# a_44234_12936# 0.0139f
C3541 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 1.81049f
C3542 a_43724_17292# a_43698_16696# 0.06762f
C3543 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.14569f
C3544 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_35177_10031# 0.18826f
C3545 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.06201f
C3546 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 10.3151f
C3547 a_38672_20477# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.37724f
C3548 a_43698_16696# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.02263f
C3549 a_28172_6250# a_29434_6250# 0.18915f
C3550 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.02575f
C3551 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.02791f
C3552 a_28606_6250# a_29158_6250# 0.16957f
C3553 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] DIN7 0.17937f
C3554 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 0.03251f
C3555 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.10397f
C3556 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.02726f
C3557 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.04304f
C3558 a_20547_20174# a_21927_20174# 0.24743f
C3559 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.09568f
C3560 a_4717_15057# VOUT 0.0236f
C3561 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 a_14055_6250# 0.07806f
C3562 VDDH a_43724_12342# 0.09227f
C3563 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 0.49734f
C3564 a_2678_11886# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.0175f
C3565 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 0.20729f
C3566 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.09163f
C3567 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.59731f
C3568 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.05765f
C3569 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 16.2949f
C3570 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_17443_7686# 0.08787f
C3571 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43698_13726# 0.06167f
C3572 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.07189f
C3573 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.08402f
C3574 a_31594_7686# a_27344_6250# 0.03764f
C3575 a_31042_7686# a_27896_6250# 0.02794f
C3576 a_31318_7686# a_27620_6250# 0.02791f
C3577 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 a_15869_6250# 0.08609f
C3578 VOUT a_6923_9707# 0.55146f
C3579 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.06132f
C3580 a_36813_19462# a_36888_19550# 0.01119f
C3581 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 0.08495f
C3582 a_37595_19462# a_36888_19786# 0.04324f
C3583 a_20932_10031# a_19000_8950# 0.06493f
C3584 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_15863_13287# 0.03337f
C3585 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_11081_12507# 0.0208f
C3586 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_44062_18805# 0.06327f
C3587 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.0436f
C3588 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] a_15224_18696# 0.03329f
C3589 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_20932_10031# 0.55228f
C3590 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 2.15445f
C3591 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.0206f
C3592 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.04341f
C3593 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.VS4 0.03261f
C3594 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.01388f
C3595 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.02583f
C3596 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.0811f
C3597 a_14331_6250# a_19000_8950# 0.08536f
C3598 a_44234_10956# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.02704f
C3599 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 0.0547f
C3600 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.09785f
C3601 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3 0.05382f
C3602 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04799f
C3603 a_34304_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.04014f
C3604 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 17.3168f
C3605 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.04736f
C3606 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.0152f
C3607 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 0.04827f
C3608 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.1802f
C3609 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.08235f
C3610 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.29969f
C3611 a_15374_19866# a_16872_18696# 0.08835f
C3612 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 a_17167_7686# 0.03977f
C3613 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.07239f
C3614 a_33634_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.06194f
C3615 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.31328f
C3616 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B a_43391_3878# 0.01136f
C3617 a_44234_11312# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.03152f
C3618 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_37410_19098# 1.01772f
C3619 a_14331_6250# a_15041_6250# 0.18706f
C3620 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.0897f
C3621 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.05787f
C3622 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_7352# 0.1344f
C3623 a_15342_18696# VDDH 0.21588f
C3624 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_16615_7686# 0.06495f
C3625 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 0.23023f
C3626 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] a_16320_18696# 0.03156f
C3627 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 a_15041_6250# 0.02791f
C3628 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB a_44234_8342# 0.08623f
C3629 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_19000_8950# 0.06137f
C3630 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.10191f
C3631 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 a_15869_6250# 0.04612f
C3632 a_4978_9535# a_4978_8388# 0.015f
C3633 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.VH3 0.04787f
C3634 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.10923f
C3635 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.09785f
C3636 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.13195f
C3637 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_20222_8950# 0.03763f
C3638 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.03386f
C3639 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.49177f
C3640 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.22369f
C3641 a_44062_20941# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.07788f
C3642 a_43724_11352# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP 0.03147f
C3643 a_44234_11312# a_43698_10756# 0.07082f
C3644 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_15041_6250# 0.16727f
C3645 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 1.57341f
C3646 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.15777f
C3647 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 1.30528f
C3648 a_35132_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.10475f
C3649 a_43724_12896# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.03597f
C3650 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.38958f
C3651 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04068f
C3652 VDDH a_43724_10362# 0.09227f
C3653 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 a_27344_6250# 0.06651f
C3654 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 0.02014f
C3655 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.35096f
C3656 a_43698_8776# a_44234_9332# 0.07082f
C3657 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 0.02017f
C3658 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.11542f
C3659 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 a_31042_7686# 0.07963f
C3660 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.02791f
C3661 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 a_30332_7686# 0.03929f
C3662 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 0.79254f
C3663 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.0975f
C3664 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.30079f
C3665 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_15353_7686# 0.21071f
C3666 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.06014f
C3667 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.03422f
C3668 a_17167_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.03944f
C3669 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 0.05973f
C3670 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.13831f
C3671 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_21099_20174# 0.11555f
C3672 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 a_15317_6250# 0.02791f
C3673 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.08388f
C3674 a_16181_7686# a_17167_7686# 0.16293f
C3675 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 9.22813f
C3676 a_15905_7686# a_17443_7686# 0.17666f
C3677 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.72875f
C3678 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.37639f
C3679 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.07477f
C3680 a_45023_21412# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.01005f
C3681 a_4415_23194# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 1.64212f
C3682 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 2.13381f
C3683 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_20076_10031# 0.02244f
C3684 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 a_15041_6250# 0.02784f
C3685 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.10026f
C3686 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.45254f
C3687 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 0.10863f
C3688 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.08837f
C3689 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 8.34443f
C3690 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_23629_18133# 0.25057f
C3691 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.01812f
C3692 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 a_31594_7686# 0.07166f
C3693 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.74385f
C3694 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 a_31042_7686# 0.03947f
C3695 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.04476f
C3696 VDDH a_12809_14150# 0.48022f
C3697 a_5111_8388# a_4978_8388# 0.03284f
C3698 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_14055_6250# 0.16545f
C3699 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.02452f
C3700 a_15353_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 0.03929f
C3701 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.09358f
C3702 a_28606_6250# a_27344_6250# 0.21112f
C3703 a_28172_6250# a_27620_6250# 0.1621f
C3704 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.02488f
C3705 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD 0.2275f
C3706 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 a_14672_18696# 0.06349f
C3707 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.04899f
C3708 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 0.01391f
C3709 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 0.02053f
C3710 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP a_43698_14716# 0.02263f
C3711 a_43698_13726# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP 0.40164f
C3712 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 0.21897f
C3713 a_34873_10031# a_36033_10031# 0.10606f
C3714 a_35177_10031# a_35757_10031# 0.05093f
C3715 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 15.219f
C3716 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 1.3535f
C3717 a_19670_8950# a_20498_8950# 0.10233f
C3718 a_19946_8950# a_20222_8950# 3.03941f
C3719 a_34873_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.20148f
C3720 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.02791f
C3721 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 1.80576f
C3722 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_22479_20174# 0.11942f
C3723 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.73909f
C3724 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.08566f
C3725 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 1.38112f
C3726 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 a_14331_6250# 0.02788f
C3727 a_19276_8950# a_18724_8950# 0.10175f
C3728 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.08559f
C3729 a_15098_19866# VDDH 0.57537f
C3730 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.02784f
C3731 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_16320_18696# 0.1193f
C3732 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.04818f
C3733 a_35177_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.06133f
C3734 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.04843f
C3735 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 0.07563f
C3736 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1896_17510# 0.06525f
C3737 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 a_29158_6250# 0.02802f
C3738 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 a_30056_7686# 0.07245f
C3739 a_44062_18449# a_44062_18805# 0.04541f
C3740 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.02797f
C3741 a_34856_8950# a_35132_8950# 3.21691f
C3742 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.02121f
C3743 top_DAC_0/top_final_switch_0.VOUT[0] a_5897_13005# 0.03196f
C3744 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 a_29434_6250# 0.04269f
C3745 a_14607_6250# a_19276_8950# 0.07793f
C3746 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.24881f
C3747 VOUT a_9353_12507# 0.04471f
C3748 VDDH top_DAC_0/top_rseg_n_dcell_0.VS4 0.47346f
C3749 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 0.09272f
C3750 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.02789f
C3751 VDDH a_43724_16856# 0.09227f
C3752 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 a_6778_12595# 0.04978f
C3753 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.1701f
C3754 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_9901_15057# 0.04959f
C3755 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 a_27896_6250# 0.03957f
C3756 VDDH a_2678_22970# 0.77537f
C3757 a_16181_7686# a_14607_6250# 0.04309f
C3758 a_15905_7686# a_15041_6250# 0.03872f
C3759 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.04851f
C3760 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_final_switch_0.VOUT[4] 0.03109f
C3761 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 a_1896_20320# 0.03145f
C3762 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.11733f
C3763 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP 0.17254f
C3764 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] a_17732_18696# 0.29618f
C3765 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_2678_11886# 0.02366f
C3766 a_43698_12736# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP 0.40164f
C3767 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_final_switch_0.VOUT[2] 0.05877f
C3768 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.05177f
C3769 a_15342_18696# a_15618_18696# 1.98501f
C3770 a_33910_8950# a_28172_6250# 0.07793f
C3771 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 1.90109f
C3772 a_36033_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.53872f
C3773 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.02787f
C3774 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN VDD 3.53251f
C3775 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.09922f
C3776 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 a_14607_6250# 0.03281f
C3777 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 a_14607_6250# 0.03556f
C3778 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.01149f
C3779 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_29780_7686# 0.54354f
C3780 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.05224f
C3781 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 0.05483f
C3782 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_36888_19550# 0.18067f
C3783 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.06145f
C3784 VDDH a_20222_8950# 0.3357f
C3785 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.02784f
C3786 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA VOUT 26.2719f
C3787 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.56882f
C3788 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.09032f
C3789 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_21375_20174# 0.17641f
C3790 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 3.83598f
C3791 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 0.32979f
C3792 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.06127f
C3793 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.11409f
C3794 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 1.3734f
C3795 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 0.02715f
C3796 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.02821f
C3797 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.05318f
C3798 a_44234_16262# a_44234_15906# 0.08026f
C3799 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.VL3 0.06414f
C3800 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 0.01926f
C3801 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.168f
C3802 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 3.95069f
C3803 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 a_16615_7686# 0.07989f
C3804 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.17101f
C3805 a_19468_10031# a_19772_10031# 0.71479f
C3806 VDDH a_1636_14353# 0.53376f
C3807 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.32704f
C3808 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 2.01261f
C3809 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.0596f
C3810 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.04858f
C3811 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.46395f
C3812 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 1.44458f
C3813 a_43698_9766# a_43724_9926# 0.02395f
C3814 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.05806f
C3815 a_29780_7686# a_31594_7686# 0.21699f
C3816 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.04173f
C3817 a_30056_7686# a_31318_7686# 0.16163f
C3818 a_29434_6250# a_31870_7686# 0.05681f
C3819 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 0.01992f
C3820 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 a_28172_6250# 0.02787f
C3821 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.59336f
C3822 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.03957f
C3823 VDDH a_43724_14322# 0.09227f
C3824 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_9332# 0.01697f
C3825 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_9353_13005# 0.0208f
C3826 a_30608_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.07998f
C3827 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 a_28606_6250# 0.08399f
C3828 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 0.9868f
C3829 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 a_14055_6250# 0.05228f
C3830 a_44062_22009# VDDH 0.04324f
C3831 a_43698_9766# a_43698_8776# 0.01563f
C3832 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.03939f
C3833 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD VOUT 0.61926f
C3834 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.05186f
C3835 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_39883_19854# 0.02806f
C3836 VOUT a_8173_15057# 0.01454f
C3837 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 0.04533f
C3838 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.09162f
C3839 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 0.1877f
C3840 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.01887f
C3841 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_16891_7686# 0.111f
C3842 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.SH[2] 19.0673f
C3843 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_15629_7686# 0.06774f
C3844 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 1.24591f
C3845 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.96691f
C3846 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_12809_14150# 0.04134f
C3847 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.05359f
C3848 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_22755_20174# 0.20842f
C3849 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 0.22947f
C3850 a_15098_19866# a_17148_18696# 0.1863f
C3851 a_24135_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 0.06449f
C3852 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.03966f
C3853 a_35453_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.2139f
C3854 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.02197f
C3855 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.05322f
C3856 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C3857 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.09553f
C3858 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.06147f
C3859 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.0543f
C3860 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_29158_6250# 0.22365f
C3861 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.60184f
C3862 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_18724_8950# 0.8009f
C3863 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_final_switch_0.VOUT[1] 0.01299f
C3864 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.01148f
C3865 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.01349f
C3866 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 0.91003f
C3867 a_33358_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.07757f
C3868 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 0.54952f
C3869 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.08493f
C3870 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 a_14615_13536# 0.08047f
C3871 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 1.89956f
C3872 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 a_15905_7686# 0.07404f
C3873 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.11433f
C3874 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 0.1216f
C3875 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.09623f
C3876 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 0.69946f
C3877 top_DAC_0/top_rseg_n_dcell_0.VH2 a_14615_13536# 0.09891f
C3878 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.02784f
C3879 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_21375_20174# 0.181f
C3880 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_final_switch_0.VOUT[3] 0.05518f
C3881 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04995f
C3882 a_15098_19866# a_15618_18696# 0.05271f
C3883 a_15374_19866# a_15342_18696# 0.04105f
C3884 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_9372# 0.03597f
C3885 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.02791f
C3886 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.50988f
C3887 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 a_14055_6250# 0.02788f
C3888 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.14625f
C3889 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 0.01797f
C3890 a_39861_22496# VDDH 1.43189f
C3891 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_19772_10031# 0.28703f
C3892 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 2.25141f
C3893 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.84185f
C3894 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1896_20320# 0.07342f
C3895 a_23859_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 0.06438f
C3896 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 a_27344_6250# 0.0453f
C3897 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.60657f
C3898 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.11881f
C3899 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.31465f
C3900 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.02715f
C3901 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 1.3157f
C3902 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 a_27620_6250# 0.02791f
C3903 a_24411_20174# a_24687_20174# 0.69559f
C3904 a_24135_20174# a_24963_20174# 0.43501f
C3905 a_14790_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.1541f
C3906 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.05182f
C3907 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.20837f
C3908 a_20547_20174# a_21099_20174# 0.15164f
C3909 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.05175f
C3910 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.02186f
C3911 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.096f
C3912 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.VL3 0.18968f
C3913 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.66863f
C3914 a_33910_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.02742f
C3915 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.48886f
C3916 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.32927f
C3917 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 0.0209f
C3918 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.0719f
C3919 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_final_switch_0.VOUT[3] 0.43345f
C3920 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 a_22203_20174# 0.04147f
C3921 a_15905_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.07456f
C3922 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_14331_6250# 0.15913f
C3923 a_43724_15866# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.08245f
C3924 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP 0.92839f
C3925 a_43698_15706# a_44234_16262# 0.07082f
C3926 a_44234_6996# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.0862f
C3927 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.01388f
C3928 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.33918f
C3929 VDDH a_43724_8382# 0.09227f
C3930 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.28496f
C3931 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.04842f
C3932 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04948f
C3933 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_22755_20174# 0.23063f
C3934 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 a_16181_7686# 0.08f
C3935 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.05782f
C3936 a_14615_14283# top_DAC_0/top_final_switch_0.VOUT[4] 0.11595f
C3937 a_15041_6250# a_17443_7686# 0.24181f
C3938 a_6778_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.11462f
C3939 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04071f
C3940 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.98866f
C3941 a_5050_12595# a_8051_10107# 0.01462f
C3942 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 0.07044f
C3943 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_27896_6250# 0.15577f
C3944 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_final_switch_0.VOUT[3] 0.04992f
C3945 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 3.75653f
C3946 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.11409f
C3947 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.59845f
C3948 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_35757_10031# 0.10876f
C3949 a_44234_16896# a_43698_16696# 0.0139f
C3950 a_38584_20389# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.02882f
C3951 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.08462f
C3952 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.08304f
C3953 a_28882_6250# a_29434_6250# 0.1847f
C3954 a_28172_6250# a_30056_7686# 0.0412f
C3955 a_28606_6250# a_29780_7686# 0.053f
C3956 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 0.0199f
C3957 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.20768f
C3958 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.15363f
C3959 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.02786f
C3960 a_20823_20174# a_22203_20174# 4.95211f
C3961 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 16.2094f
C3962 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 a_23307_20174# 0.06406f
C3963 a_21099_20174# a_21927_20174# 5.3f
C3964 a_20547_20174# a_22479_20174# 4.6659f
C3965 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_12936# 0.03855f
C3966 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 0.04802f
C3967 a_43724_12342# a_43698_11746# 0.06762f
C3968 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 0.01789f
C3969 a_11629_13005# top_DAC_0/top_final_switch_0.VOUT[4] 0.02842f
C3970 top_DAC_0/top_final_switch_0.VOUT[0] a_6445_15057# 0.01175f
C3971 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.13636f
C3972 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.08118f
C3973 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.2193f
C3974 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 0.01782f
C3975 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 0.01681f
C3976 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3 0.23498f
C3977 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.11409f
C3978 a_44255_4162# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.01264f
C3979 a_44234_9332# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.08449f
C3980 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.09515f
C3981 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09325f
C3982 a_19552_8950# a_20352_10031# 0.06482f
C3983 a_19670_8950# a_20076_10031# 0.05067f
C3984 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 4.14638f
C3985 a_31594_7686# a_27896_6250# 0.02801f
C3986 a_31870_7686# a_27620_6250# 0.04962f
C3987 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 0.03927f
C3988 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05675f
C3989 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 1.26896f
C3990 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.09644f
C3991 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 1.45085f
C3992 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.14572f
C3993 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_6923_9707# 0.5135f
C3994 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.05594f
C3995 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.14576f
C3996 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] VDDH 2.61713f
C3997 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 a_20823_20174# 0.06397f
C3998 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09746f
C3999 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_19000_8950# 0.02591f
C4000 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.VH3 0.05157f
C4001 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.04499f
C4002 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.60845f
C4003 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_11081_15057# 0.04959f
C4004 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.09146f
C4005 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.02784f
C4006 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 0.05594f
C4007 a_15098_19866# a_15374_19866# 1.77428f
C4008 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.08425f
C4009 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.0119f
C4010 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.02953f
C4011 a_34856_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.06049f
C4012 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.11672f
C4013 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 2.25734f
C4014 a_21927_20174# a_22479_20174# 0.29179f
C4015 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.21507f
C4016 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.03135f
C4017 a_44234_6996# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.07056f
C4018 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.06525f
C4019 a_34186_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.04904f
C4020 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 0.04511f
C4021 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.08314f
C4022 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.01253f
C4023 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 a_21927_20174# 0.07411f
C4024 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_27344_6250# 0.15553f
C4025 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.36625f
C4026 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 1.72824f
C4027 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_19276_8950# 0.12809f
C4028 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 0.01392f
C4029 DIN0 VDDH 0.4291f
C4030 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.49342f
C4031 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_17167_7686# 0.06372f
C4032 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_16615_7686# 0.03056f
C4033 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 0.05599f
C4034 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] a_16872_18696# 0.03108f
C4035 a_34873_10031# top_DAC_0/top_rseg_n_dcell_0.VS1 0.06091f
C4036 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44062_18805# 0.0242f
C4037 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.05772f
C4038 a_9353_15057# a_9901_15057# 0.0237f
C4039 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_34569_10031# 0.22523f
C4040 VDDH a_1896_22970# 0.74102f
C4041 a_43698_7786# VDDH 0.23565f
C4042 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.09276f
C4043 DIN0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.03542f
C4044 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.77374f
C4045 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.02611f
C4046 a_34304_8950# a_31318_7686# 0.1105f
C4047 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.7544f
C4048 VDDH a_5111_10963# 0.01434f
C4049 a_43724_10916# a_43698_10756# 0.02395f
C4050 a_44234_10956# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP 0.06668f
C4051 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.11733f
C4052 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_1896_12504# 0.02948f
C4053 VDDH a_19772_10031# 0.19531f
C4054 a_44234_12302# a_44234_11946# 0.08026f
C4055 a_24209_18133# a_20823_20174# 0.04174f
C4056 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_36888_19786# 0.02243f
C4057 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB VDD 0.6501f
C4058 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_6923_9707# 0.556f
C4059 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 0.15598f
C4060 a_43724_10916# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.03597f
C4061 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 a_27896_6250# 0.02788f
C4062 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B VDD 0.4727f
C4063 a_43698_8776# a_43724_8936# 0.02395f
C4064 VDDH a_43698_16696# 0.24624f
C4065 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.13028f
C4066 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.VS1 0.05653f
C4067 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.04506f
C4068 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.12875f
C4069 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 1.36438f
C4070 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 1.39235f
C4071 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_15905_7686# 0.11618f
C4072 DIN2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.03543f
C4073 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] VDD 0.48049f
C4074 VOUT a_9353_15057# 0.04641f
C4075 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 0.12042f
C4076 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_21651_20174# 0.11563f
C4077 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 a_15869_6250# 0.04262f
C4078 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.VS4 0.03256f
C4079 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.12207f
C4080 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 1.72334f
C4081 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 0.01015f
C4082 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 0.04875f
C4083 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.16544f
C4084 VDDH top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 2.1824f
C4085 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_33634_8950# 0.11409f
C4086 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C4087 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.VS1 0.07752f
C4088 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_44062_20941# 0.02123f
C4089 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.1268f
C4090 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.6765f
C4091 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 0.3799f
C4092 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 12.9813f
C4093 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 1.34502f
C4094 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.77287f
C4095 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 0.0315f
C4096 a_5642_9535# a_5642_8388# 0.015f
C4097 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.VH3 0.16414f
C4098 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 3.81788f
C4099 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_14607_6250# 0.27888f
C4100 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04936f
C4101 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_37410_19098# 0.13149f
C4102 a_17148_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.88189f
C4103 a_28606_6250# a_27896_6250# 0.1869f
C4104 a_29158_6250# a_27344_6250# 0.18965f
C4105 a_28882_6250# a_27620_6250# 0.15375f
C4106 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.06891f
C4107 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.20766f
C4108 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.09612f
C4109 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 a_28882_6250# 0.08549f
C4110 a_9901_13005# top_DAC_0/top_final_switch_0.VOUT[3] 0.02844f
C4111 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 a_28172_6250# 0.03925f
C4112 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.15269f
C4113 a_35453_10031# a_36033_10031# 0.05831f
C4114 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_6778_12595# 0.17535f
C4115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_17252# 0.02754f
C4116 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 0.78654f
C4117 a_20222_8950# a_20498_8950# 3.06634f
C4118 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.09972f
C4119 a_8051_10107# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 0.26604f
C4120 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.04262f
C4121 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] a_23031_20174# 0.12908f
C4122 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.04724f
C4123 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.82663f
C4124 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 a_15041_6250# 0.02791f
C4125 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 0.0119f
C4126 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.14088f
C4127 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_12936# 0.14379f
C4128 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 0.05518f
C4129 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.34747f
C4130 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_16872_18696# 0.11851f
C4131 a_35132_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.09842f
C4132 a_15317_6250# a_20222_8950# 0.08494f
C4133 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.09759f
C4134 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.01782f
C4135 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 0.04888f
C4136 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 1.57333f
C4137 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 1.94305f
C4138 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 0.02288f
C4139 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.02785f
C4140 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.15977f
C4141 top_DAC_0/top_final_switch_0.VOUT[0] a_5897_12507# 0.01061f
C4142 VOUT a_8051_10107# 0.46019f
C4143 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.15687f
C4144 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN VDD 0.26425f
C4145 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 a_17167_7686# 0.07165f
C4146 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.55369f
C4147 a_1636_14353# a_2300_14353# 0.01589f
C4148 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_9353_12507# 0.0208f
C4149 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.45991f
C4150 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.19185f
C4151 VDDH a_2678_21703# 0.75803f
C4152 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB VDD 0.51982f
C4153 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.09351f
C4154 a_15863_13536# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.02289f
C4155 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 0.65201f
C4156 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 0.01659f
C4157 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.17741f
C4158 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44471_4828# 0.01759f
C4159 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] a_18284_18696# 0.11261f
C4160 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.09997f
C4161 VDDH a_39936_22083# 0.47028f
C4162 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 0.34153f
C4163 top_DAC_0/top_rseg_n_dcell_0.VL2 VDDH 0.14809f
C4164 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 2.80645f
C4165 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_17292# 0.03597f
C4166 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 a_15593_6250# 0.05161f
C4167 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.72924f
C4168 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 a_30332_7686# 0.03985f
C4169 VOUT top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.20902f
C4170 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.02791f
C4171 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 3.10831f
C4172 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.30191f
C4173 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_11629_15057# 0.04959f
C4174 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 0.02043f
C4175 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.062f
C4176 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.10324f
C4177 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.11409f
C4178 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.11044f
C4179 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 0.05595f
C4180 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD 0.23151f
C4181 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04805f
C4182 a_44062_22009# a_44062_21653# 0.04238f
C4183 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.02906f
C4184 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] a_14948_18696# 0.04368f
C4185 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 2.75917f
C4186 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 0.72136f
C4187 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.01851f
C4188 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.11135f
C4189 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.02121f
C4190 a_39861_22496# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 0.07143f
C4191 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_final_switch_0.VOUT[3] 5.48581f
C4192 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.02784f
C4193 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.33486f
C4194 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 0.01317f
C4195 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 1.19654f
C4196 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_final_switch_0.VOUT[1] 0.59493f
C4197 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 0.90644f
C4198 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.0591f
C4199 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.20524f
C4200 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 0.0119f
C4201 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 1.15198f
C4202 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.13166f
C4203 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.2354f
C4204 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.03534f
C4205 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.63434f
C4206 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.10571f
C4207 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_30332_7686# 0.08161f
C4208 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.VS1 0.0717f
C4209 VDDH a_15593_6250# 0.64304f
C4210 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 0.1743f
C4211 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 1.72759f
C4212 a_19468_10031# a_20352_10031# 0.38399f
C4213 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.08675f
C4214 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.16815f
C4215 a_22479_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 0.04143f
C4216 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD a_11629_15057# 0.01033f
C4217 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 0.07287f
C4218 a_22479_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 0.04146f
C4219 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 0.22158f
C4220 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.04843f
C4221 a_30056_7686# a_31870_7686# 0.18599f
C4222 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 0.63647f
C4223 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 a_28882_6250# 0.02787f
C4224 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.07963f
C4225 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.01487f
C4226 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.05244f
C4227 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 a_28172_6250# 0.04346f
C4228 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 a_29158_6250# 0.04481f
C4229 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.06042f
C4230 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 a_28882_6250# 0.03927f
C4231 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 a_14607_6250# 0.04391f
C4232 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 a_28606_6250# 0.02784f
C4233 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.70581f
C4234 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.02079f
C4235 a_44234_10322# a_44234_9966# 0.08026f
C4236 top_DAC_0/top_final_switch_0.VOUT[1] a_8173_15057# 0.01175f
C4237 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 a_27620_6250# 0.03971f
C4238 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_8976# 0.01484f
C4239 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.03934f
C4240 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_17443_7686# 0.14524f
C4241 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 a_16181_7686# 0.06587f
C4242 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_15629_7686# 0.05504f
C4243 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.03934f
C4244 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 VOUT 0.03859f
C4245 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] a_23307_20174# 0.18263f
C4246 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 1.77186f
C4247 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.05535f
C4248 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.11369f
C4249 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB a_44471_4828# 0.02698f
C4250 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.06502f
C4251 a_35757_10031# a_33634_8950# 0.03997f
C4252 a_35453_10031# a_33910_8950# 0.03999f
C4253 a_35177_10031# a_34186_8950# 0.04005f
C4254 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05322f
C4255 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C4256 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 a_21375_20174# 0.06393f
C4257 a_36033_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.24408f
C4258 a_14514_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.108f
C4259 a_44234_10956# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.03855f
C4260 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 0.01623f
C4261 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 1.82582f
C4262 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_29780_7686# 0.17996f
C4263 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.09824f
C4264 a_15224_18696# a_14672_18696# 0.16068f
C4265 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 a_37022_20295# 0.02962f
C4266 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 0.05245f
C4267 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.10545f
C4268 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.07731f
C4269 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.26076f
C4270 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 0.05305f
C4271 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.02197f
C4272 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.08427f
C4273 VOUT a_11629_12507# 0.03463f
C4274 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 1.05534f
C4275 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_28606_6250# 0.05171f
C4276 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 0.8119f
C4277 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 3.48836f
C4278 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.14365f
C4279 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.18308f
C4280 a_16181_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 0.03929f
C4281 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.14076f
C4282 a_33634_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.16804f
C4283 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.06283f
C4284 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.09195f
C4285 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.10794f
C4286 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04969f
C4287 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 0.09809f
C4288 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 1.34945f
C4289 a_44234_10956# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.09046f
C4290 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.3192f
C4291 a_15863_13287# top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.03347f
C4292 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.04091f
C4293 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.02796f
C4294 VDDH a_2678_20320# 0.73328f
C4295 VDDH a_5897_15057# 0.49886f
C4296 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 a_14607_6250# 0.02789f
C4297 a_29780_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.43936f
C4298 a_5050_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 0.07275f
C4299 a_44067_22496# VDDH 1.22217f
C4300 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_20352_10031# 0.08792f
C4301 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.03532f
C4302 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.05224f
C4303 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.06751f
C4304 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.18545f
C4305 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 a_27896_6250# 0.0279f
C4306 a_43698_7786# a_43698_6796# 0.01563f
C4307 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_30332_7686# 0.12057f
C4308 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.06861f
C4309 a_24687_20174# a_24963_20174# 0.89725f
C4310 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.04859f
C4311 a_15342_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.28595f
C4312 top_DAC_0/top_rseg_n_dcell_0.SH[4] top_DAC_0/top_final_switch_0.VOUT[4] 0.05516f
C4313 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 a_23031_20174# 0.06242f
C4314 a_20547_20174# a_21651_20174# 0.33891f
C4315 a_20823_20174# a_21375_20174# 0.34196f
C4316 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.07383f
C4317 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 a_28172_6250# 0.02789f
C4318 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.02572f
C4319 a_16615_7686# a_19670_8950# 0.03954f
C4320 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.02167f
C4321 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.07603f
C4322 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 0.05127f
C4323 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.05188f
C4324 a_23859_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 1.08214f
C4325 top_DAC_0/top_rseg_n_dcell_0.SH[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.06278f
C4326 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.43454f
C4327 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.09544f
C4328 VOUT a_5050_12595# 0.52986f
C4329 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP a_43698_11746# 0.7858f
C4330 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_15041_6250# 0.32998f
C4331 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.08366f
C4332 a_16891_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.03948f
C4333 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_22970# 0.03145f
C4334 a_37022_20713# a_36888_19550# 0.014f
C4335 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04841f
C4336 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 0.05934f
C4337 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 a_14055_6250# 0.02804f
C4338 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_23307_20174# 0.15473f
C4339 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04789f
C4340 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.0673f
C4341 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.0119f
C4342 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 1.21733f
C4343 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 1.31557f
C4344 a_30332_7686# a_30608_7686# 6.3868f
C4345 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_final_switch_0.VOUT[2] 0.04711f
C4346 a_16181_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.03955f
C4347 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_final_switch_0.VOUT[4] 0.44592f
C4348 VDDH a_14615_14283# 0.05318f
C4349 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.5556f
C4350 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.01895f
C4351 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.26572f
C4352 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_33358_8950# 0.20435f
C4353 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02795f
C4354 a_31318_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.07419f
C4355 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 VDDH 0.01148f
C4356 a_43724_16856# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.08245f
C4357 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 a_15593_6250# 0.0394f
C4358 a_43698_15706# a_43698_16696# 0.01563f
C4359 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 a_14672_18696# 0.06226f
C4360 a_30608_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.03955f
C4361 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.23571f
C4362 a_29158_6250# a_29780_7686# 0.0424f
C4363 a_28882_6250# a_30056_7686# 0.028f
C4364 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.25631f
C4365 top_DAC_0/top_final_switch_0.VOUT[1] a_14615_13536# 0.07695f
C4366 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP 0.10923f
C4367 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.04462f
C4368 a_21375_20174# a_22203_20174# 0.34481f
C4369 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 0.02198f
C4370 a_21651_20174# a_21927_20174# 0.96383f
C4371 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 0.04732f
C4372 a_20823_20174# a_22755_20174# 0.17834f
C4373 a_20547_20174# a_23031_20174# 0.13399f
C4374 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 a_36888_19786# 0.5632f
C4375 a_21099_20174# a_22479_20174# 0.14104f
C4376 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN VDD 0.43723f
C4377 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN VDDH 0.01041f
C4378 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.09111f
C4379 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.02787f
C4380 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 1.79741f
C4381 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.05244f
C4382 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.07978f
C4383 a_12809_13005# top_DAC_0/top_final_switch_0.VOUT[4] 0.03376f
C4384 a_8506_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.31066f
C4385 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 3.79808f
C4386 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 1.33963f
C4387 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB a_44234_7352# 0.06676f
C4388 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.42222f
C4389 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.48656f
C4390 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.28615f
C4391 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.85005f
C4392 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.21451f
C4393 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.02715f
C4394 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 1.34745f
C4395 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.10309f
C4396 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_19772_10031# 0.23594f
C4397 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.92839f
C4398 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 a_22755_20174# 0.1103f
C4399 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.03961f
C4400 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.10172f
C4401 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A VOUT 0.95598f
C4402 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.02804f
C4403 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 a_27620_6250# 0.07812f
C4404 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 a_27344_6250# 0.13158f
C4405 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.22753f
C4406 DIN3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.01594f
C4407 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.09197f
C4408 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.08449f
C4409 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.01339f
C4410 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 1.2633f
C4411 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.05183f
C4412 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.06072f
C4413 a_43698_6796# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.78464f
C4414 a_18008_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.31744f
C4415 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 0.1099f
C4416 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.12526f
C4417 a_29780_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.01073f
C4418 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.02785f
C4419 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.04219f
C4420 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04706f
C4421 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.69962f
C4422 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_16262# 0.02704f
C4423 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.02791f
C4424 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP 0.01045f
C4425 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 0.23077f
C4426 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 0.04464f
C4427 a_23859_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.38397f
C4428 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 0.03662f
C4429 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.09f
C4430 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.16165f
C4431 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 4.13148f
C4432 a_21927_20174# a_23031_20174# 0.1325f
C4433 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB a_44234_13926# 0.08412f
C4434 a_22203_20174# a_22755_20174# 0.29618f
C4435 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04841f
C4436 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 0.05026f
C4437 a_15863_13536# top_DAC_0/top_final_switch_0.VOUT[2] 0.01137f
C4438 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15342_18696# 0.14199f
C4439 a_34580_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.04783f
C4440 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.08193f
C4441 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.2543f
C4442 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.08198f
C4443 a_44234_12302# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.03152f
C4444 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.04333f
C4445 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_27896_6250# 0.13293f
C4446 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN DIN5 0.03498f
C4447 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 0.05056f
C4448 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_12809_15057# 0.04134f
C4449 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_2678_17510# 0.0506f
C4450 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 0.21425f
C4451 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 0.01566f
C4452 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 0.02715f
C4453 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_19552_8950# 0.05781f
C4454 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_17167_7686# 0.05317f
C4455 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.09239f
C4456 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 0.09915f
C4457 a_23583_20174# a_20547_20174# 0.13315f
C4458 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_final_switch_0.VOUT[3] 0.19149f
C4459 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y a_45023_19712# 0.01032f
C4460 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 a_13779_6250# 0.04992f
C4461 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.02187f
C4462 VDDH a_43724_15866# 0.09227f
C4463 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.02784f
C4464 top_DAC_0/top_final_switch_0.VOUT[2] a_9901_14150# 0.01204f
C4465 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.1866f
C4466 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.01579f
C4467 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 0.20563f
C4468 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.01776f
C4469 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.11467f
C4470 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.89809f
C4471 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 1.22792f
C4472 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.0119f
C4473 a_44234_10956# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.14379f
C4474 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_2678_10356# 0.04179f
C4475 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.16077f
C4476 a_34580_8950# a_31594_7686# 0.08495f
C4477 a_43698_9766# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP 0.40164f
C4478 a_1896_21703# a_2678_21703# 0.02127f
C4479 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_1896_11886# 0.02948f
C4480 a_24209_18133# a_21375_20174# 0.03339f
C4481 VDDH a_20352_10031# 0.24882f
C4482 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.02163f
C4483 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.11848f
C4484 a_29780_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04787f
C4485 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD a_12809_15057# 0.01033f
C4486 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.17399f
C4487 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.4603f
C4488 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.31985f
C4489 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.1736f
C4490 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_16302# 0.03597f
C4491 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.42152f
C4492 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 0.21361f
C4493 VDDH a_13779_6250# 1.27304f
C4494 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.02775f
C4495 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.0672f
C4496 a_11081_13005# a_11629_13005# 0.0103f
C4497 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.12627f
C4498 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.19158f
C4499 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.VL2 0.54413f
C4500 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 0.06329f
C4501 top_DAC_0/top_rseg_n_dcell_0.VH2 a_22469_18133# 0.54031f
C4502 VDDH a_43724_15312# 0.09227f
C4503 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.04931f
C4504 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09511f
C4505 VOUT a_9353_14150# 0.06741f
C4506 a_23583_20174# a_21927_20174# 0.1323f
C4507 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.09478f
C4508 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.02789f
C4509 a_23049_18133# a_22203_20174# 0.06813f
C4510 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.20891f
C4511 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.12773f
C4512 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.20093f
C4513 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 0.06103f
C4514 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 0.05597f
C4515 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.3906f
C4516 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.04782f
C4517 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_34186_8950# 0.11449f
C4518 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_18724_8950# 0.10738f
C4519 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 2.46853f
C4520 a_22193_18133# a_23629_18133# 0.2151f
C4521 VOUT a_9901_15057# 0.01454f
C4522 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_9332# 0.02478f
C4523 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 3.66239f
C4524 a_43698_7786# a_44234_8342# 0.07082f
C4525 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A a_43724_8382# 0.03253f
C4526 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.04975f
C4527 a_24209_18133# a_22755_20174# 0.04127f
C4528 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.SH[4] 16.3155f
C4529 VOUT top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 0.02759f
C4530 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] a_44062_19873# 0.02123f
C4531 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.03137f
C4532 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 0.69939f
C4533 a_29434_6250# a_27620_6250# 0.17869f
C4534 a_29158_6250# a_27896_6250# 0.15373f
C4535 a_29780_7686# a_27344_6250# 0.05175f
C4536 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y a_44062_18805# 0.1286f
C4537 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.09357f
C4538 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.07524f
C4539 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 0.55841f
C4540 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 0.0686f
C4541 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 a_29434_6250# 0.22058f
C4542 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB a_44255_4614# 0.01152f
C4543 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y VDD 0.28031f
C4544 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_34569_10031# 0.26566f
C4545 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 0.02541f
C4546 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 1.03205f
C4547 a_15863_13785# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04207f
C4548 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.0119f
C4549 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.06218f
C4550 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.07891f
C4551 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.10038f
C4552 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 1.18866f
C4553 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.05413f
C4554 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.63053f
C4555 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1 0.0508f
C4556 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.80349f
C4557 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.01812f
C4558 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 15.8859f
C4559 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_final_switch_0.VOUT[0] 0.07853f
C4560 a_15905_7686# a_19552_8950# 0.11059f
C4561 a_15593_6250# a_20498_8950# 0.11034f
C4562 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_16896# 0.03152f
C4563 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.08134f
C4564 a_33358_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.10624f
C4565 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.05086f
C4566 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB a_44234_12936# 0.09046f
C4567 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.4572f
C4568 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.6007f
C4569 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 0.01616f
C4570 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.10297f
C4571 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.20013f
C4572 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.VS4 0.20368f
C4573 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.02015f
C4574 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 0.0853f
C4575 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.04469f
C4576 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 0.74155f
C4577 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD 0.2275f
C4578 a_15317_6250# a_15593_6250# 7.08969f
C4579 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 0.04477f
C4580 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.04219f
C4581 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_45343_4828# 0.01719f
C4582 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.12989f
C4583 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_8051_10107# 0.51626f
C4584 DIN1 DIN2 0.33f
C4585 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.1322f
C4586 a_44062_21653# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.06327f
C4587 a_34873_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.23085f
C4588 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 a_6778_12595# 0.1876f
C4589 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 a_14331_6250# 0.0852f
C4590 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.01848f
C4591 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.04904f
C4592 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.09809f
C4593 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 0.05463f
C4594 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 0.02015f
C4595 a_1636_13352# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.02725f
C4596 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 a_29158_6250# 0.03991f
C4597 VDDH a_39861_21457# 0.40618f
C4598 a_23049_18133# a_24209_18133# 0.20157f
C4599 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.VS1 0.07707f
C4600 a_33634_8950# a_29780_7686# 0.07803f
C4601 a_34580_8950# a_28606_6250# 0.07768f
C4602 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 0.16418f
C4603 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 0.04751f
C4604 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 a_15353_7686# 0.04539f
C4605 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.01718f
C4606 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.17264f
C4607 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.05182f
C4608 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.12781f
C4609 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 a_31318_7686# 0.07419f
C4610 a_44234_14282# a_44234_13926# 0.08026f
C4611 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.04942f
C4612 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.13343f
C4613 a_44062_22009# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.02354f
C4614 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_14615_13785# 0.02052f
C4615 a_33358_8950# a_27344_6250# 0.03917f
C4616 a_44062_21653# a_44062_21297# 0.04541f
C4617 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 2.1375f
C4618 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.12116f
C4619 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 0.05249f
C4620 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 2.21718f
C4621 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 0.02109f
C4622 a_24135_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.21924f
C4623 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.22059f
C4624 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.09211f
C4625 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 0.13043f
C4626 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.42728f
C4627 a_43698_7786# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.78464f
C4628 a_1896_22970# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 0.09901f
C4629 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.02748f
C4630 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.04856f
C4631 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_31042_7686# 0.07874f
C4632 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.14505f
C4633 VDDH a_15353_7686# 1.12574f
C4634 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.10009f
C4635 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09787f
C4636 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 10.1432f
C4637 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.05695f
C4638 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 1.27692f
C4639 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.02715f
C4640 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.2143f
C4641 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.39965f
C4642 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 4.44061f
C4643 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] a_45343_3894# 0.01081f
C4644 a_4978_11461# a_4978_10963# 0.015f
C4645 a_5111_10963# a_5642_11461# 0.02841f
C4646 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.02179f
C4647 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 1.57551f
C4648 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.02213f
C4649 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.05174f
C4650 top_DAC_0/top_final_switch_0.VOUT[2] top_DAC_0/top_final_switch_0.VOUT[4] 0.11637f
C4651 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.44932f
C4652 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04363f
C4653 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.09249f
C4654 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_44062_19517# 0.02123f
C4655 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 a_29434_6250# 0.04093f
C4656 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 a_28882_6250# 0.04017f
C4657 a_36813_19462# a_36813_19760# 0.015f
C4658 a_19772_10031# a_20076_10031# 0.26136f
C4659 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 0.32257f
C4660 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.01474f
C4661 a_17732_18696# a_18284_18696# 0.76201f
C4662 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 ROUT2 0.0484f
C4663 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_8051_10107# 0.55664f
C4664 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.11368f
C4665 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN VDD 0.77805f
C4666 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.09624f
C4667 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 a_29158_6250# 0.02785f
C4668 a_43698_7786# a_43698_8776# 0.01563f
C4669 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.22756f
C4670 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN a_44234_7986# 0.06681f
C4671 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD a_9901_15057# 0.01035f
C4672 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 0.09433f
C4673 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 0.08058f
C4674 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_19276_8950# 0.1589f
C4675 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 0.05022f
C4676 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04806f
C4677 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 0.06502f
C4678 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 a_16320_18696# 0.06351f
C4679 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 a_27620_6250# 0.03971f
C4680 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y a_44062_21653# 0.1286f
C4681 a_15863_13536# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.03462f
C4682 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.02834f
C4683 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 1.93547f
C4684 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 2.29207f
C4685 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.01222f
C4686 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 9.33133f
C4687 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] VDDH 0.18887f
C4688 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_16181_7686# 0.03035f
C4689 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.43094f
C4690 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 2.89925f
C4691 a_43698_16696# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.7858f
C4692 a_33358_8950# a_33634_8950# 2.85416f
C4693 a_27344_6250# a_27896_6250# 0.19547f
C4694 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.09024f
C4695 VDDH a_43724_7392# 0.09227f
C4696 a_15066_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.17423f
C4697 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 1.15343f
C4698 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 0.18469f
C4699 a_14948_18696# a_16320_18696# 0.09026f
C4700 a_15224_18696# a_16596_18696# 0.08858f
C4701 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 1.97838f
C4702 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_9332# 0.1344f
C4703 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 15.2414f
C4704 a_43698_9766# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.02387f
C4705 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 0.51079f
C4706 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD VOUT 0.62599f
C4707 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_29158_6250# 0.06546f
C4708 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.09811f
C4709 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 1.73519f
C4710 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.01687f
C4711 a_34186_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.32242f
C4712 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_11629_12507# 0.02171f
C4713 a_17443_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.0394f
C4714 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 0.05869f
C4715 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 a_15593_6250# 0.02785f
C4716 a_44234_11946# a_43698_11746# 0.0139f
C4717 a_43698_10756# VDDH 0.24088f
C4718 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.05177f
C4719 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.06256f
C4720 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.02611f
C4721 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.04713f
C4722 VDDH a_2678_19053# 0.72825f
C4723 VDDH a_5897_14150# 0.49013f
C4724 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 0.02555f
C4725 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH 17.253f
C4726 a_39883_19854# a_39306_20477# 0.01316f
C4727 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 0.01984f
C4728 a_1636_13352# a_1636_13708# 0.02286f
C4729 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.63972f
C4730 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.12584f
C4731 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_15224_18696# 0.17206f
C4732 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C4733 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.14448f
C4734 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_31042_7686# 0.12972f
C4735 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.01068f
C4736 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.06167f
C4737 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_19946_8950# 0.02704f
C4738 a_39861_22496# ROUT2 0.13835f
C4739 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.01148f
C4740 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] VDDH 0.89706f
C4741 a_15629_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 0.03929f
C4742 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 1.60525f
C4743 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 0.02519f
C4744 a_21099_20174# a_21651_20174# 5.44167f
C4745 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 a_28882_6250# 0.02795f
C4746 a_24963_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 0.08492f
C4747 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 a_28172_6250# 0.02789f
C4748 a_43994_22522# a_44067_22496# 0.1148f
C4749 a_16891_7686# a_19946_8950# 0.03944f
C4750 VDDH top_DAC_0/top_rseg_n_dcell_0.SH[4] 1.34727f
C4751 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.0962f
C4752 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.0119f
C4753 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.1743f
C4754 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 0.15091f
C4755 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_20823_20174# 0.03457f
C4756 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 0.12185f
C4757 a_43698_15706# a_43724_15866# 0.02395f
C4758 VOUT a_4717_12507# 0.039f
C4759 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.08957f
C4760 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.03981f
C4761 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 0.17656f
C4762 a_14514_18696# a_17732_18696# 0.10942f
C4763 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.52521f
C4764 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_2678_21703# 0.03151f
C4765 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.03512f
C4766 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_5050_12595# 0.5224f
C4767 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.02785f
C4768 a_33634_8950# a_27896_6250# 0.08536f
C4769 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.06023f
C4770 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.06158f
C4771 VOUT a_11081_15057# 0.04641f
C4772 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 a_14607_6250# 0.02787f
C4773 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.11848f
C4774 a_43724_11906# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP 0.08245f
C4775 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.07771f
C4776 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.06276f
C4777 a_30608_7686# a_31042_7686# 6.27397f
C4778 a_30332_7686# a_31318_7686# 0.16296f
C4779 a_6778_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.17806f
C4780 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.05596f
C4781 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.02793f
C4782 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.06066f
C4783 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.15563f
C4784 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.64353f
C4785 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.09256f
C4786 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.04707f
C4787 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 0.06415f
C4788 VDDH top_DAC_0/top_final_switch_0.VOUT[0] 1.7051f
C4789 a_29434_6250# a_30056_7686# 0.04346f
C4790 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_final_switch_0.VOUT[4] 0.06879f
C4791 a_23859_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 0.06438f
C4792 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.05591f
C4793 VOUT a_7625_13005# 0.02203f
C4794 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.08875f
C4795 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.10018f
C4796 a_21099_20174# a_23031_20174# 0.13237f
C4797 a_20823_20174# a_23307_20174# 0.17716f
C4798 a_21375_20174# a_22755_20174# 0.20167f
C4799 a_21651_20174# a_22479_20174# 0.14085f
C4800 top_DAC_0/top_final_switch_0.VOUT[1] a_6445_13005# 0.02851f
C4801 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.02926f
C4802 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.02791f
C4803 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 0.02446f
C4804 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_2678_10356# 0.02628f
C4805 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 0.01848f
C4806 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 a_21927_20174# 0.04143f
C4807 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 a_24963_20174# 0.04155f
C4808 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 a_21651_20174# 0.04143f
C4809 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.07772f
C4810 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.02787f
C4811 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.11733f
C4812 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.17935f
C4813 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 0.01605f
C4814 a_20498_8950# a_20352_10031# 0.0771f
C4815 a_43698_11746# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.40164f
C4816 a_19946_8950# a_20932_10031# 0.06546f
C4817 a_20222_8950# a_20656_10031# 0.06662f
C4818 a_19670_8950# a_18724_8950# 0.09051f
C4819 a_19552_8950# a_19000_8950# 0.08347f
C4820 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 17.1095f
C4821 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.06124f
C4822 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_20352_10031# 0.07634f
C4823 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 a_27620_6250# 0.02788f
C4824 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 1.7572f
C4825 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.19025f
C4826 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 a_15317_6250# 0.02794f
C4827 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.68132f
C4828 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.22966f
C4829 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.02787f
C4830 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.04912f
C4831 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 a_27896_6250# 0.04435f
C4832 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 0.41945f
C4833 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB 0.01383f
C4834 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 a_27344_6250# 0.04219f
C4835 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_19552_8950# 0.02631f
C4836 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_17252# 0.0399f
C4837 a_44234_8342# a_44234_7986# 0.08026f
C4838 VDDH a_16891_7686# 0.50696f
C4839 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] VDDH 0.99488f
C4840 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.62483f
C4841 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.06065f
C4842 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.13647f
C4843 a_33634_8950# a_34186_8950# 0.08347f
C4844 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_5050_12595# 0.56145f
C4845 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.02784f
C4846 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.15222f
C4847 a_34304_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.02655f
C4848 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 0.09572f
C4849 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.64115f
C4850 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.02792f
C4851 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.55951f
C4852 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.11698f
C4853 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.0897f
C4854 a_15317_6250# a_13779_6250# 0.18926f
C4855 a_22479_20174# a_23031_20174# 0.13449f
C4856 a_22203_20174# a_23307_20174# 0.1772f
C4857 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_final_switch_0.VOUT[2] 0.06657f
C4858 a_35132_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.05484f
C4859 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44737_4828# 0.02083f
C4860 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_9966# 0.01697f
C4861 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_15906# 0.03152f
C4862 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.096f
C4863 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.98866f
C4864 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04791f
C4865 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 a_2678_16243# 0.0585f
C4866 a_23629_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.25057f
C4867 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.06231f
C4868 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_19946_8950# 0.05276f
C4869 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_27344_6250# 0.02393f
C4870 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.05173f
C4871 a_2300_13708# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.03745f
C4872 a_24135_20174# a_20547_20174# 0.13313f
C4873 a_23583_20174# a_21099_20174# 0.13228f
C4874 a_23049_18133# a_21375_20174# 0.01726f
C4875 a_23859_20174# a_20823_20174# 0.1713f
C4876 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.03927f
C4877 a_22469_18133# a_21651_20174# 0.04303f
C4878 a_38672_20477# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.37714f
C4879 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.57206f
C4880 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_6445_13005# 0.0208f
C4881 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 a_14331_6250# 0.03601f
C4882 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.3688f
C4883 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP 0.92839f
C4884 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.27627f
C4885 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_10322# 0.02378f
C4886 a_33358_8950# a_29780_7686# 0.03937f
C4887 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 0.05149f
C4888 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.17474f
C4889 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_5897_14150# 0.04959f
C4890 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 0.02587f
C4891 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.0279f
C4892 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 1.468f
C4893 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.14582f
C4894 a_43698_9766# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.24498f
C4895 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_5111_10963# 0.12264f
C4896 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 1.73307f
C4897 a_44062_22009# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.07788f
C4898 a_34856_8950# a_31870_7686# 0.07927f
C4899 VDDH a_4978_9535# 0.73032f
C4900 DIN1 VDD 0.66672f
C4901 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.09277f
C4902 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 3.02501f
C4903 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 0.0119f
C4904 VDDH a_20932_10031# 0.2897f
C4905 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.05356f
C4906 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 0.90356f
C4907 a_2678_20320# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 0.06368f
C4908 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD 0.18445f
C4909 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.11733f
C4910 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.01469f
C4911 a_8173_13005# top_DAC_0/top_final_switch_0.VOUT[2] 0.02847f
C4912 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_final_switch_0.VOUT[1] 0.17964f
C4913 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_24209_18133# 0.42857f
C4914 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.01814f
C4915 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05095f
C4916 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_final_switch_0.VOUT[1] 0.01422f
C4917 VDDH a_14331_6250# 0.71735f
C4918 a_14790_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.15324f
C4919 a_28172_6250# a_30332_7686# 0.04243f
C4920 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 a_20547_20174# 0.08782f
C4921 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_final_switch_0.VOUT[2] 0.04984f
C4922 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.07805f
C4923 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD a_11081_15057# 0.01033f
C4924 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN a_5111_10963# 0.08766f
C4925 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.1105f
C4926 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 a_16181_7686# 0.07965f
C4927 a_24135_20174# a_21927_20174# 0.13232f
C4928 a_23583_20174# a_22479_20174# 0.13258f
C4929 a_23859_20174# a_22203_20174# 0.15608f
C4930 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.02795f
C4931 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.22406f
C4932 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.16159f
C4933 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.02785f
C4934 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.01389f
C4935 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 1.39272f
C4936 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.26339f
C4937 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 0.06415f
C4938 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.VS1 0.07172f
C4939 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.1443f
C4940 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 0.82496f
C4941 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_34580_8950# 0.11475f
C4942 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN VDD 0.46252f
C4943 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 0.55358f
C4944 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_39306_20477# 0.76695f
C4945 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.06354f
C4946 a_43698_7786# a_43724_7946# 0.02395f
C4947 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A a_44234_7986# 0.05897f
C4948 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC a_37410_19098# 0.36169f
C4949 a_33634_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.24408f
C4950 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1 0.91031f
C4951 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A a_43724_8936# 0.08029f
C4952 a_24209_18133# a_23307_20174# 0.04111f
C4953 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_final_switch_0.VOUT[0] 0.20355f
C4954 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 3.49358f
C4955 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04366f
C4956 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 a_14331_6250# 0.08495f
C4957 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1896_16243# 0.0747f
C4958 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.VL3 0.1266f
C4959 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 0.55111f
C4960 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.15103f
C4961 a_30056_7686# a_27620_6250# 0.02786f
C4962 VDDH a_31870_7686# 0.09501f
C4963 a_29780_7686# a_27896_6250# 0.04211f
C4964 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 0.85518f
C4965 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 2.60553f
C4966 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 1.19856f
C4967 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 0.11518f
C4968 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 0.18788f
C4969 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 1.8445f
C4970 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_43698_6796# 0.01234f
C4971 VDDH a_5111_8388# 1.5705f
C4972 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.16919f
C4973 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.VL3 0.05876f
C4974 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 2.0654f
C4975 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.11522f
C4976 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 a_30056_7686# 0.07439f
C4977 VOUT a_11629_15057# 0.01454f
C4978 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.05438f
C4979 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.02766f
C4980 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.04787f
C4981 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.04807f
C4982 a_43698_6796# a_43724_7392# 0.06762f
C4983 a_16181_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.08f
C4984 a_19276_8950# a_19670_8950# 0.08334f
C4985 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.21135f
C4986 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.08499f
C4987 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.10618f
C4988 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.57437f
C4989 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 ROUT1 0.03407f
C4990 a_44234_14282# a_44234_14916# 0.02262f
C4991 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 a_13779_6250# 0.04211f
C4992 top_DAC_0/top_final_switch_0.VOUT[1] VOUT 6.36642f
C4993 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_43698_15706# 0.01234f
C4994 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB VOUT 2.66242f
C4995 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_final_switch_0.VOUT[2] 0.66459f
C4996 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 VDDH 0.10974f
C4997 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 0.0651f
C4998 a_43698_12736# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP 0.02263f
C4999 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_8506_12595# 1.28111f
C5000 a_15066_18696# a_15224_18696# 0.04177f
C5001 a_14514_18696# a_14672_18696# 0.04099f
C5002 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 3.39716f
C5003 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 2.6115f
C5004 a_14790_18696# a_14948_18696# 0.04033f
C5005 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.01144f
C5006 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.02784f
C5007 a_15593_6250# a_15869_6250# 7.25194f
C5008 a_15317_6250# a_15353_7686# 0.04654f
C5009 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43698_6796# 0.06167f
C5010 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.02359f
C5011 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.0848f
C5012 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.47364f
C5013 a_43698_16696# a_44062_18093# 0.03114f
C5014 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.83161f
C5015 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.06987f
C5016 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.21309f
C5017 a_44234_9966# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.35036f
C5018 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 1.95031f
C5019 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.09778f
C5020 a_35453_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.07622f
C5021 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_17252# 0.14701f
C5022 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.17603f
C5023 a_6778_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 0.20828f
C5024 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_24135_20174# 0.06448f
C5025 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 1.73087f
C5026 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.08427f
C5027 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.02197f
C5028 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.02163f
C5029 a_23859_20174# a_24209_18133# 0.0402f
C5030 a_44234_8976# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.06552f
C5031 a_34856_8950# a_28882_6250# 0.08494f
C5032 a_33910_8950# a_30056_7686# 0.08519f
C5033 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.26823f
C5034 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.03927f
C5035 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43698_15706# 0.06167f
C5036 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 17.4112f
C5037 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.01393f
C5038 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.04304f
C5039 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.06023f
C5040 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.43649f
C5041 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.10926f
C5042 a_39861_22057# a_39936_22083# 0.01759f
C5043 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_13926# 0.02704f
C5044 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.01136f
C5045 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 a_16320_18696# 0.04264f
C5046 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.10104f
C5047 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.09649f
C5048 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 a_28606_6250# 0.11031f
C5049 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 0.01616f
C5050 a_17732_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.11658f
C5051 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.09061f
C5052 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_final_switch_0.VOUT[3] 0.0444f
C5053 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 0.21355f
C5054 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15593_6250# 0.14215f
C5055 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.01346f
C5056 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.18005f
C5057 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02787f
C5058 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.0689f
C5059 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_14282# 0.03152f
C5060 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.04851f
C5061 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.03731f
C5062 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA VOUT 21.3105f
C5063 VDDH a_15905_7686# 0.48348f
C5064 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_18008_18696# 0.07973f
C5065 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_16872_18696# 0.01853f
C5066 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.13258f
C5067 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_31594_7686# 0.07511f
C5068 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 2.08874f
C5069 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.02214f
C5070 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.02426f
C5071 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.02179f
C5072 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 a_16872_18696# 0.06954f
C5073 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 a_16596_18696# 0.09104f
C5074 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.54398f
C5075 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 0.05523f
C5076 a_37595_19462# a_37595_19760# 0.015f
C5077 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 a_29434_6250# 0.20962f
C5078 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 0.14661f
C5079 a_18008_18696# top_DAC_0/top_rseg_n_dcell_0.VL3 0.44519f
C5080 a_20076_10031# a_20352_10031# 1.72453f
C5081 a_19772_10031# a_20656_10031# 0.35686f
C5082 VDDH top_DAC_0/top_final_switch_0.VOUT[2] 1.65987f
C5083 a_15863_13287# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.04291f
C5084 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.53572f
C5085 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.05759f
C5086 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01002f
C5087 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 0.01528f
C5088 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP 0.17284f
C5089 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.09525f
C5090 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.0857f
C5091 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.01153f
C5092 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.1245f
C5093 a_44234_11946# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.02704f
C5094 a_6923_9707# a_8506_12595# 0.12855f
C5095 top_DAC_0/top_rseg_n_dcell_0.VL2 a_14615_14034# 0.04303f
C5096 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.1324f
C5097 a_34873_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.27911f
C5098 a_9901_12507# a_9353_12507# 0.0103f
C5099 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.09544f
C5100 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_43698_11746# 0.01234f
C5101 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.1499f
C5102 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 3.61778f
C5103 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 1.75263f
C5104 top_DAC_0/top_rseg_n_dcell_0.VH3 a_21099_20174# 0.01023f
C5105 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 0.1105f
C5106 top_DAC_0/top_final_switch_0.VOUT[4] a_12809_12507# 0.01061f
C5107 a_33358_8950# a_34186_8950# 0.09218f
C5108 a_36033_10031# a_34304_8950# 0.04084f
C5109 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.03009f
C5110 a_35177_10031# a_35132_8950# 0.0581f
C5111 a_35453_10031# a_34856_8950# 0.04225f
C5112 a_35757_10031# a_34580_8950# 0.04106f
C5113 a_24963_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 0.08496f
C5114 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_19670_8950# 0.09441f
C5115 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.26787f
C5116 a_15618_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.0644f
C5117 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 0.01886f
C5118 a_43698_9766# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.78464f
C5119 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 17.1369f
C5120 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 a_23307_20174# 0.05523f
C5121 a_14948_18696# a_16872_18696# 0.08863f
C5122 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.0942f
C5123 a_14672_18696# a_16596_18696# 0.09029f
C5124 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_16262# 0.03855f
C5125 a_1896_10974# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 0.02981f
C5126 a_15863_13536# top_DAC_0/top_final_switch_0.VOUT[3] 0.02881f
C5127 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_14615_13785# 0.08429f
C5128 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 1.16507f
C5129 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 0.60003f
C5130 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 0.06445f
C5131 top_DAC_0/top_final_switch_0.VOUT[1] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.07333f
C5132 a_34580_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.1983f
C5133 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.11794f
C5134 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 0.5366f
C5135 a_43698_10756# a_43698_11746# 0.01563f
C5136 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] 0.08857f
C5137 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD a_5897_15057# 0.01037f
C5138 DIN2 VDD 0.66783f
C5139 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.04651f
C5140 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 0.01318f
C5141 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 0.07764f
C5142 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3 2.18169f
C5143 a_30056_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 0.04025f
C5144 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.04839f
C5145 VDDH top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 7.284f
C5146 a_22193_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.06552f
C5147 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.04691f
C5148 a_45023_18564# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.01005f
C5149 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43698_11746# 0.06167f
C5150 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_7986# 0.01407f
C5151 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 0.02042f
C5152 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.05186f
C5153 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_44062_18093# 0.06327f
C5154 a_2300_13352# a_2300_13708# 0.02286f
C5155 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_14672_18696# 0.30878f
C5156 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.VH3 0.95191f
C5157 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_31594_7686# 0.13361f
C5158 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.05177f
C5159 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 0.03773f
C5160 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 a_20823_20174# 0.06242f
C5161 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_20498_8950# 0.22951f
C5162 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 0.01733f
C5163 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 14.8638f
C5164 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.12455f
C5165 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.09973f
C5166 a_44067_22496# ROUT2 0.08397f
C5167 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.09117f
C5168 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.14241f
C5169 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 a_28606_6250# 0.02789f
C5170 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.03697f
C5171 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_8342# 0.01484f
C5172 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_30608_7686# 0.07822f
C5173 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 a_29434_6250# 0.04652f
C5174 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 0.78921f
C5175 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 a_29158_6250# 0.07771f
C5176 a_17167_7686# a_20222_8950# 0.03939f
C5177 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 a_28882_6250# 0.02795f
C5178 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 9.82232f
C5179 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 a_21099_20174# 0.06395f
C5180 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.15699f
C5181 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1636_15118# 0.03043f
C5182 a_11629_15057# a_11081_15057# 0.0237f
C5183 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 a_28606_6250# 0.03928f
C5184 a_31318_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.03929f
C5185 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.09237f
C5186 a_7625_14150# a_8173_14150# 0.0237f
C5187 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 a_21375_20174# 0.06393f
C5188 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] a_21375_20174# 0.23227f
C5189 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.12707f
C5190 a_24963_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.2027f
C5191 a_30608_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.07963f
C5192 a_43698_15706# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP 0.02263f
C5193 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.10438f
C5194 a_14790_18696# a_18008_18696# 0.06513f
C5195 a_15066_18696# a_17732_18696# 0.21441f
C5196 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.07481f
C5197 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 0.78185f
C5198 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 a_27344_6250# 0.0433f
C5199 a_15317_6250# a_16891_7686# 0.02803f
C5200 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_4717_12507# 0.02171f
C5201 a_15593_6250# a_16615_7686# 0.02792f
C5202 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 0.03979f
C5203 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 0.01515f
C5204 VOUT a_11081_14150# 0.06741f
C5205 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 0.02114f
C5206 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP 0.08366f
C5207 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 top_DAC_0/top_final_switch_0.VOUT[3] 0.20612f
C5208 a_31042_7686# a_31318_7686# 6.39975f
C5209 a_30608_7686# a_31594_7686# 0.16293f
C5210 a_30332_7686# a_31870_7686# 0.18046f
C5211 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.99952f
C5212 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_15863_13785# 0.02534f
C5213 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_28606_6250# 0.17608f
C5214 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.04338f
C5215 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 1.41618f
C5216 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] a_44062_21653# 0.02123f
C5217 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 1.51685f
C5218 VOUT a_12809_15057# 0.04557f
C5219 VOUT a_7625_12507# 0.04471f
C5220 a_33358_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.7782f
C5221 a_21651_20174# a_23031_20174# 0.13229f
C5222 a_21375_20174# a_23307_20174# 0.20149f
C5223 a_15863_13785# top_DAC_0/top_rseg_n_dcell_0.VL3 0.31264f
C5224 top_DAC_0/top_final_switch_0.VOUT[1] a_7625_13005# 0.03215f
C5225 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 0.01457f
C5226 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.12773f
C5227 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 0.0245f
C5228 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.04267f
C5229 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 49.343f
C5230 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] a_23031_20174# 0.03037f
C5231 a_8506_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 0.28554f
C5232 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.02787f
C5233 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 8.60462f
C5234 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 0.0106f
C5235 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.04054f
C5236 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.05217f
C5237 a_20498_8950# a_20932_10031# 0.02572f
C5238 a_19946_8950# a_19000_8950# 0.08886f
C5239 a_20222_8950# a_18724_8950# 0.0986f
C5240 a_6445_14150# VOUT 0.0409f
C5241 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.06107f
C5242 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 a_19670_8950# 0.02558f
C5243 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.39896f
C5244 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.08819f
C5245 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 a_20932_10031# 0.10734f
C5246 a_15374_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.04058f
C5247 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.05159f
C5248 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_final_switch_0.VOUT[2] 0.204f
C5249 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 a_27620_6250# 0.03777f
C5250 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 a_15869_6250# 0.04597f
C5251 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 a_27896_6250# 0.02784f
C5252 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 0.10155f
C5253 a_44234_8342# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.20594f
C5254 VDDH a_17443_7686# 0.86506f
C5255 a_34580_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.01396f
C5256 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y a_44062_19873# 0.09819f
C5257 a_15041_6250# a_19946_8950# 0.07768f
C5258 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 1.22987f
C5259 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B VDD 0.29366f
C5260 VDDH a_15224_18696# 0.27978f
C5261 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.54635f
C5262 a_33634_8950# a_34580_8950# 0.08886f
C5263 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.0142f
C5264 a_33910_8950# a_34304_8950# 0.08334f
C5265 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.02784f
C5266 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.14193f
C5267 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.10032f
C5268 a_34856_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.02898f
C5269 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.08294f
C5270 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.06017f
C5271 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 0.07844f
C5272 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 0.05789f
C5273 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.07846f
C5274 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.13238f
C5275 a_24963_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.11559f
C5276 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.33109f
C5277 a_15869_6250# a_13779_6250# 0.20768f
C5278 a_22755_20174# a_23307_20174# 0.17859f
C5279 a_15317_6250# a_14331_6250# 0.15576f
C5280 a_15593_6250# a_14055_6250# 0.15272f
C5281 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 0.71908f
C5282 VDDH a_20823_20174# 0.01605f
C5283 top_DAC_0/top_rseg_n_dcell_0.VH3 a_18008_18696# 0.36592f
C5284 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] a_14672_18696# 0.02448f
C5285 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.01807f
C5286 a_14615_14283# a_14615_14034# 0.11957f
C5287 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.97326f
C5288 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.1869f
C5289 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 a_15317_6250# 0.02795f
C5290 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_20498_8950# 0.06043f
C5291 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_27896_6250# 0.05568f
C5292 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.08441f
C5293 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.09178f
C5294 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.0636f
C5295 a_23583_20174# a_21651_20174# 0.13223f
C5296 a_23859_20174# a_21375_20174# 0.17638f
C5297 a_24135_20174# a_21099_20174# 0.1323f
C5298 a_24411_20174# a_20823_20174# 0.13242f
C5299 a_24687_20174# a_20547_20174# 0.13355f
C5300 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 0.03533f
C5301 a_31042_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.07987f
C5302 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.16622f
C5303 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 0.03939f
C5304 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA a_7625_13005# 0.0208f
C5305 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 a_14672_18696# 0.05354f
C5306 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 a_15041_6250# 0.03689f
C5307 a_44234_7986# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.06328f
C5308 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.43543f
C5309 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB 0.16457f
C5310 a_23049_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.36573f
C5311 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_15317_6250# 0.36298f
C5312 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.01782f
C5313 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_4978_10963# 0.01297f
C5314 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_16262# 0.14417f
C5315 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_43698_8776# 0.01234f
C5316 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.02791f
C5317 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 a_21099_20174# 0.06395f
C5318 VDDH a_19000_8950# 0.3363f
C5319 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.03392f
C5320 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 0.21553f
C5321 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 0.02514f
C5322 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 1.81409f
C5323 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 a_16615_7686# 0.07965f
C5324 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_13779_6250# 0.27901f
C5325 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 a_22755_20174# 0.05019f
C5326 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.30168f
C5327 a_44062_18449# a_44062_18093# 0.04238f
C5328 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 0.0485f
C5329 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.34328f
C5330 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 1.62525f
C5331 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 a_27620_6250# 0.02787f
C5332 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44479_4254# 0.01259f
C5333 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 2.48633f
C5334 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.17464f
C5335 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 1.8091f
C5336 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_1896_10356# 0.02965f
C5337 VDDH a_15041_6250# 0.83743f
C5338 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.04315f
C5339 a_1636_15118# VOUT 0.01189f
C5340 a_15342_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.37508f
C5341 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.01119f
C5342 VDDH a_8173_14150# 0.49013f
C5343 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 0.0484f
C5344 a_28606_6250# a_30608_7686# 0.04042f
C5345 a_28882_6250# a_30332_7686# 0.02798f
C5346 a_28172_6250# a_31042_7686# 0.0407f
C5347 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD 0.92259f
C5348 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 0.114f
C5349 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 a_22755_20174# 0.04147f
C5350 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_9926# 0.03597f
C5351 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A VDD 1.0555f
C5352 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 a_27896_6250# 0.08515f
C5353 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.0908f
C5354 top_DAC_0/top_final_switch_0.VOUT[4] top_DAC_0/top_final_switch_0.VOUT[3] 5.50358f
C5355 a_23583_20174# a_23031_20174# 0.13358f
C5356 a_24687_20174# a_21927_20174# 0.13238f
C5357 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB VDD 0.89598f
C5358 a_24411_20174# a_22203_20174# 0.13241f
C5359 a_23859_20174# a_22755_20174# 0.15428f
C5360 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.04713f
C5361 a_24135_20174# a_22479_20174# 0.13249f
C5362 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 0.11371f
C5363 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 a_15317_6250# 0.02784f
C5364 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.02785f
C5365 a_38672_20477# a_37410_19098# 1.49212f
C5366 a_44062_20585# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.02354f
C5367 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 1.33001f
C5368 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP 0.34417f
C5369 a_44234_15272# a_44234_14916# 0.08026f
C5370 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43698_8776# 0.06167f
C5371 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_35132_8950# 0.1733f
C5372 a_19468_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.22424f
C5373 a_44234_14282# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.08438f
C5374 a_34186_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.09456f
C5375 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 1.29067f
C5376 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 0.09809f
C5377 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.08251f
C5378 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.03899f
C5379 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 1.03522f
C5380 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.14118f
C5381 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 3.43068f
C5382 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 0.04346f
C5383 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.03202f
C5384 a_17148_18696# a_15224_18696# 0.09841f
C5385 VDDH a_4978_8388# 0.79433f
C5386 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.19453f
C5387 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 0.02803f
C5388 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.38434f
C5389 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.28823f
C5390 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.04702f
C5391 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.03108f
C5392 a_16615_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.07989f
C5393 a_43698_6796# a_44234_6996# 0.0139f
C5394 a_17167_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.03944f
C5395 a_19276_8950# a_20222_8950# 0.08895f
C5396 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.02784f
C5397 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 0.15742f
C5398 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 a_14331_6250# 0.02784f
C5399 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.33061f
C5400 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_final_switch_0.VOUT[1] 0.20372f
C5401 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_14916# 0.02704f
C5402 a_15863_13785# top_DAC_0/top_rseg_n_dcell_0.VH3 0.04213f
C5403 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.0396f
C5404 a_6445_12507# a_5897_12507# 0.0103f
C5405 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.0119f
C5406 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 0.06117f
C5407 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 a_15869_6250# 0.03934f
C5408 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.04487f
C5409 a_15869_6250# a_15353_7686# 0.21158f
C5410 a_15593_6250# a_15629_7686# 0.02792f
C5411 a_15317_6250# a_15905_7686# 0.02801f
C5412 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_20076_10031# 0.24001f
C5413 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_final_switch_0.VOUT[2] 0.17964f
C5414 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 a_28172_6250# 0.03939f
C5415 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_15272# 0.03152f
C5416 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.0979f
C5417 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.05175f
C5418 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.06278f
C5419 a_36033_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.10609f
C5420 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.23994f
C5421 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN a_44234_6996# 0.07516f
C5422 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.05086f
C5423 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 1.47682f
C5424 VDDH a_17732_18696# 0.21696f
C5425 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_14514_18696# 0.07274f
C5426 a_14615_14283# top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.05354f
C5427 a_35132_8950# a_29158_6250# 0.11034f
C5428 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.01172f
C5429 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 0.05095f
C5430 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 a_31594_7686# 0.07165f
C5431 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.67152f
C5432 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.17756f
C5433 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.02784f
C5434 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 VDDH 0.20568f
C5435 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 8.31228f
C5436 a_13779_6250# a_16615_7686# 0.0317f
C5437 top_DAC_0/top_rseg_n_dcell_0.VL3 top_DAC_0/top_final_switch_0.VOUT[1] 0.03452f
C5438 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y VDD 0.41365f
C5439 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04066f
C5440 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.02029f
C5441 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_41907_22057# 0.02974f
C5442 a_43698_12736# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP 0.7858f
C5443 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.14375f
C5444 a_18284_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.57739f
C5445 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.01905f
C5446 VDDH a_43698_13726# 0.24088f
C5447 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.02791f
C5448 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15353_7686# 0.19331f
C5449 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.16177f
C5450 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 12.0047f
C5451 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 0.11461f
C5452 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02789f
C5453 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.01647f
C5454 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] 17.521f
C5455 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 0.14514f
C5456 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 1.37192f
C5457 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 0.09544f
C5458 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA a_5897_15057# 0.04959f
C5459 a_16615_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.07612f
C5460 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.36098f
C5461 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.VL3 0.68768f
C5462 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA top_DAC_0/top_final_switch_0.VOUT[1] 0.39674f
C5463 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA 13.196f
C5464 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.0977f
C5465 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 0.053f
C5466 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB a_8173_14150# 0.04994f
C5467 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 3.4669f
C5468 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 0.05183f
C5469 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.26998f
C5470 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.36163f
C5471 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09291f
C5472 top_DAC_0/top_rseg_n_dcell_0.VS1 top_DAC_0/top_final_switch_0.VOUT[4] 0.10469f
C5473 DIN1 VDDH 0.42749f
C5474 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.01034f
C5475 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 0.26736f
C5476 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.41078f
C5477 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 0.03299f
C5478 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 0.0145f
C5479 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.05053f
C5480 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.06395f
C5481 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 0.0641f
C5482 a_20352_10031# a_20656_10031# 1.3412f
C5483 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 0.08504f
C5484 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 a_30056_7686# 0.07245f
C5485 a_20076_10031# a_20932_10031# 0.0881f
C5486 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.20535f
C5487 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.02787f
C5488 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 0.26016f
C5489 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 a_14055_6250# 0.02787f
C5490 a_43698_14716# a_43724_15312# 0.06762f
C5491 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.0707f
C5492 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 a_21375_20174# 0.0516f
C5493 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.0421f
C5494 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 0.09454f
C5495 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.12612f
C5496 a_35177_10031# a_34569_10031# 0.17353f
C5497 a_35453_10031# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.08763f
C5498 top_DAC_0/top_rseg_n_dcell_0.VL2 a_14615_13536# 0.12589f
C5499 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.0119f
C5500 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_44062_19873# 0.06327f
C5501 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_13886# 0.03597f
C5502 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.06069f
C5503 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 a_28882_6250# 0.03939f
C5504 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 0.01938f
C5505 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 0.09592f
C5506 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 a_28172_6250# 0.1105f
C5507 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.03958f
C5508 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.13739f
C5509 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.1481f
C5510 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 0.02577f
C5511 a_15374_19866# a_15224_18696# 1.96272f
C5512 a_33358_8950# a_34580_8950# 0.09965f
C5513 a_35757_10031# a_35132_8950# 0.01845f
C5514 a_15098_19866# a_14948_18696# 0.21748f
C5515 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.04121f
C5516 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 a_20222_8950# 0.11773f
C5517 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.72578f
C5518 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 1.38173f
C5519 a_13779_6250# a_14055_6250# 7.36324f
C5520 a_34856_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.0268f
C5521 DIN0 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.18007f
C5522 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.02015f
C5523 a_15098_19866# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.06346f
C5524 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 a_31042_7686# 0.07987f
C5525 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.11409f
C5526 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.05999f
C5527 a_16320_18696# a_16872_18696# 0.09034f
C5528 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_final_switch_0.VOUT[3] 0.06661f
C5529 a_43698_7786# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.40011f
C5530 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] 0.04064f
C5531 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 a_14948_18696# 0.04815f
C5532 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 1.9819f
C5533 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 1.32352f
C5534 a_35132_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.1896f
C5535 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.04506f
C5536 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_20076_10031# 0.06754f
C5537 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 17.3231f
C5538 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 0.01993f
C5539 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.0706f
C5540 a_43724_12896# VDDH 0.09227f
C5541 VDDH top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 4.26993f
C5542 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 0.79196f
C5543 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_9966# 0.0248f
C5544 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A a_43724_10362# 0.03253f
C5545 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] VDD 3.68198f
C5546 a_14055_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.21631f
C5547 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.1029f
C5548 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.08972f
C5549 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 1.90818f
C5550 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] 0.11733f
C5551 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.07187f
C5552 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.97341f
C5553 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD 1.19048f
C5554 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.05025f
C5555 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.12942f
C5556 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_16596_18696# 0.21399f
C5557 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.0525f
C5558 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_19946_8950# 0.05191f
C5559 a_23031_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 0.06399f
C5560 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 a_21651_20174# 0.06393f
C5561 a_43724_11906# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.03597f
C5562 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 1.32046f
C5563 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV ROUT2 0.25958f
C5564 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 1.859f
C5565 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.11848f
C5566 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 a_29158_6250# 0.02794f
C5567 a_1896_19053# a_2678_19053# 0.02127f
C5568 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_31318_7686# 0.07576f
C5569 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.1529f
C5570 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 a_28606_6250# 0.04067f
C5571 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 a_30056_7686# 0.04025f
C5572 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.02948f
C5573 a_39861_22057# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.03219f
C5574 a_17443_7686# a_20498_8950# 0.04142f
C5575 a_15863_13287# top_DAC_0/top_final_switch_0.VOUT[1] 0.01089f
C5576 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 a_29434_6250# 0.04713f
C5577 a_22193_18133# a_20823_20174# 0.09255f
C5578 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A a_1636_14353# 0.03043f
C5579 a_11629_14150# top_DAC_0/top_final_switch_0.VOUT[3] 0.01208f
C5580 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] ROUT2 0.0162f
C5581 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 0.53743f
C5582 a_23583_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.03017f
C5583 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.02726f
C5584 top_DAC_0/top_rseg_n_dcell_0.SH[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.04779f
C5585 a_44234_7352# a_44234_7986# 0.02262f
C5586 a_15618_18696# a_17732_18696# 0.03512f
C5587 a_15342_18696# a_18008_18696# 0.17363f
C5588 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 1.23264f
C5589 a_15066_18696# a_18284_18696# 0.27847f
C5590 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 1.88113f
C5591 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.02001f
C5592 a_15869_6250# a_16891_7686# 0.03865f
C5593 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] 0.03552f
C5594 a_15317_6250# a_17443_7686# 0.05563f
C5595 a_15593_6250# a_17167_7686# 0.02797f
C5596 a_15353_7686# a_16615_7686# 0.20741f
C5597 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP 0.10923f
C5598 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.23232f
C5599 VDD top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 1.81308f
C5600 a_23629_18133# a_20547_20174# 0.06807f
C5601 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 1.61342f
C5602 a_31042_7686# a_31870_7686# 0.18186f
C5603 a_31318_7686# a_31594_7686# 6.46593f
C5604 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.04851f
C5605 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.59734f
C5606 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_29158_6250# 0.38764f
C5607 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.13293f
C5608 a_43698_14716# a_44234_14916# 0.0139f
C5609 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] 0.04329f
C5610 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44062_18093# 0.02575f
C5611 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 17.0519f
C5612 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 VDDH 0.11183f
C5613 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_7946# 0.03597f
C5614 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD VOUT 0.6262f
C5615 a_24687_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3 0.07772f
C5616 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.56413f
C5617 VOUT a_12809_14150# 0.06888f
C5618 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.20664f
C5619 a_15863_13287# top_DAC_0/top_rseg_n_dcell_0.VL3 0.35551f
C5620 top_DAC_0/top_final_switch_0.VOUT[1] a_7625_12507# 0.01061f
C5621 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 a_16596_18696# 0.0397f
C5622 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB a_7625_12507# 0.0208f
C5623 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.16266f
C5624 a_44234_10322# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.32991f
C5625 a_43698_16696# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.01132f
C5626 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.48051f
C5627 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_final_switch_0.VOUT[1] 0.01731f
C5628 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 0.1185f
C5629 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.04473f
C5630 a_15353_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.04539f
C5631 a_20498_8950# a_19000_8950# 0.10087f
C5632 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 VDDH 3.72704f
C5633 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 0.01692f
C5634 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_16891_7686# 0.11955f
C5635 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 a_15629_7686# 0.04025f
C5636 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 a_22203_20174# 0.07766f
C5637 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.11733f
C5638 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_final_switch_0.VOUT[0] 0.08765f
C5639 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.09326f
C5640 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.03991f
C5641 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_30608_7686# 0.1145f
C5642 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 0.54188f
C5643 a_23629_18133# a_21927_20174# 0.04357f
C5644 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 2.2876f
C5645 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_20498_8950# 0.20443f
C5646 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 0.47f
C5647 VDDH top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 4.40766f
C5648 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 0.6725f
C5649 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 0.32234f
C5650 VDDH a_14672_18696# 0.54064f
C5651 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 a_28606_6250# 0.03788f
C5652 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_final_switch_0.VOUT[3] 0.01325f
C5653 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 1.24741f
C5654 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 top_DAC_0/top_rseg_n_dcell_0.VH3 1.53928f
C5655 a_33634_8950# a_35132_8950# 0.10144f
C5656 a_34186_8950# a_34580_8950# 0.09177f
C5657 a_33910_8950# a_34856_8950# 0.08895f
C5658 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 0.05729f
C5659 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.04735f
C5660 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.02218f
C5661 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 0.10984f
C5662 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.17853f
C5663 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] ROUT2 0.02421f
C5664 a_13779_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.12187f
C5665 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.1319f
C5666 a_15869_6250# a_14331_6250# 0.17275f
C5667 a_15317_6250# a_15041_6250# 7.37047f
C5668 a_15629_7686# a_13779_6250# 0.03168f
C5669 a_15353_7686# a_14055_6250# 0.04204f
C5670 a_15593_6250# a_14607_6250# 0.16424f
C5671 a_30608_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.02898f
C5672 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.04792f
C5673 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 1.16961f
C5674 a_44062_20585# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.07788f
C5675 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_43698_14716# 0.01234f
C5676 top_DAC_0/top_rseg_n_dcell_0.VH3 top_DAC_0/top_rseg_n_dcell_0.VL3 2.98928f
C5677 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 1.57642f
C5678 a_14615_14034# a_14615_13785# 0.11905f
C5679 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 0.05594f
C5680 a_9353_13005# a_9901_13005# 0.0103f
C5681 a_8506_12595# a_8051_10107# 1.49673f
C5682 a_14514_18696# a_15066_18696# 0.10242f
C5683 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 a_15869_6250# 0.04707f
C5684 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 a_31318_7686# 0.07419f
C5685 VDDH a_36888_19550# 0.01826f
C5686 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.09312f
C5687 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 a_6923_9707# 0.21493f
C5688 a_24687_20174# a_21099_20174# 0.13231f
C5689 a_24135_20174# a_21651_20174# 0.13227f
C5690 a_24963_20174# a_20823_20174# 0.13307f
C5691 a_24411_20174# a_21375_20174# 0.14451f
C5692 a_29158_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.45348f
C5693 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.01212f
C5694 a_4717_15057# top_DAC_0/top_final_switch_0.VOUT[0] 0.03029f
C5695 a_15629_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.0825f
C5696 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.VS4 0.14409f
C5697 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.04811f
C5698 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 0.25882f
C5699 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.06121f
C5700 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 1.37492f
C5701 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_28172_6250# 0.15401f
C5702 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 0.0961f
C5703 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_15869_6250# 0.48286f
C5704 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 a_15224_18696# 0.04732f
C5705 a_43698_7786# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.24498f
C5706 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.09743f
C5707 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04882f
C5708 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.04847f
C5709 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.69539f
C5710 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 8.44169f
C5711 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.20262f
C5712 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 0.01944f
C5713 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.14521f
C5714 a_28882_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 0.02794f
C5715 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 0.02163f
C5716 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_14615_14034# 0.02215f
C5717 a_28172_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 0.02787f
C5718 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 0.19029f
C5719 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43698_14716# 0.06167f
C5720 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.21128f
C5721 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_13926# 0.03855f
C5722 a_22193_18133# a_24209_18133# 0.4446f
C5723 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax 1.45233f
C5724 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_14331_6250# 0.19215f
C5725 DIN2 VDDH 0.42749f
C5726 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44062_21297# 0.01675f
C5727 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 a_27344_6250# 0.04304f
C5728 a_2678_20320# a_1896_20320# 0.02127f
C5729 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_9966# 0.1344f
C5730 a_45343_4538# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.01159f
C5731 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 0.04635f
C5732 a_23859_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 0.06393f
C5733 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 a_27620_6250# 0.02787f
C5734 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 0.12231f
C5735 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 1.5609f
C5736 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.05594f
C5737 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_43698_16696# 0.29584f
C5738 a_43698_12736# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.01234f
C5739 a_1636_14353# VOUT 0.02722f
C5740 a_28882_6250# a_31042_7686# 0.02799f
C5741 a_28172_6250# a_31594_7686# 0.0504f
C5742 a_29434_6250# a_30332_7686# 0.04224f
C5743 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.03409f
C5744 a_28606_6250# a_31318_7686# 0.05423f
C5745 a_29158_6250# a_30608_7686# 0.02791f
C5746 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.05628f
C5747 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.10315f
C5748 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 top_DAC_0/top_rseg_n_dcell_0.VS1 0.07459f
C5749 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 a_34569_10031# 0.06169f
C5750 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 0.02291f
C5751 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.10068f
C5752 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.18856f
C5753 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A VDD 0.59039f
C5754 DIN4 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.01591f
C5755 a_24963_20174# a_22203_20174# 0.13327f
C5756 a_24135_20174# a_23031_20174# 0.12545f
C5757 a_23859_20174# a_23307_20174# 0.15372f
C5758 a_24687_20174# a_22479_20174# 0.13329f
C5759 a_24411_20174# a_22755_20174# 0.13313f
C5760 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 a_15869_6250# 0.04086f
C5761 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.04268f
C5762 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP a_43724_13332# 0.03147f
C5763 a_29434_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.04345f
C5764 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 a_19670_8950# 0.45875f
C5765 a_38584_20389# a_37410_19098# 0.01751f
C5766 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 9.1182f
C5767 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 0.16031f
C5768 VDDH top_DAC_0/top_final_switch_0.VOUT[3] 1.66679f
C5769 a_15863_13536# top_DAC_0/top_rseg_n_dcell_0.SH[3] 0.08809f
C5770 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.05882f
C5771 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 0.11838f
C5772 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.09286f
C5773 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 a_20547_20174# 0.01571f
C5774 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.578f
C5775 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.04259f
C5776 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.04811f
C5777 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_27344_6250# 0.8572f
C5778 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 a_21927_20174# 0.07411f
C5779 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD 0.14299f
C5780 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.02204f
C5781 a_23629_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.36919f
C5782 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD 0.21766f
C5783 a_34580_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 0.1181f
C5784 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.02298f
C5785 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] 0.32857f
C5786 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.01055f
C5787 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.06788f
C5788 top_DAC_0/top_final_switch_0.VOUT[2] a_9353_13005# 0.03212f
C5789 a_16615_7686# a_16891_7686# 6.2418f
C5790 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 3.3366f
C5791 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 a_5111_8388# 0.01452f
C5792 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.04875f
C5793 a_44234_11946# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.03855f
C5794 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] a_14948_18696# 0.11443f
C5795 a_43698_12736# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.06167f
C5796 a_17148_18696# a_14672_18696# 0.0987f
C5797 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.09548f
C5798 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.30979f
C5799 VDDH a_43724_9372# 0.09227f
C5800 ROUT1 VDD 0.68441f
C5801 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.SH[4] 0.04736f
C5802 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 0.03386f
C5803 a_27896_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 0.02788f
C5804 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.01125f
C5805 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.08136f
C5806 a_27344_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.05702f
C5807 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 0.0119f
C5808 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 a_15317_6250# 0.02795f
C5809 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44479_4170# 0.01118f
C5810 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A a_43724_6956# 0.08029f
C5811 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 0.22699f
C5812 VDDH a_6445_15057# 0.49751f
C5813 a_15869_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.04086f
C5814 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 0.07345f
C5815 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.20079f
C5816 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 a_15041_6250# 0.02785f
C5817 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 0.13121f
C5818 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.10895f
C5819 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 5.80789f
C5820 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN a_5111_8388# 0.12726f
C5821 a_15863_13287# top_DAC_0/top_rseg_n_dcell_0.VH3 0.04205f
C5822 a_14790_18696# a_16872_18696# 0.04596f
C5823 a_15618_18696# a_14672_18696# 0.04765f
C5824 a_15066_18696# a_16596_18696# 0.04642f
C5825 a_15342_18696# a_16320_18696# 0.04684f
C5826 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 0.57403f
C5827 top_DAC_0/top_rseg_n_dcell_0.VS4 top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.06264f
C5828 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 0.05777f
C5829 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 a_15863_13536# 0.16112f
C5830 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.02801f
C5831 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.13332f
C5832 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 0.63136f
C5833 a_15353_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 0.01086f
C5834 a_23583_20174# a_24135_20174# 5.57273f
C5835 a_23049_18133# a_24411_20174# 0.06945f
C5836 a_15353_7686# a_15629_7686# 6.37593f
C5837 a_15593_6250# a_16181_7686# 0.02791f
C5838 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 a_28172_6250# 0.02789f
C5839 a_15869_6250# a_15905_7686# 0.0422f
C5840 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP a_43724_14322# 0.03147f
C5841 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 0.05702f
C5842 a_43698_13726# a_44234_14282# 0.07082f
C5843 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 a_20656_10031# 0.34808f
C5844 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.04863f
C5845 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] a_44234_7986# 0.01278f
C5846 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 a_4978_11461# 0.06246f
C5847 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.47348f
C5848 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 0.02792f
C5849 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 0.05769f
C5850 a_6778_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 0.2492f
C5851 DIN4 VDD 0.67214f
C5852 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.11249f
C5853 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.07957f
C5854 a_1896_10974# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.02584f
C5855 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.02913f
C5856 a_30608_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.03222f
C5857 a_37595_19760# a_36888_19786# 0.0296f
C5858 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.02794f
C5859 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.07407f
C5860 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] a_15066_18696# 0.05817f
C5861 VDDH a_18284_18696# 0.19772f
C5862 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.09112f
C5863 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 0.03176f
C5864 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] 0.05868f
C5865 a_14615_13785# top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.05632f
C5866 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP a_43724_16302# 0.03147f
C5867 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 a_15593_6250# 0.0534f
C5868 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 a_15593_6250# 0.02794f
C5869 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.19372f
C5870 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.18193f
C5871 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 0.02394f
C5872 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.03927f
C5873 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 0.06214f
C5874 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.02784f
C5875 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.09304f
C5876 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 0.0266f
C5877 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 a_21927_20174# 0.0741f
C5878 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] a_27344_6250# 0.10609f
C5879 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 0.06197f
C5880 a_14331_6250# a_16615_7686# 0.02793f
C5881 a_13779_6250# a_17167_7686# 0.03173f
C5882 a_14055_6250# a_16891_7686# 0.02791f
C5883 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 0.0119f
C5884 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 0.68159f
C5885 a_11081_13005# top_DAC_0/top_final_switch_0.VOUT[3] 0.03209f
C5886 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.02885f
C5887 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.06438f
C5888 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 5.06241f
C5889 a_5050_12595# a_8506_12595# 0.09543f
C5890 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_40525_21457# 0.0755f
C5891 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.19079f
C5892 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_43724_14876# 0.03597f
C5893 a_43698_14716# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP 0.7858f
C5894 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.02791f
C5895 a_28172_6250# a_28606_6250# 6.24348f
C5896 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 a_15905_7686# 0.12266f
C5897 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.09058f
C5898 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.02124f
C5899 a_35132_8950# top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.03984f
C5900 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.09784f
C5901 a_6923_9707# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 5.66494f
C5902 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 2.49981f
C5903 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 1.1544f
C5904 a_17167_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.07246f
C5905 VDDH top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 0.10923f
C5906 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 0.77295f
C5907 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] 17.6537f
C5908 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 0.14327f
C5909 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_16615_7686# 0.08053f
C5910 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] 0.05912f
C5911 a_30608_7686# a_27344_6250# 0.03759f
C5912 a_30332_7686# a_27620_6250# 0.02787f
C5913 VOUT a_9901_12507# 0.03463f
C5914 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.03662f
C5915 a_20656_10031# a_20932_10031# 0.93546f
C5916 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 a_19772_10031# 0.19852f
C5917 a_15041_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.03927f
C5918 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_13926# 0.14379f
C5919 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 0.35106f
C5920 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 a_14607_6250# 0.03308f
C5921 a_27620_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 0.02786f
C5922 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB top_DAC_0/top_final_switch_0.VOUT[3] 0.20445f
C5923 a_44234_8342# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.06548f
C5924 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB DIN2 0.01828f
C5925 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 a_20076_10031# 0.15786f
C5926 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.11724f
C5927 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.05586f
C5928 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 0.02493f
C5929 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 0.02615f
C5930 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.01429f
C5931 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 0.09533f
C5932 a_35757_10031# a_34569_10031# 0.06176f
C5933 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_20823_20174# 0.032f
C5934 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.05175f
C5935 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44234_7352# 0.01488f
C5936 a_13779_6250# a_18724_8950# 0.03917f
C5937 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.13009f
C5938 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] 0.14315f
C5939 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 0.54335f
C5940 VDDH a_2678_17510# 0.72716f
C5941 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 1.96808f
C5942 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 1.1774f
C5943 a_15098_19866# a_16320_18696# 0.10129f
C5944 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.20923f
C5945 a_15374_19866# a_14672_18696# 0.1572f
C5946 a_33358_8950# a_35132_8950# 0.14481f
C5947 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 a_16615_7686# 0.03929f
C5948 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.01782f
C5949 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.28212f
C5950 a_2678_20320# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 0.05095f
C5951 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] 0.05538f
C5952 a_45015_4828# VDD 0.03791f
C5953 a_14055_6250# a_14331_6250# 7.41706f
C5954 a_13779_6250# a_14607_6250# 0.33317f
C5955 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.02139f
C5956 a_14514_18696# VDDH 0.5807f
C5957 top_DAC_0/top_final_switch_0.VOUT[0] top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA 0.59483f
C5958 a_18724_8950# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.01984f
C5959 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 0.09649f
C5960 a_14331_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 0.08519f
C5961 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.38843f
C5962 a_15593_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 0.06292f
C5963 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 a_14055_6250# 0.02787f
C5964 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_20656_10031# 0.06707f
C5965 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 0.1725f
C5966 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y a_45015_4828# 0.02202f
C5967 a_43724_10916# VDDH 0.09227f
C5968 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] a_45343_4828# 0.01631f
C5969 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A a_44234_9966# 0.05898f
C5970 a_44234_11946# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.14379f
C5971 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 1.90588f
C5972 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.01833f
C5973 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 0.32165f
C5974 a_14607_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.56697f
C5975 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 0.02493f
C5976 a_39883_19098# a_37410_19098# 0.04493f
C5977 a_43698_10756# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP 0.7858f
C5978 a_33910_8950# a_30332_7686# 0.03932f
C5979 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] a_18008_18696# 0.06145f
C5980 top_DAC_0/top_rseg_n_dcell_0.SH[3] top_DAC_0/top_final_switch_0.VOUT[4] 0.06643f
C5981 a_15066_18696# top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] 0.07973f
C5982 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] a_22203_20174# 0.03274f
C5983 a_15317_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.08551f
C5984 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 0.01393f
C5985 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 a_14055_6250# 0.15706f
C5986 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 1.15664f
C5987 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] a_44062_19873# 0.02511f
C5988 a_5111_10963# VOUT 0.01183f
C5989 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_20498_8950# 0.07294f
C5990 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.29658f
C5991 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 0.05185f
C5992 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] 0.69498f
C5993 VDDH a_15863_13536# 0.14137f
C5994 a_14615_14034# top_DAC_0/top_final_switch_0.VOUT[2] 0.06266f
C5995 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 a_16872_18696# 0.06383f
C5996 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.55748f
C5997 a_16615_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.03947f
C5998 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 a_14607_6250# 0.11032f
C5999 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 0.09994f
C6000 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 0.12119f
C6001 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] a_31870_7686# 0.08367f
C6002 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 a_29158_6250# 0.04485f
C6003 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 3.04089f
C6004 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 1.09792f
C6005 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN a_44234_15272# 0.08412f
C6006 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.54465f
C6007 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04786f
C6008 a_22193_18133# a_21375_20174# 0.05477f
C6009 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.0923f
C6010 DIN5 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.17945f
C6011 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 a_15317_6250# 0.19967f
C6012 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] 0.09076f
C6013 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 1.32022f
C6014 a_24135_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] 0.03011f
C6015 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 0.01833f
C6016 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 0.45968f
C6017 a_44234_7352# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.06689f
C6018 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 0.0191f
C6019 VDDH a_9901_14150# 0.49013f
C6020 a_15618_18696# a_18284_18696# 0.17347f
C6021 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 5.28584f
C6022 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 0.20703f
C6023 a_15905_7686# a_16615_7686# 0.17054f
C6024 a_15629_7686# a_16891_7686# 0.16163f
C6025 a_15869_6250# a_17443_7686# 0.05574f
C6026 a_15353_7686# a_17167_7686# 0.2168f
C6027 a_22469_18133# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.08701f
C6028 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 top_DAC_0/top_rseg_n_dcell_0.SH[2] 0.05175f
C6029 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB a_44234_7352# 0.08225f
C6030 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 0.01252f
C6031 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_44234_7986# 0.1344f
C6032 a_23629_18133# a_21099_20174# 0.06936f
C6033 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 1.27443f
C6034 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 a_14055_6250# 0.02784f
C6035 a_28606_6250# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 0.03939f
C6036 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] VDD 1.96314f
C6037 a_31594_7686# a_31870_7686# 6.57223f
C6038 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 2.07263f
C6039 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] a_44234_13292# 0.02704f
C6040 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.1148f
C6041 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 1.22509f
C6042 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] a_29780_7686# 0.55934f
C6043 VOUT top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B 0.65147f
C6044 VDDH VDD 5.24685f
C6045 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP a_43724_14876# 0.08245f
C6046 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax a_1896_11886# 0.02366f
C6047 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 1.97214f
C6048 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] 0.05283f
C6049 top_DAC_0/top_rseg_n_dcell_0.VL2 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 0.07746f
C6050 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 0.0555f
C6051 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD 0.11834f
C6052 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_36888_19786# 0.01362f
C6053 top_DAC_0/top_rseg_n_dcell_0.VH2 top_DAC_0/top_rseg_n_dcell_0.VL2 5.30487f
C6054 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.20641f
C6055 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 0.18431f
C6056 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD top_DAC_0/top_final_switch_0.VOUT[1] 0.59768f
C6057 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 2.15109f
C6058 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.08655f
C6059 a_44062_20229# a_44062_19873# 0.04541f
C6060 a_22193_18133# a_22755_20174# 0.09203f
C6061 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN VDD 0.45307f
C6062 a_24411_20174# top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 0.04148f
C6063 a_34873_10031# a_35177_10031# 0.26171f
C6064 a_1896_10356# top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx 0.05988f
C6065 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.0761f
C6066 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.08602f
C6067 VDDH a_7625_15057# 0.49751f
C6068 a_19552_8950# a_19946_8950# 0.09177f
C6069 a_44234_11312# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.09046f
C6070 a_8506_12595# top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 0.61545f
C6071 a_44234_6996# top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.07278f
C6072 VDDH top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 11.2804f
C6073 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] top_DAC_0/top_rseg_n_dcell_0.SH[1] 0.062f
C6074 a_29780_7686# top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 0.04526f
C6075 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 0.11409f
C6076 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.09546f
C6077 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 0.03606f
C6078 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 a_34569_10031# 0.22831f
C6079 DIN9 GND 2.58682f
C6080 DIN8 GND 2.24158f
C6081 DIN7 GND 2.21448f
C6082 DIN6 GND 2.18502f
C6083 DIN5 GND 2.16664f
C6084 DIN4 GND 2.15816f
C6085 DIN3 GND 2.13965f
C6086 DIN2 GND 2.11716f
C6087 DIN1 GND 2.1019f
C6088 DIN0 GND 2.34399f
C6089 VOUT GND 41.0058f
C6090 ROUT2 GND 13.7344f
C6091 ROUT1 GND 14.7092f
C6092 VDD GND 0.15211p
C6093 VDDH GND 0.76935p
C6094 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B GND 0.39231f
C6095 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y GND 0.3768f
C6096 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A GND 0.68099f
C6097 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y GND 0.70838f
C6098 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C GND 0.3332f
C6099 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B GND 0.32574f
C6100 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B GND 0.31137f
C6101 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A GND 0.25769f
C6102 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A GND 0.32968f
C6103 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y GND 0.45293f
C6104 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C GND 0.41678f
C6105 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B GND 0.42992f
C6106 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y GND 0.33977f
C6107 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A GND 0.73456f
C6108 a_45343_4828# GND 0.02142f $ **FLOATING
C6109 a_44471_4828# GND 0.02172f $ **FLOATING
C6110 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B GND 0.44413f
C6111 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A GND 0.49956f
C6112 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v55 GND 1.58565f
C6113 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v54 GND 1.01698f
C6114 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v53 GND 0.83396f
C6115 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v52 GND 0.84338f
C6116 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v51 GND 0.72928f
C6117 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v50 GND 0.81839f
C6118 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v49 GND 1.06253f
C6119 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v48 GND 1.66738f
C6120 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v39 GND 1.60815f
C6121 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v38 GND 1.05072f
C6122 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v37 GND 0.85279f
C6123 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v36 GND 0.85992f
C6124 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v35 GND 0.74171f
C6125 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v34 GND 0.83636f
C6126 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v33 GND 1.07608f
C6127 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v32 GND 1.72335f
C6128 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v23 GND 1.64361f
C6129 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v22 GND 1.10159f
C6130 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v21 GND 0.88377f
C6131 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v20 GND 0.90291f
C6132 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v19 GND 0.77336f
C6133 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v18 GND 0.88264f
C6134 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v17 GND 1.11637f
C6135 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v16 GND 1.84049f
C6136 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v7 GND 2.61761f
C6137 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v6 GND 1.84052f
C6138 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v5 GND 1.36319f
C6139 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v4 GND 1.54449f
C6140 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v3 GND 1.34744f
C6141 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v2 GND 2.56072f
C6142 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v1 GND 2.58685f
C6143 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 GND 1.486f
C6144 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 GND 0.92879f
C6145 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 GND 0.79566f
C6146 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 GND 0.8323f
C6147 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 GND 0.71956f
C6148 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 GND 0.79316f
C6149 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49 GND 0.97002f
C6150 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48 GND 1.65845f
C6151 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 GND 1.46001f
C6152 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 GND 0.87481f
C6153 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 GND 0.76797f
C6154 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 GND 0.79452f
C6155 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 GND 0.69232f
C6156 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 GND 0.75887f
C6157 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33 GND 0.94206f
C6158 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32 GND 1.57105f
C6159 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 GND 1.44143f
C6160 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 GND 0.85431f
C6161 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 GND 0.75086f
C6162 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 GND 0.77008f
C6163 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 GND 0.66926f
C6164 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 GND 0.73878f
C6165 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17 GND 0.92819f
C6166 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16 GND 1.52801f
C6167 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 GND 1.86046f
C6168 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 GND 0.84039f
C6169 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 GND 0.80384f
C6170 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 GND 0.77204f
C6171 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 GND 0.71421f
C6172 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 GND 0.72923f
C6173 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1 GND 0.95138f
C6174 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB GND 1.48613f
C6175 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN GND 1.2336f
C6176 a_43724_6956# GND 0.0275f
C6177 a_44234_6996# GND 0.94418f
C6178 a_44234_7352# GND 0.97967f
C6179 a_43724_7392# GND 0.02741f
C6180 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A GND 0.9729f
C6181 a_43698_6796# GND 0.37493f
C6182 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB GND 2.14419f
C6183 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN GND 1.66631f
C6184 a_43724_7946# GND 0.02732f
C6185 a_44234_7986# GND 0.97944f
C6186 a_44234_8342# GND 0.97944f
C6187 a_43724_8382# GND 0.02732f
C6188 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v63 GND 1.77222f
C6189 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v62 GND 1.00383f
C6190 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v61 GND 0.94283f
C6191 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v60 GND 0.92717f
C6192 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v59 GND 0.86196f
C6193 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v58 GND 1.47451f
C6194 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v57 GND 1.51886f
C6195 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v56 GND 2.59101f
C6196 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v47 GND 1.78935f
C6197 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v46 GND 0.999f
C6198 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v45 GND 0.9622f
C6199 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v44 GND 0.95203f
C6200 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v43 GND 0.93445f
C6201 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v42 GND 1.12363f
C6202 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v41 GND 1.58922f
C6203 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v40 GND 2.66791f
C6204 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v31 GND 1.77946f
C6205 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v30 GND 1.03387f
C6206 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v29 GND 0.98141f
C6207 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v28 GND 0.97038f
C6208 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v27 GND 0.95434f
C6209 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v26 GND 1.13854f
C6210 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v25 GND 1.60241f
C6211 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v24 GND 2.75231f
C6212 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v15 GND 1.8436f
C6213 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v14 GND 1.10941f
C6214 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v13 GND 1.06449f
C6215 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v12 GND 1.04526f
C6216 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v11 GND 1.05333f
C6217 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v10 GND 1.18974f
C6218 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v9 GND 1.70754f
C6219 top_DAC_0/top_rseg_n_dcell_0.top_segment_1_0.rseg_1_v3_1.v8 GND 3.4719f
C6220 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62 GND 1.65779f
C6221 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 GND 0.98593f
C6222 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 GND 0.96906f
C6223 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 GND 0.92766f
C6224 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 GND 1.4952f
C6225 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 GND 1.50125f
C6226 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 GND 2.51869f
C6227 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47 GND 1.53286f
C6228 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 GND 0.83546f
C6229 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 GND 0.83142f
C6230 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 GND 0.86302f
C6231 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 GND 0.8334f
C6232 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 GND 1.00167f
C6233 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 GND 1.4139f
C6234 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 GND 2.3234f
C6235 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31 GND 1.47968f
C6236 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 GND 0.79398f
C6237 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 GND 0.79447f
C6238 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 GND 0.8294f
C6239 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 GND 0.80491f
C6240 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 GND 0.96356f
C6241 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 GND 1.38045f
C6242 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 GND 2.26184f
C6243 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15 GND 1.45528f
C6244 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 GND 0.76536f
C6245 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 GND 0.79117f
C6246 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 GND 0.82395f
C6247 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 GND 0.79436f
C6248 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 GND 0.95967f
C6249 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 GND 1.37502f
C6250 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 GND 2.24954f
C6251 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A GND 0.77271f
C6252 a_43698_7786# GND 0.35068f
C6253 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB GND 1.38151f
C6254 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN GND 1.7426f
C6255 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] GND 3.54395f
C6256 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] GND 7.6635f
C6257 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] GND 3.69713f
C6258 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] GND 2.75844f
C6259 a_43724_8936# GND 0.02732f
C6260 a_44234_8976# GND 0.97944f
C6261 a_44234_9332# GND 0.97944f
C6262 a_43724_9372# GND 0.02732f
C6263 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A GND 0.76913f
C6264 a_31870_7686# GND 2.76379f
C6265 a_31594_7686# GND 1.42612f
C6266 a_31318_7686# GND 1.35431f
C6267 a_31042_7686# GND 1.27715f
C6268 a_30608_7686# GND 1.23382f
C6269 a_30332_7686# GND 1.1071f
C6270 a_30056_7686# GND 1.10378f
C6271 a_29780_7686# GND 1.83358f
C6272 a_29434_6250# GND 2.92347f
C6273 a_29158_6250# GND 1.51695f
C6274 a_28882_6250# GND 1.71491f
C6275 a_28606_6250# GND 1.98891f
C6276 a_28172_6250# GND 1.85978f
C6277 a_27896_6250# GND 1.46246f
C6278 a_27620_6250# GND 1.34968f
C6279 a_27344_6250# GND 2.32568f
C6280 a_17443_7686# GND 1.89753f
C6281 a_17167_7686# GND 0.90085f
C6282 a_16891_7686# GND 0.84018f
C6283 a_16615_7686# GND 0.8105f
C6284 a_16181_7686# GND 0.75573f
C6285 a_15905_7686# GND 0.63414f
C6286 a_15629_7686# GND 0.49296f
C6287 a_15353_7686# GND 0.6545f
C6288 a_15869_6250# GND 1.48025f
C6289 a_15593_6250# GND 0.80974f
C6290 a_15317_6250# GND 0.74476f
C6291 a_15041_6250# GND 1.03521f
C6292 a_14607_6250# GND 1.03185f
C6293 a_14331_6250# GND 0.67305f
C6294 a_14055_6250# GND 0.56947f
C6295 a_13779_6250# GND 0.69041f
C6296 a_43698_8776# GND 0.35068f
C6297 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB GND 1.70476f
C6298 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN GND 2.18999f
C6299 a_43724_9926# GND 0.02732f
C6300 a_44234_9966# GND 0.97944f
C6301 a_44234_10322# GND 0.97944f
C6302 a_43724_10362# GND 0.02732f
C6303 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A GND 0.77224f
C6304 a_35132_8950# GND 1.4146f
C6305 a_34856_8950# GND 0.75543f
C6306 a_34580_8950# GND 0.74455f
C6307 a_34304_8950# GND 0.80492f
C6308 a_34186_8950# GND 0.69668f
C6309 a_33910_8950# GND 0.71653f
C6310 a_33634_8950# GND 0.73252f
C6311 a_33358_8950# GND 1.17668f
C6312 a_36033_10031# GND 0.40395f
C6313 a_35757_10031# GND 0.39491f
C6314 a_35453_10031# GND 0.51368f
C6315 a_35177_10031# GND 1.20662f
C6316 a_34873_10031# GND 0.28185f
C6317 a_34569_10031# GND 0.39515f
C6318 a_20498_8950# GND 0.9473f
C6319 a_20222_8950# GND 0.41291f
C6320 a_19946_8950# GND 0.43734f
C6321 a_19670_8950# GND 0.40535f
C6322 a_19552_8950# GND 0.39876f
C6323 a_19276_8950# GND 0.38518f
C6324 a_19000_8950# GND 0.3768f
C6325 a_18724_8950# GND 0.5677f
C6326 a_20932_10031# GND 0.10857f
C6327 a_20656_10031# GND 0.17173f
C6328 a_20352_10031# GND 0.26688f
C6329 a_20076_10031# GND 0.84146f
C6330 a_19772_10031# GND 0.08053f
C6331 a_19468_10031# GND 0.21267f
C6332 a_43698_9766# GND 0.35068f
C6333 a_43724_10916# GND 0.02732f
C6334 a_44234_10956# GND 0.97944f
C6335 a_44234_11312# GND 0.97944f
C6336 a_43724_11352# GND 0.02732f
C6337 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP GND 0.72263f
C6338 a_43698_10756# GND 0.34573f
C6339 a_43724_11906# GND 0.02732f
C6340 a_44234_11946# GND 0.97944f
C6341 a_44234_12302# GND 0.97944f
C6342 a_43724_12342# GND 0.02732f
C6343 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP GND 0.71846f
C6344 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to2 GND 1.26949f
C6345 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to0 GND 0.80456f
C6346 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to1 GND 0.82997f
C6347 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to3 GND 2.03401f
C6348 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io1 GND 2.57321f
C6349 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.to4 GND 4.87217f
C6350 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.G1 GND 42.6114f
C6351 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_tail_0/cm_ncell1_0.io0 GND 8.66221f
C6352 a_5642_8388# GND 0.11496f $ **FLOATING
C6353 a_4978_8388# GND 0.10989f $ **FLOATING
C6354 a_5642_9535# GND 0.11145f $ **FLOATING
C6355 a_5111_8388# GND 0.63162f
C6356 a_4978_9535# GND 0.10301f $ **FLOATING
C6357 a_5642_10963# GND 0.35967f $ **FLOATING
C6358 a_4978_10963# GND 0.36693f $ **FLOATING
C6359 a_5642_11461# GND 0.38872f $ **FLOATING
C6360 a_5111_10963# GND 1.47391f
C6361 a_4978_11461# GND 0.34413f $ **FLOATING
C6362 a_2678_10356# GND 0.3141f $ **FLOATING
C6363 a_1896_10356# GND 0.31627f $ **FLOATING
C6364 a_2678_10974# GND 0.31147f $ **FLOATING
C6365 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.VTAIL2 GND 31.9875f
C6366 a_1896_10974# GND 0.31363f $ **FLOATING
C6367 a_43698_11746# GND 0.34573f
C6368 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN GND 1.76184f
C6369 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB GND 2.1668f
C6370 a_43724_12896# GND 0.02732f
C6371 a_44234_12936# GND 0.97944f
C6372 a_44234_13292# GND 0.97944f
C6373 a_43724_13332# GND 0.02732f
C6374 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP GND 0.71668f
C6375 a_43698_12736# GND 0.34573f
C6376 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB GND 2.03095f
C6377 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN GND 1.77046f
C6378 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN GND 1.69257f
C6379 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB GND 2.04707f
C6380 a_43724_13886# GND 0.02732f
C6381 a_44234_13926# GND 0.97944f
C6382 a_44234_14282# GND 0.97944f
C6383 a_43724_14322# GND 0.02732f
C6384 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP GND 0.71452f
C6385 a_43698_13726# GND 0.34573f
C6386 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN GND 1.95096f
C6387 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB GND 2.15197f
C6388 top_DAC_0/top_rseg_n_dcell_0.VS4 GND 1.44778f
C6389 top_DAC_0/top_rseg_n_dcell_0.SH[4] GND 2.30488f
C6390 top_DAC_0/top_rseg_n_dcell_0.SH[3] GND 2.30023f
C6391 a_15863_13287# GND 0.04049f
C6392 a_15863_13536# GND 0.01821f
C6393 a_15863_13785# GND 0.0393f
C6394 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb0 GND 3.66707f
C6395 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b0 GND 3.36789f
C6396 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb1 GND 4.43489f
C6397 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b1 GND 4.13168f
C6398 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb2 GND 5.96481f
C6399 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b2 GND 5.48635f
C6400 a_14615_13536# GND 0.1607f
C6401 a_14615_13785# GND 0.13123f
C6402 a_14615_14034# GND 0.12733f
C6403 a_14615_14283# GND 0.1775f
C6404 top_DAC_0/top_rseg_n_dcell_0.VS1 GND 6.64356f
C6405 top_DAC_0/top_rseg_n_dcell_0.SH[2] GND 3.55002f
C6406 top_DAC_0/top_rseg_n_dcell_0.SH[1] GND 6.74684f
C6407 a_12809_12507# GND 0.23775f $ **FLOATING
C6408 a_11629_12507# GND 0.2248f $ **FLOATING
C6409 a_12809_13005# GND 0.23111f $ **FLOATING
C6410 a_6923_9707# GND 4.02954f
C6411 a_11629_13005# GND 0.2208f $ **FLOATING
C6412 a_11081_12507# GND 0.22626f $ **FLOATING
C6413 a_9901_12507# GND 0.22553f $ **FLOATING
C6414 a_11081_13005# GND 0.2208f $ **FLOATING
C6415 a_8051_10107# GND 1.89392f
C6416 a_9901_13005# GND 0.2208f $ **FLOATING
C6417 a_9353_12507# GND 0.22485f $ **FLOATING
C6418 a_8173_12507# GND 0.22611f $ **FLOATING
C6419 a_9353_13005# GND 0.2208f $ **FLOATING
C6420 a_8506_12595# GND 1.10969f
C6421 a_8173_13005# GND 0.2208f $ **FLOATING
C6422 a_7625_12507# GND 0.22504f $ **FLOATING
C6423 a_6445_12507# GND 0.22721f $ **FLOATING
C6424 a_7625_13005# GND 0.2208f $ **FLOATING
C6425 a_6778_12595# GND 1.81371f
C6426 a_6445_13005# GND 0.2208f $ **FLOATING
C6427 a_5897_12507# GND 0.22396f $ **FLOATING
C6428 a_4717_12507# GND 0.23225f $ **FLOATING
C6429 a_5897_13005# GND 0.22049f $ **FLOATING
C6430 a_5050_12595# GND 2.14919f
C6431 a_4717_13005# GND 0.23057f $ **FLOATING
C6432 a_2678_11886# GND 0.31079f $ **FLOATING
C6433 a_1896_11886# GND 0.31296f $ **FLOATING
C6434 a_2678_12504# GND 0.31285f $ **FLOATING
C6435 a_1896_12504# GND 0.31297f $ **FLOATING
C6436 a_43724_14876# GND 0.02732f
C6437 a_44234_14916# GND 0.97944f
C6438 a_44234_15272# GND 0.97944f
C6439 a_43724_15312# GND 0.02732f
C6440 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP GND 0.71649f
C6441 a_43698_14716# GND 0.34573f
C6442 a_43724_15866# GND 0.02732f
C6443 a_44234_15906# GND 0.97944f
C6444 a_44234_16262# GND 0.98035f
C6445 a_43724_16302# GND 0.02747f
C6446 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP GND 0.71942f
C6447 a_12809_14150# GND 0.03735f $ **FLOATING
C6448 a_12809_15057# GND 0.03468f $ **FLOATING
C6449 top_DAC_0/top_final_switch_0.VOUT[4] GND 4.28985f
C6450 top_DAC_0/top_final_switch_0.VOUT[3] GND 3.40998f
C6451 top_DAC_0/top_final_switch_0.VOUT[2] GND 3.36007f
C6452 top_DAC_0/top_final_switch_0.VOUT[1] GND 3.35799f
C6453 a_4717_14150# GND 0.03708f $ **FLOATING
C6454 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPB GND 4.49065f
C6455 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_OPA GND 11.1641f
C6456 top_DAC_0/top_final_switch_0.VOUT[0] GND 4.35574f
C6457 a_4717_15057# GND 0.03501f $ **FLOATING
C6458 a_2300_13352# GND 0.27287f $ **FLOATING
C6459 a_1636_13352# GND 0.27787f $ **FLOATING
C6460 a_2300_13708# GND 0.26729f $ **FLOATING
C6461 a_1636_13708# GND 0.26729f $ **FLOATING
C6462 a_2300_14353# GND 0.06968f $ **FLOATING
C6463 a_1636_14353# GND 0.06968f $ **FLOATING
C6464 a_2300_15118# GND 0.06696f $ **FLOATING
C6465 a_1636_15118# GND 0.06696f $ **FLOATING
C6466 a_43698_15706# GND 0.34616f
C6467 a_43724_16856# GND 0.0277f
C6468 a_44234_16896# GND 0.98279f
C6469 a_44234_17252# GND 0.97824f
C6470 a_43724_17292# GND 0.02864f
C6471 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP GND 0.79071f
C6472 a_43698_16696# GND 0.53142f
C6473 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.79418f
C6474 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB GND 2.38299f
C6475 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.67704f
C6476 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB GND 2.84376f
C6477 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.643f
C6478 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN GND 2.08947f
C6479 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN GND 2.38321f
C6480 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.61395f
C6481 a_44062_18093# GND 0.73253f
C6482 a_44062_18449# GND 0.80123f
C6483 a_44062_18805# GND 0.76866f
C6484 a_44062_19161# GND 0.62805f
C6485 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.65617f
C6486 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] GND 3.84823f
C6487 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.67288f
C6488 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB GND 4.05136f
C6489 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.64256f
C6490 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] GND 4.00706f
C6491 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN GND 6.71896f
C6492 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.61568f
C6493 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC0 GND 6.16515f
C6494 a_24209_18133# GND 1.10636f
C6495 a_23629_18133# GND 0.97112f
C6496 a_23049_18133# GND 1.00054f
C6497 a_22469_18133# GND 1.20224f
C6498 top_DAC_0/top_rseg_n_dcell_0.VL2 GND 2.6263f
C6499 a_22193_18133# GND 2.35615f
C6500 top_DAC_0/top_rseg_n_dcell_0.VH2 GND 2.68525f
C6501 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[0] GND 12.8665f
C6502 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC1 GND 5.59751f
C6503 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[1] GND 11.5989f
C6504 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC2 GND 5.92507f
C6505 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[2] GND 9.96121f
C6506 top_DAC_0/top_rseg_n_dcell_0.VH3 GND 1.66107f
C6507 top_DAC_0/top_rseg_n_dcell_0.VL3 GND 1.80881f
C6508 a_18284_18696# GND 0.33888f
C6509 a_18008_18696# GND 0.19473f
C6510 a_17732_18696# GND 0.07551f
C6511 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.bb3 GND 10.0135f
C6512 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.b3 GND 9.70853f
C6513 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[4] GND 4.26794f
C6514 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[4] GND 2.70537f
C6515 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[5] GND 2.78919f
C6516 a_15618_18696# GND 0.61717f
C6517 a_15342_18696# GND 0.34164f
C6518 a_15066_18696# GND 0.37474f
C6519 a_14790_18696# GND 0.25093f
C6520 a_14514_18696# GND 0.15715f
C6521 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[5] GND 4.27305f
C6522 a_44062_19517# GND 0.62696f
C6523 a_44062_19873# GND 0.79679f
C6524 a_44062_20229# GND 0.76698f
C6525 a_44062_20585# GND 0.62705f
C6526 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.DEC3 GND 6.35874f
C6527 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC2[3] GND 11.4627f
C6528 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[3] GND 4.8343f
C6529 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.61845f
C6530 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] GND 3.5102f
C6531 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.66383f
C6532 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] GND 2.31971f
C6533 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.63305f
C6534 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] GND 2.72833f
C6535 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] GND 5.39912f
C6536 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.75299f
C6537 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[2] GND 4.41444f
C6538 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[1] GND 4.67667f
C6539 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC1[0] GND 4.59773f
C6540 a_44062_20941# GND 0.62696f
C6541 a_44062_21297# GND 0.79679f
C6542 a_44062_21653# GND 0.76698f
C6543 a_44062_22009# GND 0.71256f
C6544 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] GND 6.91015f
C6545 a_39883_19098# GND 0.21843f $ **FLOATING
C6546 a_37277_19098# GND 0.24267f $ **FLOATING
C6547 a_39883_19479# GND 0.20382f $ **FLOATING
C6548 a_37737_19479# GND 0.18912f $ **FLOATING
C6549 a_39883_19854# GND 0.20634f $ **FLOATING
C6550 a_38617_19854# GND 0.21532f $ **FLOATING
C6551 a_37595_19462# GND 0.15668f $ **FLOATING
C6552 a_36813_19462# GND 0.19962f $ **FLOATING
C6553 a_37595_19760# GND 0.19172f $ **FLOATING
C6554 a_36813_19760# GND 0.19708f $ **FLOATING
C6555 a_39768_20389# GND 0.17117f $ **FLOATING
C6556 a_38584_20389# GND 0.17006f $ **FLOATING
C6557 a_39768_20665# GND 0.17317f $ **FLOATING
C6558 a_38672_20477# GND 1.01366f
C6559 a_39306_20477# GND 0.4451f
C6560 a_37410_19098# GND 7.09932f
C6561 a_38584_20665# GND 0.17331f $ **FLOATING
C6562 a_37804_20295# GND 0.18145f $ **FLOATING
C6563 a_37022_20295# GND 0.17721f $ **FLOATING
C6564 a_37804_20713# GND 0.18276f $ **FLOATING
C6565 a_36888_19550# GND 1.43258f
C6566 a_36888_19786# GND 4.34674f
C6567 a_37022_20713# GND 0.17864f $ **FLOATING
C6568 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_5.I_HEAD GND 0.77724f
C6569 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_2.I_HEAD GND 0.8348f
C6570 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_3.I_HEAD GND 0.75334f
C6571 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_1.I_HEAD GND 1.06939f
C6572 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB2 GND 4.66799f
C6573 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_pmos_top_0/dp_pmos_0.I_HEAD GND 1.34759f
C6574 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_ncell3_0.DRAIN GND 44.3864f
C6575 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[0] GND 9.39959f
C6576 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[1] GND 8.68998f
C6577 a_24963_20174# GND 1.82982f
C6578 a_24687_20174# GND 1.24913f
C6579 a_24411_20174# GND 1.23985f
C6580 a_24135_20174# GND 1.07549f
C6581 a_23859_20174# GND 1.53863f
C6582 a_23583_20174# GND 1.0992f
C6583 a_23307_20174# GND 1.54243f
C6584 a_23031_20174# GND 1.32237f
C6585 a_22755_20174# GND 1.62006f
C6586 a_22479_20174# GND 1.38915f
C6587 a_22203_20174# GND 1.48313f
C6588 a_21927_20174# GND 1.63658f
C6589 a_21651_20174# GND 1.62945f
C6590 a_21375_20174# GND 2.27588f
C6591 a_21099_20174# GND 1.59228f
C6592 a_20823_20174# GND 1.67062f
C6593 a_20547_20174# GND 1.94548f
C6594 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.DEC0[2] GND 9.29455f
C6595 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.bb[6] GND 4.36453f
C6596 a_17148_18696# GND 0.26539f
C6597 a_16872_18696# GND 0.26002f
C6598 a_16596_18696# GND 0.29086f
C6599 a_16320_18696# GND 0.31116f
C6600 a_14672_18696# GND 0.54051f
C6601 a_14948_18696# GND 0.36296f
C6602 a_15224_18696# GND 0.35512f
C6603 a_15374_19866# GND 0.31759f
C6604 a_15098_19866# GND 0.31904f
C6605 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.b[6] GND 3.89091f
C6606 a_40525_21457# GND 0.05335f $ **FLOATING
C6607 a_39861_21457# GND 0.01074f $ **FLOATING
C6608 a_41907_22057# GND 0.01121f $ **FLOATING
C6609 a_39936_22083# GND 0.1294f
C6610 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV GND 9.50443f
C6611 a_44067_22496# GND 0.18164f $ **FLOATING
C6612 a_43994_22522# GND 0.39309f
C6613 a_39861_22496# GND 0.0387f $ **FLOATING
C6614 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV GND 19.1265f
C6615 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1 GND 2.4989f
C6616 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC GND 4.4367f
C6617 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC GND 11.6586f
C6618 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0 GND 2.18342f
C6619 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 GND 0.25356f
C6620 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 GND 0.27668f
C6621 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 GND 0.2878f
C6622 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 GND 0.34405f
C6623 top_DAC_0/top_rseg_n_dcell_0.top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 GND 1.98271f
C6624 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.V0 GND 9.78667f
C6625 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v16 GND 3.07483f
C6626 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v32 GND 3.01107f
C6627 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v1 GND 2.06217f
C6628 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v15 GND 1.52657f
C6629 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v17 GND 1.48589f
C6630 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v31 GND 1.48556f
C6631 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v33 GND 1.48168f
C6632 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v47 GND 1.55719f
C6633 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v2 GND 1.12435f
C6634 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v14 GND 0.82563f
C6635 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v18 GND 0.84609f
C6636 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v30 GND 0.80858f
C6637 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v34 GND 0.82727f
C6638 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v46 GND 0.91672f
C6639 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v3 GND 1.25062f
C6640 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v13 GND 0.85946f
C6641 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v19 GND 0.8303f
C6642 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v29 GND 0.83077f
C6643 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v35 GND 0.82365f
C6644 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v45 GND 0.89932f
C6645 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v4 GND 1.20222f
C6646 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v12 GND 0.89682f
C6647 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v20 GND 0.9106f
C6648 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v28 GND 0.87434f
C6649 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v36 GND 0.88241f
C6650 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v44 GND 1.00071f
C6651 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v5 GND 1.32479f
C6652 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v11 GND 0.93857f
C6653 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v21 GND 0.8879f
C6654 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v27 GND 0.88592f
C6655 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v37 GND 0.87598f
C6656 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v43 GND 0.96048f
C6657 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v6 GND 1.25445f
C6658 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v10 GND 0.96146f
C6659 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v22 GND 0.98448f
C6660 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v26 GND 0.9598f
C6661 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v38 GND 0.92655f
C6662 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v42 GND 1.58503f
C6663 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v7 GND 2.65934f
C6664 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v9 GND 1.38005f
C6665 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v8 GND 2.71993f
C6666 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v23 GND 1.45804f
C6667 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v25 GND 1.37054f
C6668 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v24 GND 2.32676f
C6669 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v39 GND 1.45618f
C6670 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v41 GND 1.48352f
C6671 top_DAC_0/top_rseg_n_dcell_0.top_segment_2_0.rseg_2_v3_0.v40 GND 2.34388f
C6672 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.V0 GND 2.93398f
C6673 top_DAC_0/top_rseg_n_dcell_0.top_segment_4_1.V0 GND 8.59418f
C6674 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v1 GND 1.10729f
C6675 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v15 GND 1.3484f
C6676 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v2 GND 0.9104f
C6677 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v14 GND 1.20251f
C6678 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v3 GND 0.85989f
C6679 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v13 GND 1.06531f
C6680 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v4 GND 0.94f
C6681 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v12 GND 1.23818f
C6682 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v5 GND 0.93563f
C6683 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v11 GND 1.01098f
C6684 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v6 GND 1.09411f
C6685 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v10 GND 1.50562f
C6686 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v7 GND 2.01393f
C6687 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v9 GND 1.54963f
C6688 top_DAC_0/top_rseg_n_dcell_0.top_segment_3_0.rseg_3_v3_0.v8 GND 3.06885f
C6689 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho0 GND 0.22202f
C6690 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho1 GND 0.2191f
C6691 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho2 GND 0.3605f
C6692 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho3 GND 0.62827f
C6693 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io2 GND 0.69908f
C6694 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.ho4 GND 1.27694f
C6695 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io0 GND 1.51612f
C6696 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.io1 GND 1.4754f
C6697 a_2678_16243# GND 0.03553f $ **FLOATING
C6698 a_1896_16243# GND 0.04167f $ **FLOATING
C6699 a_2678_17510# GND 0.03283f $ **FLOATING
C6700 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.B GND 5.42729f
C6701 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Bx GND 10.3408f
C6702 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.VB1 GND 5.60786f
C6703 a_1896_17510# GND 0.04167f $ **FLOATING
C6704 a_2678_19053# GND 0.03256f $ **FLOATING
C6705 a_1896_19053# GND 0.04167f $ **FLOATING
C6706 a_2678_20320# GND 0.03256f $ **FLOATING
C6707 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.A GND 2.10155f
C6708 a_1896_20320# GND 0.04167f $ **FLOATING
C6709 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/cm_pcell3_0.VB2 GND 16.0806f
C6710 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/cm_head_0/cm_pcell1_0.G1 GND 15.7829f
C6711 a_4415_23194# GND 12.5641f
C6712 a_8473_23194# GND 0.43004f
C6713 a_2678_21703# GND 0.03256f $ **FLOATING
C6714 a_1896_21703# GND 0.04167f $ **FLOATING
C6715 a_2678_22970# GND 0.03813f $ **FLOATING
C6716 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONB GND 3.47647f
C6717 top_DAC_0/top_buffer_opamp_0.opa_input_and_self_bias_0/opa_input_stage_0/opa_diffpairs_0/dp_nmos_top_0/dp_nmos_5.I_ONA GND 8.72764f
C6718 top_DAC_0/top_buffer_opamp_0.opa_folded_cascode_0.monticelli_top_0.Ax GND 2.16756f
C6719 a_1896_22970# GND 0.04724f $ **FLOATING
.ends

