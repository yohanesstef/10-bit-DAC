magic
tech sky130A
magscale 1 2
timestamp 1749375316
<< metal1 >>
rect 89 3571 149 3577
rect 89 2955 149 3511
rect 177 3395 237 3401
rect 177 2955 237 3335
rect 265 3219 325 3225
rect 265 2955 325 3159
rect 441 3131 501 3659
rect 441 3065 501 3071
rect 529 2955 589 3659
rect 617 3131 677 3659
rect 705 3219 765 3659
rect 793 3307 853 3659
rect 881 3395 941 3659
rect 969 3483 1029 3659
rect 1057 3571 1117 3659
rect 1057 3505 1117 3511
rect 969 3417 1029 3423
rect 881 3329 941 3335
rect 793 3241 853 3247
rect 705 3153 765 3159
rect 617 3065 677 3071
<< via1 >>
rect 89 3511 149 3571
rect 177 3335 237 3395
rect 265 3159 325 3219
rect 441 3071 501 3131
rect 1057 3511 1117 3571
rect 969 3423 1029 3483
rect 881 3335 941 3395
rect 793 3247 853 3307
rect 705 3159 765 3219
rect 617 3071 677 3131
<< metal2 >>
rect 83 3511 89 3571
rect 149 3511 1057 3571
rect 1117 3511 1123 3571
rect 963 3423 969 3483
rect 1029 3423 1221 3483
rect 171 3335 177 3395
rect 237 3335 881 3395
rect 941 3335 947 3395
rect 787 3247 793 3307
rect 853 3247 1221 3307
rect 259 3159 265 3219
rect 325 3159 705 3219
rect 765 3159 771 3219
rect 435 3071 441 3131
rect 501 3071 507 3131
rect 611 3071 617 3131
rect 677 3071 1221 3131
rect 441 2955 501 3071
<< end >>
