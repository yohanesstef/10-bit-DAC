magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -653 307 653
<< psubdiff >>
rect -271 583 -175 617
rect 175 583 271 617
rect -271 521 -237 583
rect 237 521 271 583
rect -271 -583 -237 -521
rect 237 -583 271 -521
rect -271 -617 -175 -583
rect 175 -617 271 -583
<< psubdiffcont >>
rect -175 583 175 617
rect -271 -521 -237 521
rect 237 -521 271 521
rect -175 -617 175 -583
<< xpolycontact >>
rect -141 55 141 487
rect -141 -487 141 -55
<< xpolyres >>
rect -141 -55 141 55
<< locali >>
rect -271 583 -175 617
rect 175 583 271 617
rect -271 521 -237 583
rect 237 521 271 583
rect -271 -583 -237 -521
rect 237 -583 271 -521
rect -271 -617 -175 -583
rect 175 -617 271 -583
<< viali >>
rect -125 72 125 469
rect -125 -469 125 -72
<< metal1 >>
rect -131 469 131 481
rect -131 72 -125 469
rect 125 72 131 469
rect -131 60 131 72
rect -131 -72 131 -60
rect -131 -469 -125 -72
rect 125 -469 131 -72
rect -131 -481 131 -469
<< properties >>
string FIXED_BBOX -254 -600 254 600
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 0.707 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 1.269k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
