magic
tech sky130A
magscale 1 2
timestamp 1749664768
<< locali >>
rect 35102 -5170 35136 -4445
rect 39256 -5170 39290 -4445
rect 36750 -5204 39063 -5170
rect 36716 -5588 36750 -5526
rect 39063 -5588 39097 -5526
rect 36716 -5622 39097 -5588
rect 34358 -6506 34392 -5622
rect 36716 -6506 36750 -5622
rect 33441 -6540 34579 -6506
rect 36555 -6540 37693 -6506
rect 39063 -6540 39097 -5622
rect 39740 -6540 40878 -6506
rect 41421 -6540 41455 -5526
rect 37443 -6924 37477 -6862
rect 39801 -6924 39835 -6862
rect 40781 -6924 40815 -6862
rect 33441 -6958 34579 -6924
rect 36555 -6958 37693 -6924
rect 39801 -6958 40815 -6924
rect 31145 -7870 31179 -6958
rect 33503 -7870 33537 -6958
rect 34259 -7870 34293 -6958
rect 31963 -7904 32653 -7870
rect 35045 -7904 35802 -7870
rect 36617 -7879 36651 -6958
rect 37443 -7879 37477 -6958
rect 38194 -7904 39063 -7870
rect 39801 -7879 39835 -6958
rect 40781 -7879 40815 -6958
rect 31963 -8322 32653 -8288
rect 35045 -8322 35802 -8288
rect 38194 -8322 39063 -8288
rect 29921 -8684 29942 -8680
<< metal1 >>
rect 33687 -5474 34291 -5414
rect 36817 -5474 37160 -5414
rect 30737 -6768 30797 -6762
rect 30737 -7992 30797 -6828
rect 33687 -7824 33747 -5474
rect 33775 -5562 34291 -5502
rect 36817 -5562 37072 -5502
rect 33775 -7736 33835 -5562
rect 33863 -5650 34291 -5590
rect 36817 -5650 36984 -5590
rect 33863 -7648 33923 -5650
rect 33951 -5738 34291 -5678
rect 36817 -5738 36896 -5678
rect 33951 -7560 34011 -5738
rect 33951 -7626 34011 -7620
rect 33863 -7714 33923 -7708
rect 33775 -7802 33835 -7796
rect 33687 -7890 33747 -7884
rect 34475 -8052 34535 -6775
rect 36836 -7472 36896 -5738
rect 36924 -7384 36984 -5650
rect 37012 -7296 37072 -5562
rect 37100 -7208 37160 -5474
rect 39921 -6470 39981 -5758
rect 40009 -6382 40069 -5764
rect 40097 -6294 40157 -5764
rect 40185 -6206 40245 -5764
rect 40273 -6118 40333 -5764
rect 40361 -6030 40421 -5764
rect 40449 -5942 40509 -5764
rect 40537 -5854 40597 -5764
rect 40537 -5920 40597 -5914
rect 40449 -6008 40509 -6002
rect 40361 -6096 40421 -6090
rect 40273 -6184 40333 -6178
rect 40185 -6272 40245 -6266
rect 40097 -6360 40157 -6354
rect 40009 -6448 40069 -6442
rect 39921 -6536 39981 -6530
rect 40229 -6768 40289 -6762
rect 37100 -7274 37160 -7268
rect 37012 -7362 37072 -7356
rect 36924 -7450 36984 -7444
rect 36836 -7538 36896 -7532
rect 37634 -8052 37694 -6775
rect 40229 -7992 40289 -6828
rect 30737 -8058 30797 -8052
rect 40229 -8058 40289 -8052
<< via1 >>
rect 30737 -6828 30797 -6768
rect 33951 -7620 34011 -7560
rect 33863 -7708 33923 -7648
rect 33775 -7796 33835 -7736
rect 33687 -7884 33747 -7824
rect 30737 -8052 30797 -7992
rect 40537 -5914 40597 -5854
rect 40449 -6002 40509 -5942
rect 40361 -6090 40421 -6030
rect 40273 -6178 40333 -6118
rect 40185 -6266 40245 -6206
rect 40097 -6354 40157 -6294
rect 40009 -6442 40069 -6382
rect 39921 -6530 39981 -6470
rect 37100 -7268 37160 -7208
rect 37012 -7356 37072 -7296
rect 36924 -7444 36984 -7384
rect 36836 -7532 36896 -7472
rect 40229 -6828 40289 -6768
rect 40229 -8052 40289 -7992
<< metal2 >>
rect 36380 -4568 41365 -4508
rect 36104 -4656 41089 -4596
rect 35828 -4744 40813 -4684
rect 35562 -4832 40537 -4772
rect 35474 -4920 40053 -4860
rect 35208 -5008 39777 -4948
rect 34932 -5096 39501 -5036
rect 34656 -5184 39225 -5124
rect 33350 -5914 40537 -5854
rect 40597 -5914 43058 -5854
rect 33074 -6002 40449 -5942
rect 40509 -6002 42782 -5942
rect 32798 -6090 40361 -6030
rect 40421 -6090 42506 -6030
rect 32522 -6178 40273 -6118
rect 40333 -6178 42230 -6118
rect 32088 -6266 40185 -6206
rect 40245 -6266 41796 -6206
rect 31812 -6354 40097 -6294
rect 40157 -6354 41520 -6294
rect 31536 -6442 40009 -6382
rect 40069 -6442 41244 -6382
rect 31260 -6530 39921 -6470
rect 39981 -6530 40968 -6470
rect 30731 -6828 30737 -6768
rect 30797 -6828 31325 -6768
rect 40223 -6828 40229 -6768
rect 40289 -6828 40961 -6768
rect 31801 -7268 37100 -7208
rect 37160 -7268 41365 -7208
rect 31525 -7356 37012 -7296
rect 37072 -7356 41089 -7296
rect 31249 -7444 36924 -7384
rect 36984 -7444 40813 -7384
rect 30973 -7532 36836 -7472
rect 36896 -7532 40537 -7472
rect 30489 -7620 33951 -7560
rect 34011 -7620 40053 -7560
rect 30213 -7708 33863 -7648
rect 33923 -7708 39777 -7648
rect 29937 -7796 33775 -7736
rect 33835 -7796 39501 -7736
rect 29661 -7884 33687 -7824
rect 33747 -7884 39225 -7824
rect 30731 -8000 30737 -7992
rect 30797 -8000 30803 -7992
rect 40223 -8000 40229 -7992
rect 40289 -8000 40295 -7992
rect 29885 -9174 29906 -9170
rect 43301 -9174 43322 -9170
use pgring_16  pgring_16_0
timestamp 1749664768
transform 1 0 -2162 0 1 -438
box 37186 -4752 41530 -3335
use pswitch_8_stage_1  pswitch_8_stage_1_0
timestamp 1749415301
transform 1 0 0 0 1 0
box 29493 -8466 32041 -7202
use pswitch_8_stage_1  pswitch_8_stage_1_1
timestamp 1749415301
transform 1 0 3082 0 1 0
box 29493 -8466 32041 -7202
use pswitch_8_stage_1  pswitch_8_stage_1_2
timestamp 1749415301
transform 1 0 6231 0 1 0
box 29493 -8466 32041 -7202
use pswitch_8_stage_1  pswitch_8_stage_1_3
timestamp 1749415301
transform 1 0 9492 0 1 0
box 29493 -8466 32041 -7202
use pswitch_8_stage_1  pswitch_8_stage_1_4
timestamp 1749415301
transform 1 0 9492 0 1 2700
box 29493 -8466 32041 -7202
use pswitch_8_stage_1_up  pswitch_8_stage_1_up_0
timestamp 1749415301
transform 1 0 1574 0 1 1346
box 29493 -9812 32041 -7194
use pswitch_8_stage_1_up  pswitch_8_stage_1_up_1
timestamp 1749415301
transform 1 0 4688 0 1 1346
box 29493 -9812 32041 -7194
use pswitch_8_stage_1_up  pswitch_8_stage_1_up_2
timestamp 1749415301
transform 1 0 7872 0 1 1346
box 29493 -9812 32041 -7194
use pswitch_8_stage_1_up  pswitch_8_stage_1_up_3
timestamp 1749415301
transform 1 0 11210 0 1 1346
box 29493 -9812 32041 -7194
use pswitch_8_stage_2  pswitch_8_stage_2_0
timestamp 1749415301
transform 1 0 0 0 1 -88
box 34280 -5650 36828 -4414
use rseg_4_routing  rseg_4_routing_0
timestamp 1749465145
transform 1 0 29988 0 1 -12125
box -103 -101 13334 3659
<< labels >>
flabel metal2 s 29885 -9170 29885 -9170 4 FreeSans 1600 0 0 0 V0
port 0 se
flabel metal2 s 43322 -9170 43322 -9170 6 FreeSans 1600 0 0 0 V63
port 1 sw
flabel metal1 s 30737 -6762 30737 -6762 4 FreeSans 800 0 0 0 DEC0
port 2 se
flabel metal1 s 34475 -7126 34475 -7126 4 FreeSans 800 0 0 0 DEC1
port 3 se
flabel metal1 s 37634 -7117 37634 -7117 4 FreeSans 800 0 0 0 DEC2
port 4 se
flabel metal1 s 40229 -7069 40229 -7069 4 FreeSans 800 0 0 0 DEC3
port 5 se
flabel metal2 s 35498 -4219 35498 -4219 4 FreeSans 480 0 0 0 b0
port 6 se
flabel metal2 s 35194 -4219 35194 -4219 4 FreeSans 480 0 0 0 bb0
port 10 se
flabel metal2 s 35192 -4043 35192 -4043 4 FreeSans 480 0 0 0 VOUT
port 14 se
flabel locali s 29921 -8680 29921 -8680 4 FreeSans 1600 0 0 0 GND
port 15 se
flabel metal2 s 38115 -4246 38115 -4246 4 FreeSans 480 0 0 0 bb2
port 12 se
flabel metal2 s 38003 -4244 38003 -4244 4 FreeSans 480 0 0 0 b2
port 8 se
flabel locali s 31161 -7270 31161 -7270 2 FreeSans 1600 0 0 0 VPB
port 16 ne
flabel metal2 s 39171 -5319 39171 -5319 4 FreeSans 480 0 0 0 bb3
port 13 se
flabel metal2 s 36614 -5332 36614 -5332 4 FreeSans 480 0 0 0 b3
port 9 se
flabel metal2 s 36285 -4253 36285 -4253 4 FreeSans 480 0 0 0 bb1
port 11 se
flabel metal2 s 36431 -4250 36431 -4250 4 FreeSans 480 0 0 0 b1
port 7 se
<< end >>
