magic
tech sky130A
magscale 1 2
timestamp 1749147130
<< pwell >>
rect -307 -755 307 755
<< psubdiff >>
rect -271 685 -175 719
rect 175 685 271 719
rect -271 623 -237 685
rect 237 623 271 685
rect -271 -685 -237 -623
rect 237 -685 271 -623
rect -271 -719 -175 -685
rect 175 -719 271 -685
<< psubdiffcont >>
rect -175 685 175 719
rect -271 -623 -237 623
rect 237 -623 271 623
rect -175 -719 175 -685
<< xpolycontact >>
rect -141 157 141 589
rect -141 -589 141 -157
<< xpolyres >>
rect -141 -157 141 157
<< locali >>
rect -271 685 -175 719
rect 175 685 271 719
rect -271 623 -237 685
rect 237 623 271 685
rect -271 -685 -237 -623
rect 237 -685 271 -623
rect -271 -719 -175 -685
rect 175 -719 271 -685
<< viali >>
rect -125 174 125 571
rect -125 -571 125 -174
<< metal1 >>
rect -131 571 131 583
rect -131 174 -125 571
rect 125 174 131 571
rect -131 162 131 174
rect -131 -174 131 -162
rect -131 -571 -125 -174
rect 125 -571 131 -174
rect -131 -583 131 -571
<< properties >>
string FIXED_BBOX -254 -702 254 702
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.733 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 2.725k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
