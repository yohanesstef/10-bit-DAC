magic
tech sky130A
magscale 1 2
timestamp 1750204660
<< nwell >>
rect -392 407 2922 534
rect -1876 -756 2922 407
rect -392 -866 2922 -756
<< mvnsubdiff >>
rect -1440 166 -574 226
rect -1440 -431 -1380 166
rect -634 -431 -574 166
rect -1440 -491 -574 -431
rect -273 -36 1975 24
rect -273 -415 -213 -36
rect 1915 -415 1975 -36
rect -273 -475 1975 -415
<< poly >>
rect -1369 -345 -1309 138
rect -705 -345 -645 138
rect -202 -387 -142 -64
rect 1844 -387 1904 -64
<< locali >>
rect -1427 179 -587 213
rect -1427 -444 -1393 179
rect -621 -444 -587 179
rect -1427 -478 -587 -444
rect -260 -23 1962 11
rect -260 -428 -226 -23
rect 1928 -428 1962 -23
rect -260 -462 1962 -428
<< metal1 >>
rect -1450 156 -564 236
rect -1450 -421 -1370 156
rect -1061 82 -953 128
rect -1288 -347 -1242 -319
rect -772 -347 -726 -319
rect -1288 -393 -726 -347
rect -644 -421 -564 156
rect -1450 -501 -564 -421
rect -283 -46 1985 34
rect -283 -405 -203 -46
rect 1905 -405 1985 -46
rect -283 -485 1985 -405
use sky130_fd_pr__pfet_g5v0d10v5_NWEVUG  sky130_fd_pr__pfet_g5v0d10v5_NWEVUG_0
timestamp 1750204660
transform 1 0 851 0 1 -225
box -1044 -202 1044 164
use sky130_fd_pr__pfet_g5v0d10v5_YDEY4G  sky130_fd_pr__pfet_g5v0d10v5_YDEY4G_0
timestamp 1750203654
transform 1 0 -1007 0 1 -103
box -353 -282 353 244
<< end >>
