magic
tech sky130A
magscale 1 2
timestamp 1750150351
<< nwell >>
rect 2267 -1100 3957 1902
<< mvnsubdiffcont >>
rect 2406 1789 3818 1823
rect 2346 -961 2380 1763
rect 3844 -961 3878 1763
rect 2406 -1021 3818 -987
<< metal1 >>
rect 2669 1682 2675 1742
rect 3135 1682 3141 1742
rect 3201 1682 3207 1742
rect 3030 1654 3076 1682
rect 3017 1594 3023 1654
rect 3083 1594 3089 1654
rect 3148 1603 3194 1682
rect 2772 491 2818 519
rect 3406 491 3452 519
rect 2772 431 2938 491
rect 3227 431 3386 491
rect 3446 431 3452 491
rect 3561 371 3621 1748
rect 2772 311 2938 371
rect 3227 311 3621 371
rect 2772 283 2818 311
rect 3406 283 3452 311
rect 3148 -792 3194 -787
rect 3030 -880 3076 -796
rect 3135 -852 3141 -792
rect 3201 -852 3207 -792
rect 3017 -940 3023 -880
rect 3083 -940 3089 -880
rect 3148 -940 3194 -852
rect 3561 -946 3621 311
rect 3649 491 3709 497
rect 3649 -946 3709 431
<< via1 >>
rect 2609 1682 2669 1742
rect 3141 1682 3201 1742
rect 2515 1594 2575 1654
rect 3023 1594 3083 1654
rect 3386 431 3446 491
rect 2515 -852 2575 -792
rect 3141 -852 3201 -792
rect 2603 -940 2663 -880
rect 3023 -940 3083 -880
rect 3649 431 3709 491
<< metal2 >>
rect 2603 1682 2609 1742
rect 2669 1682 2707 1742
rect 2509 1594 2515 1654
rect 2575 1594 3023 1654
rect 3380 431 3386 491
rect 3446 431 3649 491
rect 3709 431 3715 491
rect 2509 -852 2515 -792
rect 2575 -852 2684 -792
rect 2509 -940 2603 -880
rect 2663 -940 2684 -880
use cross_pair  cross_pair_0
timestamp 1750150351
transform 1 0 -33176 0 1 -1544
box 36114 1855 36403 2035
use fc_pmos2_2  fc_pmos2_2_0
timestamp 1750012037
transform 1 0 2707 0 1 463
box -440 -128 1250 1439
use fc_pmos2_2  fc_pmos2_2_1
timestamp 1750012037
transform 1 0 2707 0 -1 339
box -440 -128 1250 1439
<< end >>
