magic
tech sky130A
magscale 1 2
timestamp 1750900893
use hnmos_1  hnmos_1_0
timestamp 1750900893
transform 1 0 37 0 1 -2
box -41 3 235 201
use hnmos_1  hnmos_1_1
timestamp 1750900893
transform 1 0 313 0 1 -2
box -41 3 235 201
<< end >>
