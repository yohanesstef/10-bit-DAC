magic
tech sky130A
magscale 1 2
timestamp 1750845293
<< metal1 >>
rect 197 250 225 1250
rect 285 212 313 1172
use sky130_fd_pr__nfet_g5v0d10v5_ZUVY8G  sky130_fd_pr__nfet_g5v0d10v5_ZUVY8G_0
timestamp 1750845293
transform 1 0 211 0 1 681
box -278 -749 278 749
<< labels >>
flabel metal1 s 211 328 211 328 0 FreeSans 320 0 0 0 DIN
port 0 nsew
flabel metal1 s 296 722 296 722 0 FreeSans 320 0 0 0 VIN
port 1 nsew
<< end >>
