magic
tech sky130A
magscale 1 2
timestamp 1750148716
<< metal3 >>
rect -3422 2012 -2650 2040
rect -3422 1588 -2734 2012
rect -2670 1588 -2650 2012
rect -3422 1560 -2650 1588
rect -2410 2012 -1638 2040
rect -2410 1588 -1722 2012
rect -1658 1588 -1638 2012
rect -2410 1560 -1638 1588
rect -1398 2012 -626 2040
rect -1398 1588 -710 2012
rect -646 1588 -626 2012
rect -1398 1560 -626 1588
rect -386 2012 386 2040
rect -386 1588 302 2012
rect 366 1588 386 2012
rect -386 1560 386 1588
rect 626 2012 1398 2040
rect 626 1588 1314 2012
rect 1378 1588 1398 2012
rect 626 1560 1398 1588
rect 1638 2012 2410 2040
rect 1638 1588 2326 2012
rect 2390 1588 2410 2012
rect 1638 1560 2410 1588
rect 2650 2012 3422 2040
rect 2650 1588 3338 2012
rect 3402 1588 3422 2012
rect 2650 1560 3422 1588
rect -3422 1292 -2650 1320
rect -3422 868 -2734 1292
rect -2670 868 -2650 1292
rect -3422 840 -2650 868
rect -2410 1292 -1638 1320
rect -2410 868 -1722 1292
rect -1658 868 -1638 1292
rect -2410 840 -1638 868
rect -1398 1292 -626 1320
rect -1398 868 -710 1292
rect -646 868 -626 1292
rect -1398 840 -626 868
rect -386 1292 386 1320
rect -386 868 302 1292
rect 366 868 386 1292
rect -386 840 386 868
rect 626 1292 1398 1320
rect 626 868 1314 1292
rect 1378 868 1398 1292
rect 626 840 1398 868
rect 1638 1292 2410 1320
rect 1638 868 2326 1292
rect 2390 868 2410 1292
rect 1638 840 2410 868
rect 2650 1292 3422 1320
rect 2650 868 3338 1292
rect 3402 868 3422 1292
rect 2650 840 3422 868
rect -3422 572 -2650 600
rect -3422 148 -2734 572
rect -2670 148 -2650 572
rect -3422 120 -2650 148
rect -2410 572 -1638 600
rect -2410 148 -1722 572
rect -1658 148 -1638 572
rect -2410 120 -1638 148
rect -1398 572 -626 600
rect -1398 148 -710 572
rect -646 148 -626 572
rect -1398 120 -626 148
rect -386 572 386 600
rect -386 148 302 572
rect 366 148 386 572
rect -386 120 386 148
rect 626 572 1398 600
rect 626 148 1314 572
rect 1378 148 1398 572
rect 626 120 1398 148
rect 1638 572 2410 600
rect 1638 148 2326 572
rect 2390 148 2410 572
rect 1638 120 2410 148
rect 2650 572 3422 600
rect 2650 148 3338 572
rect 3402 148 3422 572
rect 2650 120 3422 148
rect -3422 -148 -2650 -120
rect -3422 -572 -2734 -148
rect -2670 -572 -2650 -148
rect -3422 -600 -2650 -572
rect -2410 -148 -1638 -120
rect -2410 -572 -1722 -148
rect -1658 -572 -1638 -148
rect -2410 -600 -1638 -572
rect -1398 -148 -626 -120
rect -1398 -572 -710 -148
rect -646 -572 -626 -148
rect -1398 -600 -626 -572
rect -386 -148 386 -120
rect -386 -572 302 -148
rect 366 -572 386 -148
rect -386 -600 386 -572
rect 626 -148 1398 -120
rect 626 -572 1314 -148
rect 1378 -572 1398 -148
rect 626 -600 1398 -572
rect 1638 -148 2410 -120
rect 1638 -572 2326 -148
rect 2390 -572 2410 -148
rect 1638 -600 2410 -572
rect 2650 -148 3422 -120
rect 2650 -572 3338 -148
rect 3402 -572 3422 -148
rect 2650 -600 3422 -572
rect -3422 -868 -2650 -840
rect -3422 -1292 -2734 -868
rect -2670 -1292 -2650 -868
rect -3422 -1320 -2650 -1292
rect -2410 -868 -1638 -840
rect -2410 -1292 -1722 -868
rect -1658 -1292 -1638 -868
rect -2410 -1320 -1638 -1292
rect -1398 -868 -626 -840
rect -1398 -1292 -710 -868
rect -646 -1292 -626 -868
rect -1398 -1320 -626 -1292
rect -386 -868 386 -840
rect -386 -1292 302 -868
rect 366 -1292 386 -868
rect -386 -1320 386 -1292
rect 626 -868 1398 -840
rect 626 -1292 1314 -868
rect 1378 -1292 1398 -868
rect 626 -1320 1398 -1292
rect 1638 -868 2410 -840
rect 1638 -1292 2326 -868
rect 2390 -1292 2410 -868
rect 1638 -1320 2410 -1292
rect 2650 -868 3422 -840
rect 2650 -1292 3338 -868
rect 3402 -1292 3422 -868
rect 2650 -1320 3422 -1292
rect -3422 -1588 -2650 -1560
rect -3422 -2012 -2734 -1588
rect -2670 -2012 -2650 -1588
rect -3422 -2040 -2650 -2012
rect -2410 -1588 -1638 -1560
rect -2410 -2012 -1722 -1588
rect -1658 -2012 -1638 -1588
rect -2410 -2040 -1638 -2012
rect -1398 -1588 -626 -1560
rect -1398 -2012 -710 -1588
rect -646 -2012 -626 -1588
rect -1398 -2040 -626 -2012
rect -386 -1588 386 -1560
rect -386 -2012 302 -1588
rect 366 -2012 386 -1588
rect -386 -2040 386 -2012
rect 626 -1588 1398 -1560
rect 626 -2012 1314 -1588
rect 1378 -2012 1398 -1588
rect 626 -2040 1398 -2012
rect 1638 -1588 2410 -1560
rect 1638 -2012 2326 -1588
rect 2390 -2012 2410 -1588
rect 1638 -2040 2410 -2012
rect 2650 -1588 3422 -1560
rect 2650 -2012 3338 -1588
rect 3402 -2012 3422 -1588
rect 2650 -2040 3422 -2012
<< via3 >>
rect -2734 1588 -2670 2012
rect -1722 1588 -1658 2012
rect -710 1588 -646 2012
rect 302 1588 366 2012
rect 1314 1588 1378 2012
rect 2326 1588 2390 2012
rect 3338 1588 3402 2012
rect -2734 868 -2670 1292
rect -1722 868 -1658 1292
rect -710 868 -646 1292
rect 302 868 366 1292
rect 1314 868 1378 1292
rect 2326 868 2390 1292
rect 3338 868 3402 1292
rect -2734 148 -2670 572
rect -1722 148 -1658 572
rect -710 148 -646 572
rect 302 148 366 572
rect 1314 148 1378 572
rect 2326 148 2390 572
rect 3338 148 3402 572
rect -2734 -572 -2670 -148
rect -1722 -572 -1658 -148
rect -710 -572 -646 -148
rect 302 -572 366 -148
rect 1314 -572 1378 -148
rect 2326 -572 2390 -148
rect 3338 -572 3402 -148
rect -2734 -1292 -2670 -868
rect -1722 -1292 -1658 -868
rect -710 -1292 -646 -868
rect 302 -1292 366 -868
rect 1314 -1292 1378 -868
rect 2326 -1292 2390 -868
rect 3338 -1292 3402 -868
rect -2734 -2012 -2670 -1588
rect -1722 -2012 -1658 -1588
rect -710 -2012 -646 -1588
rect 302 -2012 366 -1588
rect 1314 -2012 1378 -1588
rect 2326 -2012 2390 -1588
rect 3338 -2012 3402 -1588
<< mimcap >>
rect -3382 1960 -2982 2000
rect -3382 1640 -3342 1960
rect -3022 1640 -2982 1960
rect -3382 1600 -2982 1640
rect -2370 1960 -1970 2000
rect -2370 1640 -2330 1960
rect -2010 1640 -1970 1960
rect -2370 1600 -1970 1640
rect -1358 1960 -958 2000
rect -1358 1640 -1318 1960
rect -998 1640 -958 1960
rect -1358 1600 -958 1640
rect -346 1960 54 2000
rect -346 1640 -306 1960
rect 14 1640 54 1960
rect -346 1600 54 1640
rect 666 1960 1066 2000
rect 666 1640 706 1960
rect 1026 1640 1066 1960
rect 666 1600 1066 1640
rect 1678 1960 2078 2000
rect 1678 1640 1718 1960
rect 2038 1640 2078 1960
rect 1678 1600 2078 1640
rect 2690 1960 3090 2000
rect 2690 1640 2730 1960
rect 3050 1640 3090 1960
rect 2690 1600 3090 1640
rect -3382 1240 -2982 1280
rect -3382 920 -3342 1240
rect -3022 920 -2982 1240
rect -3382 880 -2982 920
rect -2370 1240 -1970 1280
rect -2370 920 -2330 1240
rect -2010 920 -1970 1240
rect -2370 880 -1970 920
rect -1358 1240 -958 1280
rect -1358 920 -1318 1240
rect -998 920 -958 1240
rect -1358 880 -958 920
rect -346 1240 54 1280
rect -346 920 -306 1240
rect 14 920 54 1240
rect -346 880 54 920
rect 666 1240 1066 1280
rect 666 920 706 1240
rect 1026 920 1066 1240
rect 666 880 1066 920
rect 1678 1240 2078 1280
rect 1678 920 1718 1240
rect 2038 920 2078 1240
rect 1678 880 2078 920
rect 2690 1240 3090 1280
rect 2690 920 2730 1240
rect 3050 920 3090 1240
rect 2690 880 3090 920
rect -3382 520 -2982 560
rect -3382 200 -3342 520
rect -3022 200 -2982 520
rect -3382 160 -2982 200
rect -2370 520 -1970 560
rect -2370 200 -2330 520
rect -2010 200 -1970 520
rect -2370 160 -1970 200
rect -1358 520 -958 560
rect -1358 200 -1318 520
rect -998 200 -958 520
rect -1358 160 -958 200
rect -346 520 54 560
rect -346 200 -306 520
rect 14 200 54 520
rect -346 160 54 200
rect 666 520 1066 560
rect 666 200 706 520
rect 1026 200 1066 520
rect 666 160 1066 200
rect 1678 520 2078 560
rect 1678 200 1718 520
rect 2038 200 2078 520
rect 1678 160 2078 200
rect 2690 520 3090 560
rect 2690 200 2730 520
rect 3050 200 3090 520
rect 2690 160 3090 200
rect -3382 -200 -2982 -160
rect -3382 -520 -3342 -200
rect -3022 -520 -2982 -200
rect -3382 -560 -2982 -520
rect -2370 -200 -1970 -160
rect -2370 -520 -2330 -200
rect -2010 -520 -1970 -200
rect -2370 -560 -1970 -520
rect -1358 -200 -958 -160
rect -1358 -520 -1318 -200
rect -998 -520 -958 -200
rect -1358 -560 -958 -520
rect -346 -200 54 -160
rect -346 -520 -306 -200
rect 14 -520 54 -200
rect -346 -560 54 -520
rect 666 -200 1066 -160
rect 666 -520 706 -200
rect 1026 -520 1066 -200
rect 666 -560 1066 -520
rect 1678 -200 2078 -160
rect 1678 -520 1718 -200
rect 2038 -520 2078 -200
rect 1678 -560 2078 -520
rect 2690 -200 3090 -160
rect 2690 -520 2730 -200
rect 3050 -520 3090 -200
rect 2690 -560 3090 -520
rect -3382 -920 -2982 -880
rect -3382 -1240 -3342 -920
rect -3022 -1240 -2982 -920
rect -3382 -1280 -2982 -1240
rect -2370 -920 -1970 -880
rect -2370 -1240 -2330 -920
rect -2010 -1240 -1970 -920
rect -2370 -1280 -1970 -1240
rect -1358 -920 -958 -880
rect -1358 -1240 -1318 -920
rect -998 -1240 -958 -920
rect -1358 -1280 -958 -1240
rect -346 -920 54 -880
rect -346 -1240 -306 -920
rect 14 -1240 54 -920
rect -346 -1280 54 -1240
rect 666 -920 1066 -880
rect 666 -1240 706 -920
rect 1026 -1240 1066 -920
rect 666 -1280 1066 -1240
rect 1678 -920 2078 -880
rect 1678 -1240 1718 -920
rect 2038 -1240 2078 -920
rect 1678 -1280 2078 -1240
rect 2690 -920 3090 -880
rect 2690 -1240 2730 -920
rect 3050 -1240 3090 -920
rect 2690 -1280 3090 -1240
rect -3382 -1640 -2982 -1600
rect -3382 -1960 -3342 -1640
rect -3022 -1960 -2982 -1640
rect -3382 -2000 -2982 -1960
rect -2370 -1640 -1970 -1600
rect -2370 -1960 -2330 -1640
rect -2010 -1960 -1970 -1640
rect -2370 -2000 -1970 -1960
rect -1358 -1640 -958 -1600
rect -1358 -1960 -1318 -1640
rect -998 -1960 -958 -1640
rect -1358 -2000 -958 -1960
rect -346 -1640 54 -1600
rect -346 -1960 -306 -1640
rect 14 -1960 54 -1640
rect -346 -2000 54 -1960
rect 666 -1640 1066 -1600
rect 666 -1960 706 -1640
rect 1026 -1960 1066 -1640
rect 666 -2000 1066 -1960
rect 1678 -1640 2078 -1600
rect 1678 -1960 1718 -1640
rect 2038 -1960 2078 -1640
rect 1678 -2000 2078 -1960
rect 2690 -1640 3090 -1600
rect 2690 -1960 2730 -1640
rect 3050 -1960 3090 -1640
rect 2690 -2000 3090 -1960
<< mimcapcontact >>
rect -3342 1640 -3022 1960
rect -2330 1640 -2010 1960
rect -1318 1640 -998 1960
rect -306 1640 14 1960
rect 706 1640 1026 1960
rect 1718 1640 2038 1960
rect 2730 1640 3050 1960
rect -3342 920 -3022 1240
rect -2330 920 -2010 1240
rect -1318 920 -998 1240
rect -306 920 14 1240
rect 706 920 1026 1240
rect 1718 920 2038 1240
rect 2730 920 3050 1240
rect -3342 200 -3022 520
rect -2330 200 -2010 520
rect -1318 200 -998 520
rect -306 200 14 520
rect 706 200 1026 520
rect 1718 200 2038 520
rect 2730 200 3050 520
rect -3342 -520 -3022 -200
rect -2330 -520 -2010 -200
rect -1318 -520 -998 -200
rect -306 -520 14 -200
rect 706 -520 1026 -200
rect 1718 -520 2038 -200
rect 2730 -520 3050 -200
rect -3342 -1240 -3022 -920
rect -2330 -1240 -2010 -920
rect -1318 -1240 -998 -920
rect -306 -1240 14 -920
rect 706 -1240 1026 -920
rect 1718 -1240 2038 -920
rect 2730 -1240 3050 -920
rect -3342 -1960 -3022 -1640
rect -2330 -1960 -2010 -1640
rect -1318 -1960 -998 -1640
rect -306 -1960 14 -1640
rect 706 -1960 1026 -1640
rect 1718 -1960 2038 -1640
rect 2730 -1960 3050 -1640
<< metal4 >>
rect -2750 2012 -2654 2028
rect -3343 1960 -3021 1961
rect -3343 1640 -3342 1960
rect -3022 1640 -3021 1960
rect -3343 1639 -3021 1640
rect -2750 1588 -2734 2012
rect -2670 1588 -2654 2012
rect -1738 2012 -1642 2028
rect -2331 1960 -2009 1961
rect -2331 1640 -2330 1960
rect -2010 1640 -2009 1960
rect -2331 1639 -2009 1640
rect -2750 1572 -2654 1588
rect -1738 1588 -1722 2012
rect -1658 1588 -1642 2012
rect -726 2012 -630 2028
rect -1319 1960 -997 1961
rect -1319 1640 -1318 1960
rect -998 1640 -997 1960
rect -1319 1639 -997 1640
rect -1738 1572 -1642 1588
rect -726 1588 -710 2012
rect -646 1588 -630 2012
rect 286 2012 382 2028
rect -307 1960 15 1961
rect -307 1640 -306 1960
rect 14 1640 15 1960
rect -307 1639 15 1640
rect -726 1572 -630 1588
rect 286 1588 302 2012
rect 366 1588 382 2012
rect 1298 2012 1394 2028
rect 705 1960 1027 1961
rect 705 1640 706 1960
rect 1026 1640 1027 1960
rect 705 1639 1027 1640
rect 286 1572 382 1588
rect 1298 1588 1314 2012
rect 1378 1588 1394 2012
rect 2310 2012 2406 2028
rect 1717 1960 2039 1961
rect 1717 1640 1718 1960
rect 2038 1640 2039 1960
rect 1717 1639 2039 1640
rect 1298 1572 1394 1588
rect 2310 1588 2326 2012
rect 2390 1588 2406 2012
rect 3322 2012 3418 2028
rect 2729 1960 3051 1961
rect 2729 1640 2730 1960
rect 3050 1640 3051 1960
rect 2729 1639 3051 1640
rect 2310 1572 2406 1588
rect 3322 1588 3338 2012
rect 3402 1588 3418 2012
rect 3322 1572 3418 1588
rect -2750 1292 -2654 1308
rect -3343 1240 -3021 1241
rect -3343 920 -3342 1240
rect -3022 920 -3021 1240
rect -3343 919 -3021 920
rect -2750 868 -2734 1292
rect -2670 868 -2654 1292
rect -1738 1292 -1642 1308
rect -2331 1240 -2009 1241
rect -2331 920 -2330 1240
rect -2010 920 -2009 1240
rect -2331 919 -2009 920
rect -2750 852 -2654 868
rect -1738 868 -1722 1292
rect -1658 868 -1642 1292
rect -726 1292 -630 1308
rect -1319 1240 -997 1241
rect -1319 920 -1318 1240
rect -998 920 -997 1240
rect -1319 919 -997 920
rect -1738 852 -1642 868
rect -726 868 -710 1292
rect -646 868 -630 1292
rect 286 1292 382 1308
rect -307 1240 15 1241
rect -307 920 -306 1240
rect 14 920 15 1240
rect -307 919 15 920
rect -726 852 -630 868
rect 286 868 302 1292
rect 366 868 382 1292
rect 1298 1292 1394 1308
rect 705 1240 1027 1241
rect 705 920 706 1240
rect 1026 920 1027 1240
rect 705 919 1027 920
rect 286 852 382 868
rect 1298 868 1314 1292
rect 1378 868 1394 1292
rect 2310 1292 2406 1308
rect 1717 1240 2039 1241
rect 1717 920 1718 1240
rect 2038 920 2039 1240
rect 1717 919 2039 920
rect 1298 852 1394 868
rect 2310 868 2326 1292
rect 2390 868 2406 1292
rect 3322 1292 3418 1308
rect 2729 1240 3051 1241
rect 2729 920 2730 1240
rect 3050 920 3051 1240
rect 2729 919 3051 920
rect 2310 852 2406 868
rect 3322 868 3338 1292
rect 3402 868 3418 1292
rect 3322 852 3418 868
rect -2750 572 -2654 588
rect -3343 520 -3021 521
rect -3343 200 -3342 520
rect -3022 200 -3021 520
rect -3343 199 -3021 200
rect -2750 148 -2734 572
rect -2670 148 -2654 572
rect -1738 572 -1642 588
rect -2331 520 -2009 521
rect -2331 200 -2330 520
rect -2010 200 -2009 520
rect -2331 199 -2009 200
rect -2750 132 -2654 148
rect -1738 148 -1722 572
rect -1658 148 -1642 572
rect -726 572 -630 588
rect -1319 520 -997 521
rect -1319 200 -1318 520
rect -998 200 -997 520
rect -1319 199 -997 200
rect -1738 132 -1642 148
rect -726 148 -710 572
rect -646 148 -630 572
rect 286 572 382 588
rect -307 520 15 521
rect -307 200 -306 520
rect 14 200 15 520
rect -307 199 15 200
rect -726 132 -630 148
rect 286 148 302 572
rect 366 148 382 572
rect 1298 572 1394 588
rect 705 520 1027 521
rect 705 200 706 520
rect 1026 200 1027 520
rect 705 199 1027 200
rect 286 132 382 148
rect 1298 148 1314 572
rect 1378 148 1394 572
rect 2310 572 2406 588
rect 1717 520 2039 521
rect 1717 200 1718 520
rect 2038 200 2039 520
rect 1717 199 2039 200
rect 1298 132 1394 148
rect 2310 148 2326 572
rect 2390 148 2406 572
rect 3322 572 3418 588
rect 2729 520 3051 521
rect 2729 200 2730 520
rect 3050 200 3051 520
rect 2729 199 3051 200
rect 2310 132 2406 148
rect 3322 148 3338 572
rect 3402 148 3418 572
rect 3322 132 3418 148
rect -2750 -148 -2654 -132
rect -3343 -200 -3021 -199
rect -3343 -520 -3342 -200
rect -3022 -520 -3021 -200
rect -3343 -521 -3021 -520
rect -2750 -572 -2734 -148
rect -2670 -572 -2654 -148
rect -1738 -148 -1642 -132
rect -2331 -200 -2009 -199
rect -2331 -520 -2330 -200
rect -2010 -520 -2009 -200
rect -2331 -521 -2009 -520
rect -2750 -588 -2654 -572
rect -1738 -572 -1722 -148
rect -1658 -572 -1642 -148
rect -726 -148 -630 -132
rect -1319 -200 -997 -199
rect -1319 -520 -1318 -200
rect -998 -520 -997 -200
rect -1319 -521 -997 -520
rect -1738 -588 -1642 -572
rect -726 -572 -710 -148
rect -646 -572 -630 -148
rect 286 -148 382 -132
rect -307 -200 15 -199
rect -307 -520 -306 -200
rect 14 -520 15 -200
rect -307 -521 15 -520
rect -726 -588 -630 -572
rect 286 -572 302 -148
rect 366 -572 382 -148
rect 1298 -148 1394 -132
rect 705 -200 1027 -199
rect 705 -520 706 -200
rect 1026 -520 1027 -200
rect 705 -521 1027 -520
rect 286 -588 382 -572
rect 1298 -572 1314 -148
rect 1378 -572 1394 -148
rect 2310 -148 2406 -132
rect 1717 -200 2039 -199
rect 1717 -520 1718 -200
rect 2038 -520 2039 -200
rect 1717 -521 2039 -520
rect 1298 -588 1394 -572
rect 2310 -572 2326 -148
rect 2390 -572 2406 -148
rect 3322 -148 3418 -132
rect 2729 -200 3051 -199
rect 2729 -520 2730 -200
rect 3050 -520 3051 -200
rect 2729 -521 3051 -520
rect 2310 -588 2406 -572
rect 3322 -572 3338 -148
rect 3402 -572 3418 -148
rect 3322 -588 3418 -572
rect -2750 -868 -2654 -852
rect -3343 -920 -3021 -919
rect -3343 -1240 -3342 -920
rect -3022 -1240 -3021 -920
rect -3343 -1241 -3021 -1240
rect -2750 -1292 -2734 -868
rect -2670 -1292 -2654 -868
rect -1738 -868 -1642 -852
rect -2331 -920 -2009 -919
rect -2331 -1240 -2330 -920
rect -2010 -1240 -2009 -920
rect -2331 -1241 -2009 -1240
rect -2750 -1308 -2654 -1292
rect -1738 -1292 -1722 -868
rect -1658 -1292 -1642 -868
rect -726 -868 -630 -852
rect -1319 -920 -997 -919
rect -1319 -1240 -1318 -920
rect -998 -1240 -997 -920
rect -1319 -1241 -997 -1240
rect -1738 -1308 -1642 -1292
rect -726 -1292 -710 -868
rect -646 -1292 -630 -868
rect 286 -868 382 -852
rect -307 -920 15 -919
rect -307 -1240 -306 -920
rect 14 -1240 15 -920
rect -307 -1241 15 -1240
rect -726 -1308 -630 -1292
rect 286 -1292 302 -868
rect 366 -1292 382 -868
rect 1298 -868 1394 -852
rect 705 -920 1027 -919
rect 705 -1240 706 -920
rect 1026 -1240 1027 -920
rect 705 -1241 1027 -1240
rect 286 -1308 382 -1292
rect 1298 -1292 1314 -868
rect 1378 -1292 1394 -868
rect 2310 -868 2406 -852
rect 1717 -920 2039 -919
rect 1717 -1240 1718 -920
rect 2038 -1240 2039 -920
rect 1717 -1241 2039 -1240
rect 1298 -1308 1394 -1292
rect 2310 -1292 2326 -868
rect 2390 -1292 2406 -868
rect 3322 -868 3418 -852
rect 2729 -920 3051 -919
rect 2729 -1240 2730 -920
rect 3050 -1240 3051 -920
rect 2729 -1241 3051 -1240
rect 2310 -1308 2406 -1292
rect 3322 -1292 3338 -868
rect 3402 -1292 3418 -868
rect 3322 -1308 3418 -1292
rect -2750 -1588 -2654 -1572
rect -3343 -1640 -3021 -1639
rect -3343 -1960 -3342 -1640
rect -3022 -1960 -3021 -1640
rect -3343 -1961 -3021 -1960
rect -2750 -2012 -2734 -1588
rect -2670 -2012 -2654 -1588
rect -1738 -1588 -1642 -1572
rect -2331 -1640 -2009 -1639
rect -2331 -1960 -2330 -1640
rect -2010 -1960 -2009 -1640
rect -2331 -1961 -2009 -1960
rect -2750 -2028 -2654 -2012
rect -1738 -2012 -1722 -1588
rect -1658 -2012 -1642 -1588
rect -726 -1588 -630 -1572
rect -1319 -1640 -997 -1639
rect -1319 -1960 -1318 -1640
rect -998 -1960 -997 -1640
rect -1319 -1961 -997 -1960
rect -1738 -2028 -1642 -2012
rect -726 -2012 -710 -1588
rect -646 -2012 -630 -1588
rect 286 -1588 382 -1572
rect -307 -1640 15 -1639
rect -307 -1960 -306 -1640
rect 14 -1960 15 -1640
rect -307 -1961 15 -1960
rect -726 -2028 -630 -2012
rect 286 -2012 302 -1588
rect 366 -2012 382 -1588
rect 1298 -1588 1394 -1572
rect 705 -1640 1027 -1639
rect 705 -1960 706 -1640
rect 1026 -1960 1027 -1640
rect 705 -1961 1027 -1960
rect 286 -2028 382 -2012
rect 1298 -2012 1314 -1588
rect 1378 -2012 1394 -1588
rect 2310 -1588 2406 -1572
rect 1717 -1640 2039 -1639
rect 1717 -1960 1718 -1640
rect 2038 -1960 2039 -1640
rect 1717 -1961 2039 -1960
rect 1298 -2028 1394 -2012
rect 2310 -2012 2326 -1588
rect 2390 -2012 2406 -1588
rect 3322 -1588 3418 -1572
rect 2729 -1640 3051 -1639
rect 2729 -1960 2730 -1640
rect 3050 -1960 3051 -1640
rect 2729 -1961 3051 -1960
rect 2310 -2028 2406 -2012
rect 3322 -2012 3338 -1588
rect 3402 -2012 3418 -1588
rect 3322 -2028 3418 -2012
<< properties >>
string FIXED_BBOX 2650 1560 3130 2040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.0 l 2.0 val 9.52 carea 2.00 cperi 0.19 nx 7 ny 6 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
