magic
tech sky130A
magscale 1 2
timestamp 1751021419
<< nwell >>
rect -3098 5083 -2883 13397
<< metal1 >>
rect -3151 12991 -2366 13176
rect -3151 12806 -2360 12991
rect -3154 10640 -2369 10825
rect -2682 7950 -2622 8044
rect -3232 5142 -2903 5172
rect -3232 5020 -2987 5142
rect -2931 5020 -2903 5142
rect -3232 5008 -2903 5020
rect -2682 2006 -2622 7890
rect -5386 -145 -5063 1009
rect -4371 828 -4365 888
rect -4305 828 -4299 888
rect -4369 -596 -4363 -474
rect -4307 -596 -4301 -474
rect -2682 -541 -2622 1946
rect -2594 8038 -2534 8044
rect -2594 1886 -2534 7978
rect -2594 1820 -2534 1826
rect -2506 3964 -2447 4064
rect -2418 4058 -2358 4064
rect -2506 3938 -2446 3964
rect -2506 497 -2446 3878
rect -2506 431 -2446 437
rect -2418 585 -2358 3998
rect -2682 -601 -2647 -541
rect -2587 -601 -2579 -541
rect -2418 -546 -2358 525
rect -2529 -606 -2521 -546
rect -2461 -606 -2358 -546
rect -3519 -2195 -2921 -1795
rect -3519 -3848 -3119 -2195
rect -3278 -4683 -3272 -4630
rect -3150 -4683 -3144 -4630
<< via1 >>
rect -2682 7890 -2622 7950
rect -2987 5020 -2931 5142
rect -2682 1946 -2622 2006
rect -4365 828 -4305 888
rect -4194 -404 -4138 -282
rect -4363 -596 -4307 -474
rect -2594 7978 -2534 8038
rect -2255 6419 -2195 6479
rect -2594 1826 -2534 1886
rect -2418 3998 -2358 4058
rect -2506 3878 -2446 3938
rect -2506 437 -2446 497
rect -721 3147 -661 3207
rect -2255 1388 -2195 1448
rect -2418 525 -2358 585
rect -2647 -601 -2587 -541
rect -2255 148 -2195 208
rect -2521 -606 -2461 -546
rect -4868 -1524 -4808 -1464
rect -3272 -4683 -3150 -4627
<< metal2 >>
rect -4020 8126 -3960 8188
rect -4020 8066 -1954 8126
rect -2688 7978 -2594 8038
rect -2534 7978 -2056 8038
rect -2688 7890 -2682 7950
rect -2622 7890 -2051 7950
rect -4736 7306 -3090 7308
rect -4736 7250 -3221 7306
rect -3099 7250 -3090 7306
rect -4736 7248 -3090 7250
rect -2846 6477 -2255 6479
rect -2846 6421 -2837 6477
rect -2715 6421 -2255 6477
rect -2846 6419 -2255 6421
rect -2195 6419 -2189 6479
rect -5488 6230 -3090 6232
rect -5488 6174 -3221 6230
rect -3099 6174 -3090 6230
rect -5488 6172 -3090 6174
rect -2996 5020 -2987 5142
rect -2931 5020 -2922 5142
rect -3696 3998 -2418 4058
rect -2358 3998 -2352 4058
rect -3696 3878 -2506 3938
rect -2446 3878 -2352 3938
rect -727 3147 -721 3207
rect -661 3205 -331 3207
rect -661 3149 -427 3205
rect -341 3149 -331 3205
rect -661 3147 -331 3149
rect -3696 1946 -2682 2006
rect -2622 1946 -2528 2006
rect -3696 1826 -2594 1886
rect -2534 1826 -2528 1886
rect -3230 1446 -2255 1448
rect -3230 1390 -3221 1446
rect -3099 1390 -2255 1446
rect -3230 1388 -2255 1390
rect -2195 1388 -2189 1448
rect -4372 972 -4296 982
rect -4372 888 -4362 972
rect -4306 888 -4296 972
rect -4372 860 -4365 888
rect -4305 860 -4296 888
rect -4365 822 -4305 828
rect -2512 525 -2418 585
rect -2358 525 -2052 585
rect -7297 470 -5466 472
rect -7297 414 -5532 470
rect -5476 414 -5466 470
rect -2512 437 -2506 497
rect -2446 437 -2052 497
rect -7297 412 -5466 414
rect -5888 148 -2255 208
rect -2195 148 -2189 208
rect -4203 -404 -4194 -282
rect -4138 -404 -4129 -282
rect -4372 -596 -4363 -474
rect -4307 -596 -4298 -474
rect -2655 -601 -2647 -541
rect -2587 -601 -2579 -541
rect -2529 -606 -2521 -546
rect -2461 -606 -2453 -546
rect -6545 -958 -5466 -956
rect -6545 -1014 -5532 -958
rect -5476 -1014 -5466 -958
rect -6545 -1016 -5466 -1014
rect -5542 -1466 -4868 -1464
rect -5542 -1522 -5532 -1466
rect -5476 -1522 -4868 -1466
rect -5542 -1524 -4868 -1522
rect -4808 -1524 -4802 -1464
rect -3281 -4683 -3272 -4627
rect -3150 -4683 -3141 -4627
<< via2 >>
rect -3221 7250 -3099 7306
rect -2837 6421 -2715 6477
rect -3221 6174 -3099 6230
rect -2987 5020 -2931 5142
rect -427 3149 -341 3205
rect -3221 1390 -3099 1446
rect -4362 888 -4306 972
rect -4362 860 -4306 888
rect -5532 414 -5476 470
rect -4194 -404 -4138 -282
rect -4363 -596 -4307 -474
rect -2645 -599 -2589 -543
rect -2519 -604 -2463 -548
rect -5532 -1014 -5476 -958
rect -5532 -1522 -5476 -1466
rect -3272 -4683 -3150 -4627
<< metal3 >>
rect -3226 7306 -3094 7311
rect -3226 7250 -3221 7306
rect -3099 7250 -3094 7306
rect -3226 6230 -3094 7250
rect -3226 6174 -3221 6230
rect -3099 6174 -3094 6230
rect -3226 1446 -3094 6174
rect -2842 6477 -2710 6482
rect -2842 6421 -2837 6477
rect -2715 6421 -2710 6477
rect -3226 1390 -3221 1446
rect -3099 1390 -3094 1446
rect -3226 982 -3094 1390
rect -4368 972 -3094 982
rect -4368 860 -4362 972
rect -4306 860 -3094 972
rect -4368 850 -3094 860
rect -3034 5142 -2902 5173
rect -3034 5020 -2987 5142
rect -2931 5020 -2902 5142
rect -5537 470 -5471 480
rect -5537 414 -5532 470
rect -5476 414 -5471 470
rect -5537 -958 -5471 414
rect -3034 -277 -2902 5020
rect -4203 -282 -2902 -277
rect -4203 -404 -4194 -282
rect -4138 -404 -2902 -282
rect -4203 -409 -2902 -404
rect -2842 -469 -2710 6421
rect -4372 -474 -2710 -469
rect -4372 -596 -4363 -474
rect -4307 -596 -2710 -474
rect -432 3205 -336 3210
rect -432 3149 -427 3205
rect -341 3149 -336 3205
rect -4372 -601 -2710 -596
rect -2650 -543 -2584 -533
rect -2650 -599 -2645 -543
rect -2589 -599 -2584 -543
rect -5537 -1014 -5532 -958
rect -5476 -1014 -5471 -958
rect -5537 -1466 -5471 -1014
rect -5537 -1522 -5532 -1466
rect -5476 -1522 -5471 -1466
rect -5537 -1532 -5471 -1522
rect -2650 -4538 -2584 -599
rect -2524 -548 -2458 -538
rect -2524 -604 -2519 -548
rect -2463 -604 -2458 -548
rect -2524 -4382 -2458 -604
rect -2524 -4478 -1333 -4382
rect -3288 -4627 -3119 -4622
rect -3288 -4683 -3272 -4627
rect -3150 -4683 -3119 -4627
rect -2650 -4634 -2347 -4538
rect -3288 -4718 -3119 -4683
rect -2443 -5990 -2347 -4634
rect -1429 -5838 -1333 -4478
rect -1429 -5902 -1412 -5838
rect -1348 -5902 -1333 -5838
rect -1429 -5903 -1333 -5902
rect -1429 -6168 -1333 -6152
rect -1429 -6232 -1412 -6168
rect -1348 -6232 -1333 -6168
rect -1429 -6710 -1333 -6232
rect -7048 -6806 -1333 -6710
rect -432 -7430 -336 3149
rect -496 -7526 -336 -7430
<< via3 >>
rect -1412 -5902 -1348 -5838
rect -1412 -6232 -1348 -6168
<< metal4 >>
rect -1429 -5838 -1333 -5837
rect -1429 -5902 -1412 -5838
rect -1348 -5902 -1333 -5838
rect -1429 -6168 -1333 -5902
rect -1429 -6232 -1412 -6168
rect -1348 -6232 -1333 -6168
rect -1429 -6233 -1333 -6232
use fcm_bias_ncell  fcm_bias_ncell_0
timestamp 1750066031
transform 1 0 -5053 0 1 400
box -36 -571 956 635
use fcm_bias_pcell  fcm_bias_pcell_0
timestamp 1750065844
transform 1 0 -5274 0 1 -1612
box 155 -1155 1207 1391
use opa_cap  opa_cap_0
timestamp 1750150226
transform 1 0 -7388 0 1 -15196
box -5008 6398 7908 10478
use opa_folded_cascode  opa_folded_cascode_0
timestamp 1750150351
transform 1 0 -2404 0 1 7738
box -543 -9959 2211 5484
use opa_input_and_self_bias  opa_input_and_self_bias_0
timestamp 1751017459
transform 1 0 -12418 0 1 -3832
box -44 -886 9367 17230
<< labels >>
flabel metal1 s -3668 2688 -3608 2748 0 FreeSans 320 0 0 0 N_IN
port 5 nsew
flabel metal1 s -691 3347 -631 3407 0 FreeSans 320 0 0 0 VOUT
port 6 nsew
flabel metal3 s -12283 13306 -12223 13366 0 FreeSans 800 0 0 0 ROUT
port 7 nsew
flabel metal1 s -2761 13050 -2701 13110 0 FreeSans 1600 0 0 0 VDDA
port 8 nsew
flabel metal1 s -3361 -3012 -3301 -2952 0 FreeSans 1600 0 0 0 GNDA
port 9 nsew
flabel metal2 s -12298 2532 -12238 2592 0 FreeSans 320 0 0 0 P_IN[0]
port 0 nsew
flabel metal2 s -12298 2620 -12238 2680 0 FreeSans 320 0 0 0 P_IN[1]
port 1 nsew
flabel metal2 s -12298 2708 -12238 2768 0 FreeSans 320 0 0 0 P_IN[2]
port 2 nsew
flabel metal2 s -12298 2796 -12238 2856 0 FreeSans 320 0 0 0 P_IN[3]
port 3 nsew
flabel metal2 s -12298 2884 -12238 2944 0 FreeSans 320 0 0 0 P_IN[4]
port 4 nsew
<< end >>
