magic
tech sky130A
timestamp 1749560624
<< metal1 >>
rect 770 -11382 800 -11308
rect 814 -11382 844 -11308
rect 858 -11382 888 -11308
rect 902 -11382 932 -11308
<< end >>
