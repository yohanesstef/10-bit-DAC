magic
tech sky130A
magscale 1 2
timestamp 1749523501
<< error_s >>
rect 1120 758 1126 764
rect 1174 758 1180 764
rect 1114 752 1120 758
rect 1180 752 1186 758
rect 1114 698 1120 704
rect 1180 698 1186 704
rect 1120 692 1126 698
rect 1174 692 1180 698
rect 844 670 850 676
rect 898 670 904 676
rect 838 664 844 670
rect 904 664 910 670
rect 838 610 844 616
rect 904 610 910 616
rect 844 604 850 610
rect 898 604 904 610
rect 568 582 574 588
rect 622 582 628 588
rect 562 576 568 582
rect 628 576 634 582
rect 562 522 568 528
rect 628 522 634 528
rect 568 516 574 522
rect 622 516 628 522
rect 292 494 298 500
rect 346 494 352 500
rect 286 488 292 494
rect 352 488 358 494
rect 286 434 292 440
rect 352 434 358 440
rect 292 428 298 434
rect 346 428 352 434
rect 16 406 22 412
rect 70 406 76 412
rect 10 400 16 406
rect 76 400 82 406
rect 10 346 16 352
rect 76 346 82 352
rect 16 340 22 346
rect 70 340 76 346
<< nwell >>
rect -156 -170 1564 438
<< mvnsubdiff >>
rect -90 360 1498 372
rect -90 326 18 360
rect 1390 326 1498 360
rect -90 314 1498 326
rect -90 264 -32 314
rect -90 4 -78 264
rect -44 4 -32 264
rect -90 -46 -32 4
rect 1440 264 1498 314
rect 1440 4 1452 264
rect 1486 4 1498 264
rect 1440 -46 1498 4
rect -90 -58 1498 -46
rect -90 -92 18 -58
rect 1390 -92 1498 -58
rect -90 -104 1498 -92
<< mvnsubdiffcont >>
rect 18 326 1390 360
rect -78 4 -44 264
rect 1452 4 1486 264
rect 18 -92 1390 -58
<< locali >>
rect -78 326 18 360
rect 1390 326 1486 360
rect -78 264 -44 326
rect -78 -58 -44 4
rect 1452 264 1486 326
rect 1452 -58 1486 4
rect -78 -92 18 -58
rect 1390 -92 1486 -58
<< metal1 >>
rect 1120 758 1180 764
rect 844 670 904 676
rect 568 582 628 588
rect 292 494 352 500
rect 16 406 76 412
rect 16 56 76 346
rect 292 56 352 434
rect 568 56 628 522
rect 844 56 904 610
rect 1120 56 1180 698
<< via1 >>
rect 1120 698 1180 758
rect 844 610 904 670
rect 568 522 628 582
rect 292 434 352 494
rect 16 346 76 406
use hpmos_1  hpmos_1_1 ~/10-bit-DAC/mag
timestamp 1749230053
transform 1 0 -774 0 1 3211
box 1856 -3221 2204 -2971
use hpmos_4  hpmos_4_0 ~/10-bit-DAC/mag
timestamp 1749384553
transform 1 0 -400 0 1 -41
box 378 31 1554 281
<< end >>
