magic
tech sky130A
magscale 1 2
timestamp 1749289931
<< metal1 >>
rect 9957 -15154 10017 -14830
rect 9944 -15740 10017 -15154
rect 10045 -15802 10105 -14830
rect 10032 -16388 10105 -15802
rect 10133 -16450 10193 -14830
rect 10058 -17036 10193 -16450
rect 10221 -17098 10281 -14830
rect 10099 -17360 10281 -17098
<< end >>
