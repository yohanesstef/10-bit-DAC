magic
tech sky130A
magscale 1 2
timestamp 1749057406
<< pwell >>
rect -307 -1068 307 1068
<< psubdiff >>
rect -271 998 -175 1032
rect 175 998 271 1032
rect -271 936 -237 998
rect 237 936 271 998
rect -271 -998 -237 -936
rect 237 -998 271 -936
rect -271 -1032 -175 -998
rect 175 -1032 271 -998
<< psubdiffcont >>
rect -175 998 175 1032
rect -271 -936 -237 936
rect 237 -936 271 936
rect -175 -1032 175 -998
<< xpolycontact >>
rect -141 470 141 902
rect -141 -902 141 -470
<< xpolyres >>
rect -141 -470 141 470
<< locali >>
rect -271 998 -175 1032
rect 175 998 271 1032
rect -271 936 -237 998
rect 237 936 271 998
rect -271 -998 -237 -936
rect 237 -998 271 -936
rect -271 -1032 -175 -998
rect 175 -1032 271 -998
<< viali >>
rect -125 487 125 884
rect -125 -884 125 -487
<< metal1 >>
rect -131 884 131 896
rect -131 487 -125 884
rect 125 487 131 884
rect -131 475 131 487
rect -131 -487 131 -475
rect -131 -884 -125 -487
rect 125 -884 131 -487
rect -131 -896 131 -884
<< properties >>
string FIXED_BBOX -254 -1015 254 1015
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 4.859 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 7.159k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
