magic
tech sky130A
magscale 1 2
timestamp 1749007001
<< xpolycontact >>
rect -141 516 141 948
rect -141 -948 141 -516
<< xpolyres >>
rect -141 -516 141 516
<< viali >>
rect -125 533 125 930
rect -125 -930 125 -533
<< metal1 >>
rect -131 930 131 942
rect -131 533 -125 930
rect 125 533 131 930
rect -131 521 131 533
rect -131 -533 131 -521
rect -131 -930 -125 -533
rect 125 -930 131 -533
rect -131 -942 131 -930
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 5.32 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 7.813k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
