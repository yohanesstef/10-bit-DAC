magic
tech sky130A
magscale 1 2
timestamp 1749057406
<< pwell >>
rect -307 -914 307 914
<< psubdiff >>
rect -271 844 -175 878
rect 175 844 271 878
rect -271 782 -237 844
rect 237 782 271 844
rect -271 -844 -237 -782
rect 237 -844 271 -782
rect -271 -878 -175 -844
rect 175 -878 271 -844
<< psubdiffcont >>
rect -175 844 175 878
rect -271 -782 -237 782
rect 237 -782 271 782
rect -175 -878 175 -844
<< xpolycontact >>
rect -141 316 141 748
rect -141 -748 141 -316
<< xpolyres >>
rect -141 -316 141 316
<< locali >>
rect -271 844 -175 878
rect 175 844 271 878
rect -271 782 -237 844
rect 237 782 271 844
rect -271 -844 -237 -782
rect 237 -844 271 -782
rect -271 -878 -175 -844
rect 175 -878 271 -844
<< viali >>
rect -125 333 125 730
rect -125 -730 125 -333
<< metal1 >>
rect -131 730 131 742
rect -131 333 -125 730
rect 125 333 131 730
rect -131 321 131 333
rect -131 -333 131 -321
rect -131 -730 -125 -333
rect 125 -730 131 -333
rect -131 -742 131 -730
<< properties >>
string FIXED_BBOX -254 -861 254 861
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 3.321 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 4.977k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
