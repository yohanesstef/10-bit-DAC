magic
tech sky130A
magscale 1 2
timestamp 1751017459
<< locali >>
rect 49 3650 8723 3730
rect 49 -40 7023 40
<< metal2 >>
rect 4745 6445 6152 6447
rect 4745 6389 6086 6445
rect 6142 6389 6152 6445
rect 4745 6387 6152 6389
rect 4623 6357 7880 6359
rect 4623 6301 7814 6357
rect 7870 6301 7880 6357
rect 4623 6299 7880 6301
rect 3921 6093 5368 6095
rect 3921 6037 3931 6093
rect 3987 6037 5368 6093
rect 3921 6035 5368 6037
rect 2620 5917 4956 5919
rect 2620 5861 2630 5917
rect 2686 5861 4956 5917
rect 2620 5859 4956 5861
rect 892 5830 949 5831
rect 892 5774 902 5830
rect 958 5774 968 5830
rect 892 5771 949 5774
rect 892 5105 922 5107
rect 892 5049 902 5105
rect 958 5049 968 5105
rect 892 5047 922 5049
rect 2620 5017 3128 5019
rect 2620 4961 2630 5017
rect 2686 4961 3128 5017
rect 2620 4959 3128 4961
rect 3926 4841 3997 4843
rect 3921 4785 3931 4841
rect 3987 4785 3997 4841
rect 3926 4783 3997 4785
rect 4747 4577 7880 4579
rect 4747 4521 7814 4577
rect 7870 4521 7880 4577
rect 4747 4519 7880 4521
rect 4629 4489 6152 4491
rect 4629 4433 6086 4489
rect 6142 4433 6152 4489
rect 4629 4431 6152 4433
rect 902 2695 958 2705
rect 902 2629 958 2639
rect 2630 2695 2686 2705
rect 2630 2629 2686 2639
rect 4358 2695 4414 2705
rect 4358 2629 4414 2639
rect 6086 2695 6142 2705
rect 6086 2629 6142 2639
rect 7814 2695 7870 2705
rect 7814 2629 7870 2639
rect 902 643 958 653
rect 902 577 958 587
rect 2630 643 2686 653
rect 2630 577 2686 587
rect 4358 643 4414 653
rect 4358 577 4414 587
rect 6086 643 6142 653
rect 6086 577 6142 587
rect 7814 643 7870 653
rect 7814 577 7870 587
rect 892 -271 902 -215
rect 958 -271 968 -215
rect 2966 -655 4424 -653
rect 2966 -711 4358 -655
rect 4414 -711 4424 -655
rect 2966 -713 4424 -711
rect 2620 -799 2630 -743
rect 2686 -799 2696 -743
rect 3183 -1183 7145 -1181
rect 3183 -1239 7079 -1183
rect 7135 -1239 7145 -1183
rect 3183 -1241 7145 -1239
rect 3889 -1271 6152 -1269
rect 3889 -1327 6086 -1271
rect 6142 -1327 6152 -1271
rect 3889 -1329 6152 -1327
rect 3255 -1819 6152 -1817
rect 3255 -1875 6086 -1819
rect 6142 -1875 6152 -1819
rect 3255 -1877 6152 -1875
rect 3889 -1907 7145 -1905
rect 3889 -1963 7079 -1907
rect 7135 -1963 7145 -1907
rect 3889 -1965 7145 -1963
rect 2620 -2347 2737 -2345
rect 2620 -2403 2630 -2347
rect 2686 -2403 2737 -2347
rect 2620 -2405 2737 -2403
rect 4348 -2491 4358 -2435
rect 4414 -2491 4424 -2435
rect 892 -2875 1561 -2873
rect 892 -2931 902 -2875
rect 958 -2931 1561 -2875
rect 892 -2933 1561 -2931
<< via2 >>
rect 6086 6389 6142 6445
rect 7814 6301 7870 6357
rect 3931 6037 3987 6093
rect 2630 5861 2686 5917
rect 902 5774 958 5830
rect 902 5049 958 5105
rect 2630 4961 2686 5017
rect 3931 4785 3987 4841
rect 7814 4521 7870 4577
rect 6086 4433 6142 4489
rect 902 2639 958 2695
rect 2630 2639 2686 2695
rect 4358 2639 4414 2695
rect 6086 2639 6142 2695
rect 7814 2639 7870 2695
rect 902 587 958 643
rect 2630 587 2686 643
rect 4358 587 4414 643
rect 6086 587 6142 643
rect 7814 587 7870 643
rect 902 -271 958 -215
rect 4358 -711 4414 -655
rect 2630 -799 2686 -743
rect 7079 -1239 7135 -1183
rect 6086 -1327 6142 -1271
rect 6086 -1875 6142 -1819
rect 7079 -1963 7135 -1907
rect 2630 -2403 2686 -2347
rect 4358 -2491 4414 -2435
rect 902 -2931 958 -2875
<< metal3 >>
rect 2625 5917 2691 7179
rect 6081 6445 6147 6450
rect 6081 6389 6086 6445
rect 6142 6389 6147 6445
rect 2625 5861 2630 5917
rect 2686 5861 2691 5917
rect 897 5830 963 5840
rect 897 5774 902 5830
rect 958 5774 963 5830
rect 897 5105 963 5774
rect 897 5049 902 5105
rect 958 5049 963 5105
rect 897 2695 963 5049
rect 897 2639 902 2695
rect 958 2639 963 2695
rect 897 2629 963 2639
rect 2625 5017 2691 5861
rect 2625 4961 2630 5017
rect 2686 4961 2691 5017
rect 2625 2695 2691 4961
rect 3926 6093 3992 6103
rect 3926 6037 3931 6093
rect 3987 6037 3992 6093
rect 3926 4841 3992 6037
rect 3926 4785 3931 4841
rect 3987 4785 3992 4841
rect 3926 3724 3992 4785
rect 6081 4489 6147 6389
rect 6081 4433 6086 4489
rect 6142 4433 6147 4489
rect 3926 3658 4419 3724
rect 2625 2639 2630 2695
rect 2686 2639 2691 2695
rect 2625 2629 2691 2639
rect 4353 2695 4419 3658
rect 4353 2639 4358 2695
rect 4414 2639 4419 2695
rect 4353 2629 4419 2639
rect 6081 2695 6147 4433
rect 6081 2639 6086 2695
rect 6142 2639 6147 2695
rect 6081 2629 6147 2639
rect 7809 6357 7875 6362
rect 7809 6301 7814 6357
rect 7870 6301 7875 6357
rect 7809 4577 7875 6301
rect 7809 4521 7814 4577
rect 7870 4521 7875 4577
rect 7809 2695 7875 4521
rect 7809 2639 7814 2695
rect 7870 2639 7875 2695
rect 7809 2629 7875 2639
rect 897 643 963 653
rect 897 587 902 643
rect 958 587 963 643
rect 897 -215 963 587
rect 897 -271 902 -215
rect 958 -271 963 -215
rect 897 -2875 963 -271
rect 2625 643 2691 653
rect 2625 587 2630 643
rect 2686 587 2691 643
rect 2625 -743 2691 587
rect 2625 -799 2630 -743
rect 2686 -799 2691 -743
rect 2625 -2347 2691 -799
rect 2625 -2403 2630 -2347
rect 2686 -2403 2691 -2347
rect 2625 -2413 2691 -2403
rect 4353 643 4419 653
rect 4353 587 4358 643
rect 4414 587 4419 643
rect 4353 -655 4419 587
rect 4353 -711 4358 -655
rect 4414 -711 4419 -655
rect 4353 -2435 4419 -711
rect 6081 643 6147 653
rect 6081 587 6086 643
rect 6142 587 6147 643
rect 6081 -1271 6147 587
rect 7809 643 7875 653
rect 7809 587 7814 643
rect 7870 587 7875 643
rect 7809 -1 7875 587
rect 6081 -1327 6086 -1271
rect 6142 -1327 6147 -1271
rect 6081 -1819 6147 -1327
rect 6081 -1875 6086 -1819
rect 6142 -1875 6147 -1819
rect 6081 -1880 6147 -1875
rect 7074 -67 7875 -1
rect 7074 -1183 7140 -67
rect 7074 -1239 7079 -1183
rect 7135 -1239 7140 -1183
rect 7074 -1907 7140 -1239
rect 7074 -1963 7079 -1907
rect 7135 -1963 7140 -1907
rect 7074 -1973 7140 -1963
rect 4353 -2491 4358 -2435
rect 4414 -2491 4419 -2435
rect 4353 -2501 4419 -2491
rect 897 -2931 902 -2875
rect 958 -2931 963 -2875
rect 897 -2941 963 -2931
use cm_head  cm_head_0
timestamp 1750075212
transform 1 0 434 0 1 7160
box -464 -3509 8900 2316
use cm_tail  cm_tail_0
timestamp 1750079478
transform 1 0 35 0 1 -5092
box -35 -39 7037 5101
use opa_diffpairs  opa_diffpairs_0
timestamp 1751017459
transform 1 0 33 0 1 316
box -63 -325 8797 3413
<< end >>
