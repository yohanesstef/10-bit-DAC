magic
tech sky130A
magscale 1 2
timestamp 1748936551
<< pwell >>
rect -307 -673 307 673
<< psubdiff >>
rect -271 603 -175 637
rect 175 603 271 637
rect -271 541 -237 603
rect 237 541 271 603
rect -271 -603 -237 -541
rect 237 -603 271 -541
rect -271 -637 -175 -603
rect 175 -637 271 -603
<< psubdiffcont >>
rect -175 603 175 637
rect -271 -541 -237 541
rect 237 -541 271 541
rect -175 -637 175 -603
<< xpolycontact >>
rect -141 75 141 507
rect -141 -507 141 -75
<< xpolyres >>
rect -141 -75 141 75
<< locali >>
rect -271 603 -175 637
rect 175 603 271 637
rect -271 541 -237 603
rect 237 541 271 603
rect -271 -603 -237 -541
rect 237 -603 271 -541
rect -271 -637 -175 -603
rect 175 -637 271 -603
<< viali >>
rect -125 92 125 489
rect -125 -489 125 -92
<< metal1 >>
rect -131 489 131 501
rect -131 92 -125 489
rect 125 92 131 489
rect -131 80 131 92
rect -131 -92 131 -80
rect -131 -489 -125 -92
rect 125 -489 131 -92
rect -131 -501 131 -489
<< properties >>
string FIXED_BBOX -254 -620 254 620
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 0.913 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 1.561k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
