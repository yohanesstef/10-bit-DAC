magic
tech sky130A
magscale 1 2
timestamp 1750156376
<< nwell >>
rect -4665 11508 4744 14208
<< mvnsubdiffcont >>
rect -4526 14095 4605 14129
rect -4586 12875 -4552 14069
rect 4631 12875 4665 14069
rect -4586 12841 4665 12875
rect -4586 11647 -4552 12841
rect 4631 11647 4665 12841
rect -4526 11587 4605 11621
<< viali >>
rect -4586 14095 -4526 14129
rect -4526 14095 4605 14129
rect 4605 14095 4665 14129
rect -4586 14069 -4552 14095
rect -4586 12875 -4552 14069
rect 4631 14069 4665 14095
rect 4631 12875 4665 14069
rect -4586 12841 4665 12875
rect -4586 11647 -4552 12841
rect -4586 11621 -4552 11647
rect 4631 11647 4665 12841
rect 4631 11621 4665 11647
rect -4586 11587 -4526 11621
rect -4526 11587 4605 11621
rect 4605 11587 4665 11621
<< via1 >>
rect 4530 12730 4590 12790
<< metal2 >>
rect 4530 12790 4590 12929
rect 4530 12724 4590 12730
use cm_pcell3_cell  cm_pcell3_cell_0
timestamp 1750156376
transform 1 0 -14 0 1 9178
box -4651 3584 4758 5030
use cm_pcell3_cell  cm_pcell3_cell_1
timestamp 1750156376
transform -1 0 93 0 1 7924
box -4651 3584 4758 5030
<< labels >>
flabel metal1 s -4511 13990 -4451 14050 0 FreeSans 320 0 0 0 VB1
port 0 nsew
flabel metal1 s 9 13603 69 13663 0 FreeSans 320 0 0 0 VB2
port 1 nsew
flabel metal1 s -4511 12261 -4451 12321 0 FreeSans 320 0 0 0 ROUT
port 2 nsew
flabel locali s -4586 14095 -4552 14129 0 FreeSans 320 0 0 0 VDDA
port 3 nsew
<< end >>
