magic
tech sky130A
magscale 1 2
timestamp 1750150351
<< metal2 >>
rect 1437 1791 1876 1851
rect 3165 1791 3604 1851
rect 4893 1791 5332 1851
rect 6621 1791 7060 1851
rect 8349 1791 8756 1851
rect 1844 1077 2139 1137
rect 3572 1077 3867 1137
rect 5300 1077 5595 1137
rect 7028 1077 7323 1137
rect 1844 957 2139 1017
rect 3572 957 3867 1017
rect 5300 957 5595 1017
rect 7028 957 7323 1017
rect 1437 155 1876 215
rect 3165 155 3604 215
rect 4893 155 5332 215
rect 6621 155 7060 215
rect 8349 155 8756 215
use dp_pmos  dp_pmos_0
timestamp 1750150351
transform 1 0 -35092 0 1 -19
box 35082 4 37002 2128
use dp_pmos  dp_pmos_1
timestamp 1750150351
transform 1 0 -33364 0 1 -19
box 35082 4 37002 2128
use dp_pmos  dp_pmos_2
timestamp 1750150351
transform 1 0 -29908 0 1 -19
box 35082 4 37002 2128
use dp_pmos  dp_pmos_3
timestamp 1750150351
transform 1 0 -31636 0 1 -19
box 35082 4 37002 2128
use dp_pmos  dp_pmos_5
timestamp 1750150351
transform 1 0 -28180 0 1 -19
box 35082 4 37002 2128
<< end >>
