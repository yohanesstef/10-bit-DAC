magic
tech sky130A
magscale 1 2
timestamp 1749550684
<< error_s >>
rect 31782 -7200 31788 -7194
rect 31836 -7200 31842 -7194
rect 31776 -7206 31782 -7200
rect 31842 -7206 31848 -7200
rect 31776 -7260 31782 -7254
rect 31842 -7260 31848 -7254
rect 31782 -7266 31788 -7260
rect 31836 -7266 31842 -7260
rect 31506 -7288 31512 -7282
rect 31560 -7288 31566 -7282
rect 31500 -7294 31506 -7288
rect 31566 -7294 31572 -7288
rect 31500 -7348 31506 -7342
rect 31566 -7348 31572 -7342
rect 31506 -7354 31512 -7348
rect 31560 -7354 31566 -7348
rect 31230 -7376 31236 -7370
rect 31284 -7376 31290 -7370
rect 31224 -7382 31230 -7376
rect 31290 -7382 31296 -7376
rect 31224 -7436 31230 -7430
rect 31290 -7436 31296 -7430
rect 31230 -7442 31236 -7436
rect 31284 -7442 31290 -7436
rect 30954 -7464 30960 -7458
rect 31008 -7464 31014 -7458
rect 30948 -7470 30954 -7464
rect 31014 -7470 31020 -7464
rect 30948 -7524 30954 -7518
rect 31014 -7524 31020 -7518
rect 30954 -7530 30960 -7524
rect 31008 -7530 31014 -7524
rect 30520 -7552 30526 -7546
rect 30574 -7552 30580 -7546
rect 30514 -7558 30520 -7552
rect 30580 -7558 30586 -7552
rect 30514 -7612 30520 -7606
rect 30580 -7612 30586 -7606
rect 30520 -7618 30526 -7612
rect 30574 -7618 30580 -7612
rect 30244 -7640 30250 -7634
rect 30298 -7640 30304 -7634
rect 30238 -7646 30244 -7640
rect 30304 -7646 30310 -7640
rect 30238 -7700 30244 -7694
rect 30304 -7700 30310 -7694
rect 30244 -7706 30250 -7700
rect 30298 -7706 30304 -7700
rect 29968 -7728 29974 -7722
rect 30022 -7728 30028 -7722
rect 29962 -7734 29968 -7728
rect 30028 -7734 30034 -7728
rect 29962 -7788 29968 -7782
rect 30028 -7788 30034 -7782
rect 29968 -7794 29974 -7788
rect 30022 -7794 30028 -7788
rect 29692 -7816 29698 -7810
rect 29746 -7816 29752 -7810
rect 29686 -7822 29692 -7816
rect 29752 -7822 29758 -7816
rect 29686 -7876 29692 -7870
rect 29752 -7876 29758 -7870
rect 29692 -7882 29698 -7876
rect 29746 -7882 29752 -7876
<< metal1 >>
rect 31782 -7200 31842 -7194
rect 31506 -7288 31566 -7282
rect 31230 -7376 31290 -7370
rect 30954 -7464 31014 -7458
rect 30520 -7552 30580 -7546
rect 30244 -7640 30304 -7634
rect 29968 -7728 30028 -7722
rect 29692 -7816 29752 -7810
rect 29692 -8000 29752 -7876
rect 29968 -8000 30028 -7788
rect 30244 -8000 30304 -7700
rect 30520 -8000 30580 -7612
rect 30954 -8000 31014 -7524
rect 31230 -8000 31290 -7436
rect 31506 -8000 31566 -7348
rect 31782 -8000 31842 -7260
rect 29875 -8378 29935 -8000
rect 30151 -8290 30211 -8000
rect 30427 -8202 30487 -8000
rect 30703 -8199 30753 -8000
rect 30427 -8262 30665 -8202
rect 30151 -8350 30577 -8290
rect 29875 -8438 30489 -8378
rect 30429 -9812 30489 -8438
rect 30517 -9812 30577 -8350
rect 30605 -9812 30665 -8262
rect 30693 -9812 30753 -8199
rect 30781 -8199 30831 -8000
rect 30781 -9812 30841 -8199
rect 31047 -8202 31107 -8000
rect 30869 -8262 31107 -8202
rect 30869 -9812 30929 -8262
rect 31323 -8290 31383 -8000
rect 30957 -8350 31383 -8290
rect 30957 -9812 31017 -8350
rect 31599 -8378 31659 -8000
rect 31045 -8438 31659 -8378
rect 31045 -9812 31105 -8438
<< via1 >>
rect 31782 -7260 31842 -7200
rect 31506 -7348 31566 -7288
rect 31230 -7436 31290 -7376
rect 30954 -7524 31014 -7464
rect 30520 -7612 30580 -7552
rect 30244 -7700 30304 -7640
rect 29968 -7788 30028 -7728
rect 29692 -7876 29752 -7816
use hnmos_8  hnmos_8_8
timestamp 1749548291
transform 1 0 29660 0 -1 -7984
box -137 -180 2351 358
<< end >>
