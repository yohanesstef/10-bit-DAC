magic
tech sky130A
magscale 1 2
timestamp 1750845293
<< pwell >>
rect -278 -749 278 749
<< mvnmos >>
rect -50 407 50 491
rect -50 167 50 251
rect -50 -73 50 11
rect -50 -313 50 -229
rect -50 -553 50 -469
<< mvndiff >>
rect -108 479 -50 491
rect -108 419 -96 479
rect -62 419 -50 479
rect -108 407 -50 419
rect 50 479 108 491
rect 50 419 62 479
rect 96 419 108 479
rect 50 407 108 419
rect -108 239 -50 251
rect -108 179 -96 239
rect -62 179 -50 239
rect -108 167 -50 179
rect 50 239 108 251
rect 50 179 62 239
rect 96 179 108 239
rect 50 167 108 179
rect -108 -1 -50 11
rect -108 -61 -96 -1
rect -62 -61 -50 -1
rect -108 -73 -50 -61
rect 50 -1 108 11
rect 50 -61 62 -1
rect 96 -61 108 -1
rect 50 -73 108 -61
rect -108 -241 -50 -229
rect -108 -301 -96 -241
rect -62 -301 -50 -241
rect -108 -313 -50 -301
rect 50 -241 108 -229
rect 50 -301 62 -241
rect 96 -301 108 -241
rect 50 -313 108 -301
rect -108 -481 -50 -469
rect -108 -541 -96 -481
rect -62 -541 -50 -481
rect -108 -553 -50 -541
rect 50 -481 108 -469
rect 50 -541 62 -481
rect 96 -541 108 -481
rect 50 -553 108 -541
<< mvndiffc >>
rect -96 419 -62 479
rect 62 419 96 479
rect -96 179 -62 239
rect 62 179 96 239
rect -96 -61 -62 -1
rect 62 -61 96 -1
rect -96 -301 -62 -241
rect 62 -301 96 -241
rect -96 -541 -62 -481
rect 62 -541 96 -481
<< mvpsubdiff >>
rect -242 701 242 713
rect -242 667 -134 701
rect 134 667 242 701
rect -242 655 242 667
rect -242 605 -184 655
rect -242 -605 -230 605
rect -196 -605 -184 605
rect 184 605 242 655
rect -242 -655 -184 -605
rect 184 -605 196 605
rect 230 -605 242 605
rect 184 -655 242 -605
rect -242 -667 242 -655
rect -242 -701 -134 -667
rect 134 -701 242 -667
rect -242 -713 242 -701
<< mvpsubdiffcont >>
rect -134 667 134 701
rect -230 -605 -196 605
rect 196 -605 230 605
rect -134 -701 134 -667
<< poly >>
rect -50 563 50 579
rect -50 529 -34 563
rect 34 529 50 563
rect -50 491 50 529
rect -50 381 50 407
rect -50 323 50 339
rect -50 289 -34 323
rect 34 289 50 323
rect -50 251 50 289
rect -50 141 50 167
rect -50 83 50 99
rect -50 49 -34 83
rect 34 49 50 83
rect -50 11 50 49
rect -50 -99 50 -73
rect -50 -157 50 -141
rect -50 -191 -34 -157
rect 34 -191 50 -157
rect -50 -229 50 -191
rect -50 -339 50 -313
rect -50 -397 50 -381
rect -50 -431 -34 -397
rect 34 -431 50 -397
rect -50 -469 50 -431
rect -50 -579 50 -553
<< polycont >>
rect -34 529 34 563
rect -34 289 34 323
rect -34 49 34 83
rect -34 -191 34 -157
rect -34 -431 34 -397
<< locali >>
rect -230 667 -134 701
rect 134 667 230 701
rect -230 605 -196 667
rect 196 605 230 667
rect -50 529 -34 563
rect 34 529 50 563
rect -96 479 -62 495
rect -96 403 -62 419
rect 62 479 96 495
rect 62 403 96 419
rect -50 289 -34 323
rect 34 289 50 323
rect -96 239 -62 255
rect -96 163 -62 179
rect 62 239 96 255
rect 62 163 96 179
rect -50 49 -34 83
rect 34 49 50 83
rect -96 -1 -62 15
rect -96 -77 -62 -61
rect 62 -1 96 15
rect 62 -77 96 -61
rect -50 -191 -34 -157
rect 34 -191 50 -157
rect -96 -241 -62 -225
rect -96 -317 -62 -301
rect 62 -241 96 -225
rect 62 -317 96 -301
rect -50 -431 -34 -397
rect 34 -431 50 -397
rect -96 -481 -62 -465
rect -96 -557 -62 -541
rect 62 -481 96 -465
rect 62 -557 96 -541
rect -230 -667 -196 -605
rect 196 -667 230 -605
rect -230 -701 -134 -667
rect 134 -701 230 -667
<< viali >>
rect -26 529 26 563
rect -96 419 -62 479
rect 62 419 96 479
rect -26 289 26 323
rect -96 179 -62 239
rect 62 179 96 239
rect -26 49 26 83
rect -96 -61 -62 -1
rect 62 -61 96 -1
rect -26 -191 26 -157
rect -96 -301 -62 -241
rect 62 -301 96 -241
rect -26 -431 26 -397
rect -96 -541 -62 -481
rect 62 -541 96 -481
<< metal1 >>
rect -38 563 38 569
rect -38 529 -26 563
rect 26 529 38 563
rect -38 523 38 529
rect -102 479 -56 491
rect -102 419 -96 479
rect -62 419 -56 479
rect -102 407 -56 419
rect 56 479 102 491
rect 56 419 62 479
rect 96 419 102 479
rect 56 407 102 419
rect -38 323 38 329
rect -38 289 -26 323
rect 26 289 38 323
rect -38 283 38 289
rect -102 239 -56 251
rect -102 179 -96 239
rect -62 179 -56 239
rect -102 167 -56 179
rect 56 239 102 251
rect 56 179 62 239
rect 96 179 102 239
rect 56 167 102 179
rect -38 83 38 89
rect -38 49 -26 83
rect 26 49 38 83
rect -38 43 38 49
rect -102 -1 -56 11
rect -102 -61 -96 -1
rect -62 -61 -56 -1
rect -102 -73 -56 -61
rect 56 -1 102 11
rect 56 -61 62 -1
rect 96 -61 102 -1
rect 56 -73 102 -61
rect -38 -157 38 -151
rect -38 -191 -26 -157
rect 26 -191 38 -157
rect -38 -197 38 -191
rect -102 -241 -56 -229
rect -102 -301 -96 -241
rect -62 -301 -56 -241
rect -102 -313 -56 -301
rect 56 -241 102 -229
rect 56 -301 62 -241
rect 96 -301 102 -241
rect 56 -313 102 -301
rect -38 -397 38 -391
rect -38 -431 -26 -397
rect 26 -431 38 -397
rect -38 -437 38 -431
rect -102 -481 -56 -469
rect -102 -541 -96 -481
rect -62 -541 -56 -481
rect -102 -553 -56 -541
rect 56 -481 102 -469
rect 56 -541 62 -481
rect 96 -541 102 -481
rect 56 -553 102 -541
<< properties >>
string FIXED_BBOX -213 -684 213 684
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.420 l 0.50 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
