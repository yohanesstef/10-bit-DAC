magic
tech sky130A
magscale 1 2
timestamp 1750150351
<< pwell >>
rect 1143 1631 2701 1666
<< mvpsubdiff >>
rect 1143 1631 2701 1666
<< locali >>
rect 1156 1618 2688 1679
<< metal1 >>
rect 2371 1917 2431 2368
rect 2371 1851 2431 1857
rect 685 1449 745 1455
rect 685 1383 745 1389
rect 773 1449 833 1455
rect 773 1383 833 1389
<< via1 >>
rect 2371 1857 2431 1917
rect 685 1389 745 1449
rect 773 1389 833 1449
<< metal2 >>
rect 2371 1917 2431 1923
rect 685 1857 1319 1917
rect 685 1449 745 1857
rect 685 1383 745 1389
rect 773 1769 1319 1829
rect 773 1449 833 1769
rect 2371 1741 2431 1857
rect 1892 1681 2431 1741
rect 1892 1640 1952 1681
rect 773 1383 833 1389
use fc_ncell1  fc_ncell1_0
timestamp 1750150351
transform 1 0 451 0 1 1103
box 94 -748 2848 564
use fc_ncell2  fc_ncell2_0
timestamp 1750150351
transform 1 0 1152 0 1 2476
box -45 -846 1585 816
<< end >>
