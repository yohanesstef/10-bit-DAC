magic
tech sky130A
magscale 1 2
timestamp 1750203392
<< mvpsubdiff >>
rect 1805 1925 3273 1985
rect 1805 1612 1865 1925
rect 3213 1612 3273 1925
rect 1805 1552 3273 1612
<< poly >>
rect 1876 1660 1936 1894
rect 3142 1660 3202 1894
<< locali >>
rect 1818 1938 3260 1972
rect 1818 1599 1852 1938
rect 3226 1599 3260 1938
rect 1818 1565 3260 1599
rect 1818 1564 1875 1565
<< metal1 >>
rect 1795 1915 3283 1995
rect 1795 1622 1875 1915
rect 3075 1622 3121 1686
rect 3203 1622 3283 1915
rect 1795 1542 3283 1622
use sky130_fd_pr__nfet_g5v0d10v5_SZ2N2S  sky130_fd_pr__nfet_g5v0d10v5_SZ2N2S_0
timestamp 1750202493
transform 1 0 2539 0 1 1777
box -588 -117 588 117
<< end >>
