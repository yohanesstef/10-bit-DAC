magic
tech sky130A
magscale 1 2
timestamp 1749890363
<< error_s >>
rect 6050 2542 6056 2548
rect 6104 2542 6110 2548
rect 7554 2542 7560 2548
rect 7608 2542 7614 2548
rect 6044 2536 6050 2542
rect 6110 2536 6116 2542
rect 7548 2536 7554 2542
rect 7614 2536 7620 2542
rect 6044 2482 6050 2488
rect 6110 2482 6116 2488
rect 7548 2482 7554 2488
rect 7614 2482 7620 2488
rect 6050 2476 6056 2482
rect 6104 2476 6110 2482
rect 7554 2476 7560 2482
rect 7608 2476 7614 2482
rect 5298 2454 5304 2460
rect 5352 2454 5358 2460
rect 6802 2454 6808 2460
rect 6856 2454 6862 2460
rect 8306 2454 8312 2460
rect 8360 2454 8366 2460
rect 5292 2448 5298 2454
rect 5358 2448 5364 2454
rect 6796 2448 6802 2454
rect 6862 2448 6868 2454
rect 8300 2448 8306 2454
rect 8366 2448 8372 2454
rect 5292 2394 5298 2400
rect 5358 2394 5364 2400
rect 6796 2394 6802 2400
rect 6862 2394 6868 2400
rect 8300 2394 8306 2400
rect 8366 2394 8372 2400
rect 5298 2388 5304 2394
rect 5352 2388 5358 2394
rect 6802 2388 6808 2394
rect 6856 2388 6862 2394
rect 8306 2388 8312 2394
rect 8360 2388 8366 2394
rect 7930 2190 7936 2196
rect 7984 2190 7990 2196
rect 7924 2184 7930 2190
rect 7990 2184 7996 2190
rect 7924 2130 7930 2136
rect 7990 2130 7996 2136
rect 7930 2124 7936 2130
rect 7984 2124 7990 2130
rect 7178 2102 7184 2108
rect 7232 2102 7238 2108
rect 8623 2102 8629 2108
rect 8677 2102 8683 2108
rect 7172 2096 7178 2102
rect 7238 2096 7244 2102
rect 8617 2096 8623 2102
rect 8683 2096 8689 2102
rect 7172 2042 7178 2048
rect 7238 2042 7244 2048
rect 8617 2042 8623 2048
rect 8683 2042 8689 2048
rect 7178 2036 7184 2042
rect 7232 2036 7238 2042
rect 8623 2036 8629 2042
rect 8677 2036 8683 2042
rect 6426 2014 6432 2020
rect 6480 2014 6486 2020
rect 6420 2008 6426 2014
rect 6486 2008 6492 2014
rect 6420 1954 6426 1960
rect 6486 1954 6492 1960
rect 6426 1948 6432 1954
rect 6480 1948 6486 1954
rect 5674 1926 5680 1932
rect 5728 1926 5734 1932
rect 5668 1920 5674 1926
rect 5734 1920 5740 1926
rect 5668 1866 5674 1872
rect 5734 1866 5740 1872
rect 5674 1860 5680 1866
rect 5728 1860 5734 1866
<< metal1 >>
rect 8623 2102 8683 2108
rect 8623 2036 8683 2042
<< via1 >>
rect 6050 2482 6110 2542
rect 7554 2482 7614 2542
rect 5298 2394 5358 2454
rect 6802 2394 6862 2454
rect 8306 2394 8366 2454
rect 7930 2130 7990 2190
rect 7178 2042 7238 2102
rect 8623 2042 8683 2102
rect 6426 1954 6486 2014
rect 5674 1866 5734 1926
use cm_pcell1_cell  cm_pcell1_cell_0
timestamp 1749890363
transform 1 0 4905 0 1 1555
box -35 -10 4729 1308
<< end >>
