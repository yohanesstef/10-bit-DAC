magic
tech sky130A
magscale 1 2
timestamp 1749890363
<< metal1 >>
rect 325 -392 489 -317
rect 701 -392 865 -317
rect 1077 -392 1241 -317
rect 1453 -392 1611 -317
use cm_pcell1_4  cm_pcell1_4_0
timestamp 1749890363
transform 1 0 -14 0 1 -323
box -21 1 1625 678
use cm_pcell1_4  cm_pcell1_4_1
timestamp 1749890363
transform 1 0 -14 0 -1 -283
box -21 1 1625 678
<< end >>
