magic
tech sky130A
magscale 1 2
timestamp 1749147130
<< pwell >>
rect -307 -822 307 822
<< psubdiff >>
rect -271 752 -175 786
rect 175 752 271 786
rect -271 690 -237 752
rect 237 690 271 752
rect -271 -752 -237 -690
rect 237 -752 271 -690
rect -271 -786 -175 -752
rect 175 -786 271 -752
<< psubdiffcont >>
rect -175 752 175 786
rect -271 -690 -237 690
rect 237 -690 271 690
rect -175 -786 175 -752
<< xpolycontact >>
rect -141 224 141 656
rect -141 -656 141 -224
<< xpolyres >>
rect -141 -224 141 224
<< locali >>
rect -271 752 -175 786
rect 175 752 271 786
rect -271 690 -237 752
rect 237 690 271 752
rect -271 -752 -237 -690
rect 237 -752 271 -690
rect -271 -786 -175 -752
rect 175 -786 271 -752
<< viali >>
rect -125 241 125 638
rect -125 -638 125 -241
<< metal1 >>
rect -131 638 131 650
rect -131 241 -125 638
rect 125 241 131 638
rect -131 229 131 241
rect -131 -241 131 -229
rect -131 -638 -125 -241
rect 125 -638 131 -241
rect -131 -650 131 -638
<< properties >>
string FIXED_BBOX -254 -769 254 769
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 2.399 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 3.669k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
