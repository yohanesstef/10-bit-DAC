magic
tech sky130A
magscale 1 2
timestamp 1749538868
<< metal1 >>
rect 18462 -23125 18522 -21181
rect 18550 -22477 18610 -21181
rect 18638 -21829 18698 -21181
rect 18726 -21443 18731 -21181
rect 18731 -21505 19147 -21443
rect 19701 -21505 19761 -21181
rect 19678 -21767 19761 -21505
rect 19257 -21829 19678 -21767
rect 18638 -22091 18726 -21829
rect 18726 -22153 19147 -22091
rect 19789 -22153 19849 -21181
rect 19678 -22415 19849 -22153
rect 19257 -22477 19678 -22415
rect 18550 -22739 18726 -22477
rect 18726 -22801 19147 -22739
rect 19877 -22801 19937 -21181
rect 19678 -23063 19937 -22801
rect 19257 -23125 19678 -23063
rect 18462 -23387 18726 -23125
rect 18726 -23449 19142 -23387
use sky130_fd_pr__res_xhigh_po_1p41_238JSU  sky130_fd_pr__res_xhigh_po_1p41_238JSU_0
timestamp 1749123380
transform 0 -1 19202 1 0 -23904
box -141 -487 141 487
use sky130_fd_pr__res_xhigh_po_1p41_238LSU  sky130_fd_pr__res_xhigh_po_1p41_238LSU_0
timestamp 1748944356
transform 0 -1 19202 1 0 -23580
box -141 -487 141 487
use sky130_fd_pr__res_xhigh_po_1p41_C5Z94V  sky130_fd_pr__res_xhigh_po_1p41_C5Z94V_0
timestamp 1748944356
transform 0 -1 19202 1 0 -21636
box -141 -482 141 482
use sky130_fd_pr__res_xhigh_po_1p41_HUJR2Q  sky130_fd_pr__res_xhigh_po_1p41_HUJR2Q_0
timestamp 1749201400
transform 0 -1 19202 1 0 -20988
box -141 -477 141 477
use sky130_fd_pr__res_xhigh_po_1p41_C5Z94V  XR58
timestamp 1748944356
transform 0 -1 19202 1 0 -23256
box -141 -482 141 482
use sky130_fd_pr__res_xhigh_po_1p41_C5Z94V  XR59
timestamp 1748944356
transform 0 -1 19202 1 0 -22932
box -141 -482 141 482
use sky130_fd_pr__res_xhigh_po_1p41_C5Z94V  XR60
timestamp 1748944356
transform 0 -1 19202 1 0 -22608
box -141 -482 141 482
use sky130_fd_pr__res_xhigh_po_1p41_C5Z94V  XR61
timestamp 1748944356
transform 0 -1 19202 1 0 -22284
box -141 -482 141 482
use sky130_fd_pr__res_xhigh_po_1p41_C5Z94V  XR62
timestamp 1748944356
transform 0 -1 19202 1 0 -21960
box -141 -482 141 482
use sky130_fd_pr__res_xhigh_po_1p41_HUJT2Q  XR64
timestamp 1748944356
transform 0 -1 19202 1 0 -21312
box -141 -477 141 477
<< end >>
