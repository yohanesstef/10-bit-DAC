magic
tech sky130A
magscale 1 2
timestamp 1750771847
<< pwell >>
rect -56 -638 1418 626
<< metal1 >>
rect 84 398 144 492
rect 84 -438 144 338
rect 84 -504 144 -498
rect 172 486 232 492
rect 172 -350 232 426
rect 599 398 645 486
rect 704 426 710 486
rect 770 426 776 486
rect 586 338 592 398
rect 652 338 658 398
rect 599 232 645 338
rect 717 232 763 426
rect 341 84 387 112
rect 975 84 1021 112
rect 341 24 537 84
rect 826 24 955 84
rect 1015 24 1021 84
rect 341 -96 537 -36
rect 826 -96 955 -36
rect 1015 -96 1021 -36
rect 341 -124 387 -96
rect 975 -124 1021 -96
rect 599 -350 645 -244
rect 586 -410 592 -350
rect 652 -410 658 -350
rect 172 -504 232 -410
rect 599 -498 645 -410
rect 717 -438 763 -239
rect 704 -498 710 -438
rect 770 -498 776 -438
<< via1 >>
rect 84 338 144 398
rect 84 -498 144 -438
rect 172 426 232 486
rect 710 426 770 486
rect 592 338 652 398
rect 955 24 1015 84
rect 955 -96 1015 -36
rect 172 -410 232 -350
rect 592 -410 652 -350
rect 710 -498 770 -438
<< metal2 >>
rect 78 426 172 486
rect 232 426 710 486
rect 770 426 776 486
rect 78 338 84 398
rect 144 338 592 398
rect 652 338 776 398
rect 949 24 955 84
rect 1015 24 1284 84
rect 949 -96 955 -36
rect 1015 -96 1284 -36
rect 78 -410 172 -350
rect 232 -410 592 -350
rect 652 -410 776 -350
rect 78 -498 84 -438
rect 144 -498 710 -438
rect 770 -498 776 -438
use cm2_ncell2_ncell  cm2_ncell2_ncell_0
timestamp 1750771847
transform 1 0 -1062 0 1 -181
box 1032 175 2454 781
use cm2_ncell2_ncell  cm2_ncell2_ncell_1
timestamp 1750771847
transform -1 0 2424 0 -1 169
box 1032 175 2454 781
use cross_pair  cross_pair_0
timestamp 1750150351
transform 1 0 -35577 0 1 -1951
box 36114 1855 36403 2035
<< end >>
