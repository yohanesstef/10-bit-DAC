* PEX produced on Tue Jun 24 20:55:49 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from top_bias_lvsf_dec.ext - technology: sky130A

.subckt bias_lvsf_posim ROUT VBPLV VBNLV VBPDEC VBNDEC VDDA GNDA
X0 cm2_pcell_0.cm2_pcell2_0.S4.t3 cm2_pcell_0.cm2_pcell2_0.S0.t6 VDDA.t45 VDDA.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X1 cm2_pcell_0.cm2_pcell2_0.S2.t1 cm2_pcell_0.D0.t6 VBPDEC.t4 VDDA.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X2 VBNDEC.t5 cm2_pcell_0.D0.t7 cm2_pcell_0.cm2_pcell2_0.S4.t1 VDDA.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X3 GNDA.t8 a_4080_n2791.t3 a_4080_n2791.t4 GNDA.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X4 cm2_pcell_0.cm2_pcell2_0.S0.t4 cm2_pcell_0.cm2_pcell2_0.S0.t3 VDDA.t44 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X5 VBPDEC.t1 VBPDEC.t0 a_4602_n3479.t1 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X6 a_11186_n55.t3 ROUT.t4 cm2_pcell_0.D0.t5 VDDA.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X7 cm2_pcell_0.D1.t3 cm2_pcell_0.D1.t2 a_4080_n2791.t0 GNDA.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X8 VDDA.t34 VDDA.t32 VDDA.t33 VDDA.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X9 VDDA.t43 cm2_pcell_0.cm2_pcell2_0.S0.t1 cm2_pcell_0.cm2_pcell2_0.S0.t2 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X10 cm2_pcell_0.cm2_pcell2_0.S4.t0 cm2_pcell_0.D0.t8 VBNDEC.t4 VDDA.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X11 VBPDEC.t5 cm2_pcell_0.D0.t9 cm2_pcell_0.cm2_pcell2_0.S2.t0 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X12 VDDA.t31 VDDA.t29 VDDA.t30 VDDA.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X13 VBPLV.t1 cm2_pcell_0.D1.t6 a_4080_n3027.t1 GNDA.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X14 a_6498_n2100.t2 VBNLV.t2 VBNLV.t3 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X15 a_6498_n2100.t0 VBNLV.t6 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=5.3
X16 a_11186_n55.t1 ROUT.t2 ROUT.t3 VDDA.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X17 a_5864_n2100.t0 VBNDEC.t6 GNDA.t15 GNDA.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1769 pd=1.8 as=0.1769 ps=1.8 w=0.61 l=9.7
X18 cm2_pcell_0.cm2_pcell2_0.S3.t3 cm2_pcell_0.cm2_pcell2_0.S0.t7 VDDA.t42 VDDA.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X19 a_4080_n3027.t3 a_4080_n2791.t6 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X20 GNDA.t5 a_4080_n2791.t7 a_4080_n3027.t2 GNDA.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X21 VDDA.t28 VDDA.t26 VDDA.t27 VDDA.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X22 cm2_pcell_0.D0.t4 cm2_pcell_0.D0.t3 cm2_pcell_0.cm2_pcell2_0.S0.t5 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X23 VDDA.t25 VDDA.t23 VDDA.t24 VDDA.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X24 cm2_pcell_0.cm2_pcell2_0.S1.t1 cm2_pcell_0.D0.t10 cm2_pcell_0.D1.t5 VDDA.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X25 VBNLV.t4 cm2_pcell_0.D0.t11 cm2_pcell_0.cm2_pcell2_0.S3.t1 VDDA.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X26 cm2_pcell_0.cm2_pcell2_0.S2.t3 cm2_pcell_0.cm2_pcell2_0.S0.t8 VDDA.t41 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X27 a_5864_n2100.t2 VBNDEC.t2 VBNDEC.t3 GNDA.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X28 VDDA.t40 cm2_pcell_0.cm2_pcell2_0.S0.t9 cm2_pcell_0.cm2_pcell2_0.S4.t2 VDDA.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X29 VBNDEC.t1 VBNDEC.t0 a_5864_n2100.t1 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X30 VDDA.t6 VBPLV.t6 a_7128_n494.t2 VDDA.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9.2
X31 a_11186_n55.t0 ROUT.t0 ROUT.t1 VDDA.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X32 a_7128_n494.t1 VBPLV.t2 VBPLV.t3 VDDA.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=1
X33 VDDA.t39 cm2_pcell_0.cm2_pcell2_0.S0.t10 cm2_pcell_0.cm2_pcell2_0.S2.t2 VDDA.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X34 VDDA.t22 VDDA.t20 VDDA.t21 VDDA.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X35 a_6498_n2100.t1 VBNLV.t0 VBNLV.t1 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X36 a_4080_n2791.t2 a_4080_n2791.t1 GNDA.t4 GNDA.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X37 VDDA.t19 VDDA.t17 VDDA.t18 VDDA.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X38 VDDA.t38 cm2_pcell_0.cm2_pcell2_0.S0.t11 cm2_pcell_0.cm2_pcell2_0.S1.t3 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X39 cm2_pcell_0.cm2_pcell2_0.S3.t0 cm2_pcell_0.D0.t12 VBNLV.t5 VDDA.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X40 cm2_pcell_0.D1.t4 cm2_pcell_0.D0.t13 cm2_pcell_0.cm2_pcell2_0.S1.t0 VDDA.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X41 VDDA.t37 cm2_pcell_0.cm2_pcell2_0.S0.t12 cm2_pcell_0.cm2_pcell2_0.S3.t2 VDDA.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X42 VDDA.t16 VDDA.t13 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X43 a_4080_n3027.t0 cm2_pcell_0.D1.t7 VBPLV.t0 GNDA.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X44 cm2_pcell_0.cm2_pcell2_0.S1.t2 cm2_pcell_0.cm2_pcell2_0.S0.t13 VDDA.t36 VDDA.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X45 cm2_pcell_0.D0.t2 cm2_pcell_0.D0.t1 cm2_pcell_0.cm2_pcell2_0.S0.t0 VDDA.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X46 VDDA.t12 VDDA.t9 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X47 a_4080_n2791.t5 cm2_pcell_0.D1.t0 cm2_pcell_0.D1.t1 GNDA.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X48 VBPLV.t5 VBPLV.t4 a_7128_n494.t0 VDDA.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=1
X49 a_4602_n3479.t3 a_4602_n3479.t2 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1856 pd=1.86 as=0.1856 ps=1.86 w=0.64 l=12
X50 a_11186_n55.t2 ROUT.t5 cm2_pcell_0.D0.t0 VDDA.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X51 a_4602_n3479.t0 VBPDEC.t2 VBPDEC.t3 GNDA.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
R0 cm2_pcell_0.cm2_pcell2_0.S0.n6 cm2_pcell_0.cm2_pcell2_0.S0.t7 142.488
R1 cm2_pcell_0.cm2_pcell2_0.S0.n5 cm2_pcell_0.cm2_pcell2_0.S0.t6 142.488
R2 cm2_pcell_0.cm2_pcell2_0.S0.n2 cm2_pcell_0.cm2_pcell2_0.S0.t9 142.488
R3 cm2_pcell_0.cm2_pcell2_0.S0.n1 cm2_pcell_0.cm2_pcell2_0.S0.t12 142.488
R4 cm2_pcell_0.cm2_pcell2_0.S0.n6 cm2_pcell_0.cm2_pcell2_0.S0.t11 141.704
R5 cm2_pcell_0.cm2_pcell2_0.S0.n5 cm2_pcell_0.cm2_pcell2_0.S0.t10 141.704
R6 cm2_pcell_0.cm2_pcell2_0.S0.n2 cm2_pcell_0.cm2_pcell2_0.S0.t8 141.704
R7 cm2_pcell_0.cm2_pcell2_0.S0.n1 cm2_pcell_0.cm2_pcell2_0.S0.t13 141.704
R8 cm2_pcell_0.cm2_pcell2_0.S0.n8 cm2_pcell_0.cm2_pcell2_0.S0.t3 139.454
R9 cm2_pcell_0.cm2_pcell2_0.S0.n4 cm2_pcell_0.cm2_pcell2_0.S0.t1 139.454
R10 cm2_pcell_0.cm2_pcell2_0.S0.n12 cm2_pcell_0.cm2_pcell2_0.S0.t0 135.305
R11 cm2_pcell_0.cm2_pcell2_0.S0.n0 cm2_pcell_0.cm2_pcell2_0.S0.t4 135.246
R12 cm2_pcell_0.cm2_pcell2_0.S0.n10 cm2_pcell_0.cm2_pcell2_0.S0.t2 135.246
R13 cm2_pcell_0.cm2_pcell2_0.S0 cm2_pcell_0.cm2_pcell2_0.S0.t5 135.244
R14 cm2_pcell_0.cm2_pcell2_0.S0.n12 cm2_pcell_0.cm2_pcell2_0.S0.n11 12.38
R15 cm2_pcell_0.cm2_pcell2_0.S0.n11 cm2_pcell_0.cm2_pcell2_0.S0.n0 5.038
R16 cm2_pcell_0.cm2_pcell2_0.S0.n11 cm2_pcell_0.cm2_pcell2_0.S0.n10 4.5005
R17 cm2_pcell_0.cm2_pcell2_0.S0.n8 cm2_pcell_0.cm2_pcell2_0.S0.n7 2.2505
R18 cm2_pcell_0.cm2_pcell2_0.S0.n4 cm2_pcell_0.cm2_pcell2_0.S0.n3 2.2505
R19 cm2_pcell_0.cm2_pcell2_0.S0.n9 cm2_pcell_0.cm2_pcell2_0.S0.n4 0.842167
R20 cm2_pcell_0.cm2_pcell2_0.S0.n9 cm2_pcell_0.cm2_pcell2_0.S0.n8 0.842167
R21 cm2_pcell_0.cm2_pcell2_0.S0.n7 cm2_pcell_0.cm2_pcell2_0.S0.n5 0.783833
R22 cm2_pcell_0.cm2_pcell2_0.S0.n7 cm2_pcell_0.cm2_pcell2_0.S0.n6 0.783833
R23 cm2_pcell_0.cm2_pcell2_0.S0.n3 cm2_pcell_0.cm2_pcell2_0.S0.n1 0.783833
R24 cm2_pcell_0.cm2_pcell2_0.S0.n3 cm2_pcell_0.cm2_pcell2_0.S0.n2 0.783833
R25 cm2_pcell_0.cm2_pcell2_0.S0.n9 cm2_pcell_0.cm2_pcell2_0.S0.n0 0.26925
R26 cm2_pcell_0.cm2_pcell2_0.S0.n10 cm2_pcell_0.cm2_pcell2_0.S0.n9 0.26925
R27 cm2_pcell_0.cm2_pcell2_0.S0 cm2_pcell_0.cm2_pcell2_0.S0.n12 0.063
R28 VDDA.n51 VDDA.n50 5941.3
R29 VDDA.n7 VDDA.n3 5939.4
R30 VDDA.n50 VDDA.n9 3072.35
R31 VDDA.n46 VDDA.n9 2375.56
R32 VDDA.n63 VDDA.n62 1349.17
R33 VDDA.n52 VDDA.n2 1182.12
R34 VDDA.n52 VDDA.n1 1182.12
R35 VDDA.n60 VDDA.n2 1181.74
R36 VDDA.n63 VDDA.n0 739.817
R37 VDDA.n61 VDDA.n0 718.591
R38 VDDA.n9 VDDA.n3 672.484
R39 VDDA.n62 VDDA.n61 383.473
R40 VDDA.n62 VDDA.n1 366.202
R41 VDDA.n55 VDDA.t6 227.737
R42 VDDA.n8 VDDA.n7 177.855
R43 VDDA.t14 VDDA.n46 162.96
R44 VDDA.n23 VDDA.t17 139.454
R45 VDDA.n11 VDDA.t13 139.454
R46 VDDA.n16 VDDA.t20 139.454
R47 VDDA.n18 VDDA.t9 139.454
R48 VDDA.n29 VDDA.t29 139.454
R49 VDDA.n34 VDDA.t32 139.454
R50 VDDA.n37 VDDA.t23 139.454
R51 VDDA.n40 VDDA.t26 139.454
R52 VDDA.n10 VDDA.t15 135.312
R53 VDDA.n10 VDDA.t16 135.312
R54 VDDA.n24 VDDA.t19 135.312
R55 VDDA.n15 VDDA.t22 135.312
R56 VDDA.n15 VDDA.t21 135.312
R57 VDDA.n17 VDDA.t11 135.312
R58 VDDA.n17 VDDA.t12 135.312
R59 VDDA.n35 VDDA.t34 135.312
R60 VDDA.n33 VDDA.t33 135.312
R61 VDDA.n28 VDDA.t30 135.312
R62 VDDA.n36 VDDA.t25 135.312
R63 VDDA.n36 VDDA.t24 135.312
R64 VDDA.n39 VDDA.t28 135.312
R65 VDDA.n39 VDDA.t27 135.312
R66 VDDA.n12 VDDA.t18 134.712
R67 VDDA.n12 VDDA.t42 134.712
R68 VDDA.n13 VDDA.t38 134.712
R69 VDDA.n13 VDDA.t44 134.712
R70 VDDA.n14 VDDA.t39 134.712
R71 VDDA.n14 VDDA.t45 134.712
R72 VDDA.n27 VDDA.t37 134.712
R73 VDDA.n27 VDDA.t31 134.712
R74 VDDA.n25 VDDA.t40 134.712
R75 VDDA.n25 VDDA.t41 134.712
R76 VDDA.n26 VDDA.t43 134.712
R77 VDDA.n26 VDDA.t36 134.712
R78 VDDA.n47 VDDA.t10 119.24
R79 VDDA.t10 VDDA.t4 113.218
R80 VDDA.t4 VDDA.t35 113.218
R81 VDDA.t35 VDDA.t7 113.218
R82 VDDA.t7 VDDA.t8 113.218
R83 VDDA.t8 VDDA.t2 113.218
R84 VDDA.t2 VDDA.t14 113.218
R85 VDDA.n48 VDDA.t1 111.41
R86 VDDA.n46 VDDA.n45 92.5005
R87 VDDA.n49 VDDA.t3 86.5389
R88 VDDA.n49 VDDA.t5 83.5887
R89 VDDA.t0 VDDA.n47 82.5045
R90 VDDA.t1 VDDA.t0 77.6867
R91 VDDA.t5 VDDA.n48 57.8135
R92 VDDA.n61 VDDA.n60 54.2123
R93 VDDA.n50 VDDA.n49 49.5835
R94 VDDA.n51 VDDA.n8 33.4588
R95 VDDA.n60 VDDA.n3 6.85235
R96 VDDA.n47 VDDA.n3 6.85235
R97 VDDA.n52 VDDA.n51 6.85235
R98 VDDA.n48 VDDA.t3 6.73471
R99 VDDA VDDA.n63 6.4005
R100 VDDA.n53 VDDA.n4 4.87081
R101 VDDA.n54 VDDA.n53 4.87081
R102 VDDA.n59 VDDA.n4 4.86925
R103 VDDA.n45 VDDA.n44 4.6505
R104 VDDA.n57 VDDA.n56 3.41925
R105 VDDA.n42 VDDA.n41 3.13175
R106 VDDA.n41 VDDA.n38 3.0505
R107 VDDA.n7 VDDA.n2 2.93701
R108 VDDA.n50 VDDA.n1 2.93701
R109 VDDA.n55 VDDA.n6 2.5573
R110 VDDA.n43 VDDA.n35 1.79104
R111 VDDA.n28 VDDA.n5 1.79104
R112 VDDA.n58 VDDA.n57 1.12706
R113 VDDA.n45 VDDA.n0 1.07517
R114 VDDA.t3 VDDA.n8 1.0395
R115 VDDA.n22 VDDA.n21 0.985808
R116 VDDA.n31 VDDA.n30 0.947451
R117 VDDA.n21 VDDA.n20 0.91925
R118 VDDA.n32 VDDA.n31 0.91925
R119 VDDA.n57 VDDA.n6 0.806458
R120 VDDA.n38 VDDA.n6 0.789247
R121 VDDA.n56 VDDA.n55 0.788
R122 VDDA.n33 VDDA.n32 0.534794
R123 VDDA.n20 VDDA.n19 0.516125
R124 VDDA.n53 VDDA.n52 0.358192
R125 VDDA.n60 VDDA.n59 0.358192
R126 VDDA.n21 VDDA.n13 0.255835
R127 VDDA.n20 VDDA.n14 0.255835
R128 VDDA.n32 VDDA.n25 0.255835
R129 VDDA.n31 VDDA.n26 0.255835
R130 VDDA.n58 VDDA.n5 0.241125
R131 VDDA.n43 VDDA.n42 0.241125
R132 VDDA.n30 VDDA.n27 0.227634
R133 VDDA.n59 VDDA.n58 0.189563
R134 VDDA.n19 VDDA.n18 0.185122
R135 VDDA.n38 VDDA.n37 0.185122
R136 VDDA.n41 VDDA.n40 0.185122
R137 VDDA.n22 VDDA.n12 0.168945
R138 VDDA.n23 VDDA.n11 0.168674
R139 VDDA.n23 VDDA.n22 0.153097
R140 VDDA.n4 VDDA.n2 0.152959
R141 VDDA.n54 VDDA.n1 0.152959
R142 VDDA.n44 VDDA.n24 0.147294
R143 VDDA.n19 VDDA.n5 0.141125
R144 VDDA.n24 VDDA.n23 0.105208
R145 VDDA.n34 VDDA.n33 0.105208
R146 VDDA.n35 VDDA.n34 0.105208
R147 VDDA.n29 VDDA.n28 0.105208
R148 VDDA.n30 VDDA.n29 0.086539
R149 VDDA.n19 VDDA.n16 0.0379178
R150 VDDA.n42 VDDA 0.0270625
R151 VDDA.n44 VDDA.n43 0.013
R152 VDDA.n11 VDDA.n10 0.00995724
R153 VDDA.n16 VDDA.n15 0.00995724
R154 VDDA.n18 VDDA.n17 0.00995724
R155 VDDA.n37 VDDA.n36 0.00995724
R156 VDDA.n40 VDDA.n39 0.00995724
R157 VDDA.n56 VDDA.n54 0.009875
R158 cm2_pcell_0.cm2_pcell2_0.S4 cm2_pcell_0.cm2_pcell2_0.S4.t1 158.145
R159 cm2_pcell_0.cm2_pcell2_0.S4.n0 cm2_pcell_0.cm2_pcell2_0.S4.t3 142.477
R160 cm2_pcell_0.cm2_pcell2_0.S4.n0 cm2_pcell_0.cm2_pcell2_0.S4.t2 140.496
R161 cm2_pcell_0.cm2_pcell2_0.S4.n1 cm2_pcell_0.cm2_pcell2_0.S4.t0 140.082
R162 cm2_pcell_0.cm2_pcell2_0.S4.n1 cm2_pcell_0.cm2_pcell2_0.S4.n0 7.35744
R163 cm2_pcell_0.cm2_pcell2_0.S4 cm2_pcell_0.cm2_pcell2_0.S4.n1 0.0463333
R164 cm2_pcell_0.D0.n7 cm2_pcell_0.D0.t8 142.488
R165 cm2_pcell_0.D0.n1 cm2_pcell_0.D0.t12 142.488
R166 cm2_pcell_0.D0.n0 cm2_pcell_0.D0.t7 142.488
R167 cm2_pcell_0.D0.n7 cm2_pcell_0.D0.t9 141.704
R168 cm2_pcell_0.D0.n1 cm2_pcell_0.D0.t13 141.704
R169 cm2_pcell_0.D0.n0 cm2_pcell_0.D0.t6 141.704
R170 cm2_pcell_0.D0.n6 cm2_pcell_0.D0.t10 141.704
R171 cm2_pcell_0.D0.n5 cm2_pcell_0.D0.t11 141.704
R172 cm2_pcell_0.D0.n3 cm2_pcell_0.D0.t3 139.454
R173 cm2_pcell_0.D0.n9 cm2_pcell_0.D0.t1 139.454
R174 cm2_pcell_0.D0.n4 cm2_pcell_0.D0.t5 135.329
R175 cm2_pcell_0.D0.n11 cm2_pcell_0.D0.t2 135.231
R176 cm2_pcell_0.D0.n11 cm2_pcell_0.D0.t4 135.231
R177 cm2_pcell_0.D0.n4 cm2_pcell_0.D0.t0 134.444
R178 cm2_pcell_0.D0.n5 cm2_pcell_0.D0.n4 6.41092
R179 cm2_pcell_0.cm2_pcell2_0.D0 cm2_pcell_0.D0.n11 4.563
R180 cm2_pcell_0.D0.n3 cm2_pcell_0.D0.n2 2.2505
R181 cm2_pcell_0.D0.n9 cm2_pcell_0.D0.n8 2.2505
R182 cm2_pcell_0.D0.n10 cm2_pcell_0.D0.n3 0.829667
R183 cm2_pcell_0.D0.n10 cm2_pcell_0.D0.n9 0.829667
R184 cm2_pcell_0.D0.n2 cm2_pcell_0.D0.n0 0.783833
R185 cm2_pcell_0.D0.n2 cm2_pcell_0.D0.n1 0.783833
R186 cm2_pcell_0.D0.n6 cm2_pcell_0.D0.n5 0.783833
R187 cm2_pcell_0.D0.n8 cm2_pcell_0.D0.n6 0.783833
R188 cm2_pcell_0.D0.n8 cm2_pcell_0.D0.n7 0.783833
R189 cm2_pcell_0.D0.n11 cm2_pcell_0.D0.n10 0.224458
R190 VBPDEC.n3 VBPDEC.t1 221.851
R191 VBPDEC.n1 VBPDEC.t3 221.851
R192 VBPDEC.n6 VBPDEC.t4 140.061
R193 VBPDEC.n7 VBPDEC.t5 139.566
R194 VBPDEC.n0 VBPDEC.t2 108.365
R195 VBPDEC.n4 VBPDEC.t0 108.365
R196 VBPDEC.n5 VBPDEC.n0 15.3463
R197 VBPDEC.n6 VBPDEC.n5 8.1267
R198 VBPDEC.n3 VBPDEC.n2 5.86092
R199 VBPDEC.n2 VBPDEC.n1 4.95104
R200 VBPDEC.n5 VBPDEC.n4 4.79425
R201 VBPDEC VBPDEC.n6 1.21717
R202 VBPDEC.n1 VBPDEC.n0 0.557293
R203 VBPDEC.n4 VBPDEC.n3 0.546515
R204 VBPDEC VBPDEC.n7 0.08175
R205 VBPDEC.n7 VBPDEC 0.063
R206 VBPDEC.n2 VBPDEC 0.0525833
R207 cm2_pcell_0.cm2_pcell2_0.S2 cm2_pcell_0.cm2_pcell2_0.S2.t1 158.273
R208 cm2_pcell_0.cm2_pcell2_0.S2.n0 cm2_pcell_0.cm2_pcell2_0.S2.t2 141.358
R209 cm2_pcell_0.cm2_pcell2_0.S2.n1 cm2_pcell_0.cm2_pcell2_0.S2.t0 140.304
R210 cm2_pcell_0.cm2_pcell2_0.S2.n0 cm2_pcell_0.cm2_pcell2_0.S2.t3 139.566
R211 cm2_pcell_0.cm2_pcell2_0.S2.n1 cm2_pcell_0.cm2_pcell2_0.S2.n0 8.02027
R212 cm2_pcell_0.cm2_pcell2_0.S2 cm2_pcell_0.cm2_pcell2_0.S2.n1 0.063
R213 VBNDEC.n3 VBNDEC.t3 221.851
R214 VBNDEC.n2 VBNDEC.t1 221.851
R215 VBNDEC.n8 VBNDEC.t4 140.244
R216 VBNDEC.n7 VBNDEC.t5 140.056
R217 VBNDEC.n4 VBNDEC.t2 108.365
R218 VBNDEC.n1 VBNDEC.t0 108.365
R219 VBNDEC.n5 VBNDEC.n4 15.0927
R220 VBNDEC.n0 VBNDEC.t6 13.3032
R221 VBNDEC.n3 VBNDEC.n2 11.1702
R222 VBNDEC.n7 VBNDEC.n6 4.63108
R223 VBNDEC.n6 VBNDEC.n0 3.9493
R224 VBNDEC.n6 VBNDEC.n5 3.4105
R225 VBNDEC.n8 VBNDEC.n7 2.67342
R226 VBNDEC.n5 VBNDEC.n1 2.25675
R227 VBNDEC.n2 VBNDEC.n1 0.546515
R228 VBNDEC.n4 VBNDEC.n3 0.527402
R229 VBNDEC VBNDEC.n8 0.063
R230 VBNDEC.n0 VBNDEC 0.0498421
R231 a_4080_n2791.n4 a_4080_n2791.t5 239.399
R232 a_4080_n2791.t0 a_4080_n2791.n4 227.651
R233 a_4080_n2791.n0 a_4080_n2791.t2 222.332
R234 a_4080_n2791.n2 a_4080_n2791.t4 222.332
R235 a_4080_n2791.n1 a_4080_n2791.t7 111.007
R236 a_4080_n2791.n3 a_4080_n2791.t6 111.007
R237 a_4080_n2791.n0 a_4080_n2791.t1 108.365
R238 a_4080_n2791.n2 a_4080_n2791.t3 108.365
R239 a_4080_n2791.n1 a_4080_n2791.n0 2.64217
R240 a_4080_n2791.n3 a_4080_n2791.n2 2.64217
R241 a_4080_n2791.n3 a_4080_n2791.n1 0.817167
R242 a_4080_n2791.n4 a_4080_n2791.n3 0.302583
R243 GNDA.n4 GNDA.n3 1179.3
R244 GNDA.t11 GNDA.t0 547.01
R245 GNDA.t3 GNDA.t6 256.649
R246 GNDA.t1 GNDA.t2 232.725
R247 GNDA.n3 GNDA.t9 231.637
R248 GNDA.n10 GNDA.t12 222.284
R249 GNDA.n2 GNDA.t4 222.023
R250 GNDA.n2 GNDA.t5 221.905
R251 GNDA.n12 GNDA.t8 221.851
R252 GNDA.n12 GNDA.t7 221.851
R253 GNDA.n8 GNDA.t15 221.738
R254 GNDA.n3 GNDA.t14 179.436
R255 GNDA.n7 GNDA.t10 127.977
R256 GNDA.t0 GNDA.t1 102.225
R257 GNDA.t6 GNDA.t11 102.225
R258 GNDA.t2 GNDA.t13 52.2002
R259 GNDA.t14 GNDA.t3 47.8502
R260 GNDA.n9 GNDA.n7 4.538
R261 GNDA.n15 GNDA.n14 4.39425
R262 GNDA.n9 GNDA.n8 3.34894
R263 GNDA.n15 GNDA.n0 1.64425
R264 GNDA.n10 GNDA.n9 1.50919
R265 GNDA.n11 GNDA.n10 1.49623
R266 GNDA.n4 GNDA.n0 0.956486
R267 GNDA.n13 GNDA.n0 0.59425
R268 GNDA.n6 GNDA.n1 0.59425
R269 GNDA.n14 GNDA.n13 0.59425
R270 GNDA.n11 GNDA.n1 0.461438
R271 GNDA.n14 GNDA.n11 0.311437
R272 GNDA.n8 GNDA.n1 0.227062
R273 GNDA.n7 GNDA.n6 0.164562
R274 GNDA.n13 GNDA.n12 0.159799
R275 GNDA.n5 GNDA.n2 0.091223
R276 GNDA.n5 GNDA.n4 0.0648892
R277 GNDA GNDA.n15 0.0270625
R278 GNDA.n6 GNDA.n5 0.0141985
R279 a_4602_n3479.t1 a_4602_n3479.n1 229.328
R280 a_4602_n3479.n1 a_4602_n3479.t0 226.986
R281 a_4602_n3479.n0 a_4602_n3479.t3 127.692
R282 a_4602_n3479.n1 a_4602_n3479.n0 12.484
R283 a_4602_n3479.n0 a_4602_n3479.t2 10.584
R284 ROUT.n1 ROUT.t3 134.847
R285 ROUT.n2 ROUT.t1 134.246
R286 ROUT.n1 ROUT.n0 8.36161
R287 ROUT.t4 ROUT.t5 5.8809
R288 ROUT.t2 ROUT.t4 5.0615
R289 ROUT.n0 ROUT.t0 2.9407
R290 ROUT.n0 ROUT.t2 2.9407
R291 ROUT.n2 ROUT.n1 0.601043
R292 ROUT ROUT.n2 0.402674
R293 a_11186_n55.n0 a_11186_n55.t2 135.572
R294 a_11186_n55.n1 a_11186_n55.t0 135.572
R295 a_11186_n55.n0 a_11186_n55.t3 134.246
R296 a_11186_n55.t1 a_11186_n55.n1 134.246
R297 a_11186_n55.n1 a_11186_n55.n0 1.1418
R298 cm2_pcell_0.D1.n4 cm2_pcell_0.D1.t1 221.851
R299 cm2_pcell_0.D1.n2 cm2_pcell_0.D1.t3 221.851
R300 cm2_pcell_0.D1.n0 cm2_pcell_0.D1.t5 140.625
R301 cm2_pcell_0.D1.n0 cm2_pcell_0.D1.t4 140.244
R302 cm2_pcell_0.D1.n3 cm2_pcell_0.D1.t6 113.648
R303 cm2_pcell_0.D1.n1 cm2_pcell_0.D1.t7 113.648
R304 cm2_pcell_0.D1.n3 cm2_pcell_0.D1.t0 108.365
R305 cm2_pcell_0.D1.n1 cm2_pcell_0.D1.t2 108.365
R306 cm2_pcell_0.cm2_pcell2_0.D1 cm2_pcell_0.D1.n5 12.9957
R307 cm2_pcell_0.D1.n5 cm2_pcell_0.D1.n4 1.60385
R308 cm2_pcell_0.D1.n4 cm2_pcell_0.D1.n3 0.557293
R309 cm2_pcell_0.D1.n2 cm2_pcell_0.D1.n1 0.557293
R310 cm2_pcell_0.D1.n5 cm2_pcell_0.D1.n2 0.266714
R311 cm2_pcell_0.cm2_pcell2_0.D1 cm2_pcell_0.D1.n0 0.063
R312 a_4080_n3027.n1 a_4080_n3027.t1 239.831
R313 a_4080_n3027.t0 a_4080_n3027.n1 226.853
R314 a_4080_n3027.n0 a_4080_n3027.t2 223.633
R315 a_4080_n3027.n0 a_4080_n3027.t3 221.851
R316 a_4080_n3027.n1 a_4080_n3027.n0 5.73071
R317 VBPLV.n4 VBPLV.t0 232.263
R318 VBPLV.n4 VBPLV.t1 222.117
R319 VBPLV.n0 VBPLV.t2 139.454
R320 VBPLV.n1 VBPLV.t4 139.454
R321 VBPLV.n0 VBPLV.t3 135.197
R322 VBPLV.n2 VBPLV.t5 134.625
R323 VBPLV.n3 VBPLV.t6 17.157
R324 VBPLV VBPLV.n4 11.263
R325 VBPLV.n3 VBPLV.n2 4.5005
R326 VBPLV VBPLV.n3 1.10467
R327 VBPLV.n1 VBPLV.n0 0.701587
R328 VBPLV.n2 VBPLV.n1 0.51454
R329 VBNLV.n1 VBNLV.t3 222.043
R330 VBNLV.n1 VBNLV.t1 222.043
R331 VBNLV.n5 VBNLV.t4 140.061
R332 VBNLV.n6 VBNLV.t5 139.566
R333 VBNLV.n2 VBNLV.t2 108.754
R334 VBNLV.n3 VBNLV.t0 108.365
R335 VBNLV.n0 VBNLV.t6 20.8855
R336 VBNLV.n4 VBNLV.n3 7.91883
R337 VBNLV.n5 VBNLV.n4 5.02291
R338 VBNLV.n4 VBNLV.n0 3.68368
R339 VBNLV.n6 VBNLV.n5 3.40258
R340 VBNLV.n3 VBNLV.n2 0.310917
R341 VBNLV.n2 VBNLV.n1 0.224458
R342 VBNLV VBNLV.n6 0.063
R343 VBNLV.n0 VBNLV 0.0498421
R344 a_6498_n2100.t0 a_6498_n2100.n0 239.25
R345 a_6498_n2100.n0 a_6498_n2100.t2 222.119
R346 a_6498_n2100.n0 a_6498_n2100.t1 222.119
R347 a_5864_n2100.t0 a_5864_n2100.n0 233.361
R348 a_5864_n2100.n0 a_5864_n2100.t1 229.339
R349 a_5864_n2100.n0 a_5864_n2100.t2 227.399
R350 cm2_pcell_0.cm2_pcell2_0.S3.n1 cm2_pcell_0.cm2_pcell2_0.S3.t0 157.346
R351 cm2_pcell_0.cm2_pcell2_0.S3.n0 cm2_pcell_0.cm2_pcell2_0.S3.t3 142.179
R352 cm2_pcell_0.cm2_pcell2_0.S3.n0 cm2_pcell_0.cm2_pcell2_0.S3.t2 140.314
R353 cm2_pcell_0.cm2_pcell2_0.S3.n2 cm2_pcell_0.cm2_pcell2_0.S3.t1 140.065
R354 cm2_pcell_0.cm2_pcell2_0.S3.n1 cm2_pcell_0.cm2_pcell2_0.S3.n0 7.42011
R355 cm2_pcell_0.cm2_pcell2_0.S3 cm2_pcell_0.cm2_pcell2_0.S3.n2 0.063
R356 cm2_pcell_0.cm2_pcell2_0.S3.n2 cm2_pcell_0.cm2_pcell2_0.S3.n1 0.0171667
R357 cm2_pcell_0.cm2_pcell2_0.S1.n1 cm2_pcell_0.cm2_pcell2_0.S1.t0 157.49
R358 cm2_pcell_0.cm2_pcell2_0.S1.n0 cm2_pcell_0.cm2_pcell2_0.S1.t3 142.079
R359 cm2_pcell_0.cm2_pcell2_0.S1.n1 cm2_pcell_0.cm2_pcell2_0.S1.t1 140.304
R360 cm2_pcell_0.cm2_pcell2_0.S1.n0 cm2_pcell_0.cm2_pcell2_0.S1.t2 139.327
R361 cm2_pcell_0.cm2_pcell2_0.S1.n1 cm2_pcell_0.cm2_pcell2_0.S1.n0 7.54544
R362 cm2_pcell_0.cm2_pcell2_0.S1 cm2_pcell_0.cm2_pcell2_0.S1.n1 0.063
R363 a_7128_n494.n0 a_7128_n494.t2 356.854
R364 a_7128_n494.n0 a_7128_n494.t0 15.3866
R365 a_7128_n494.t1 a_7128_n494.n0 15.3866
C0 VBPDEC cm2_pcell_0.cm2_pcell2_0.S4 0.0483f
C1 a_7075_n3098# VBNDEC 0.02736f
C2 VDDA cm2_pcell_0.cm2_pcell2_0.S3 2.05072f
C3 VDDA a_7053_n520# 0.3015f
C4 cm2_pcell_0.cm2_pcell2_0.S1 VBPLV 0.01639f
C5 VBPLV ROUT 0.25958f
C6 cm2_pcell_0.cm2_pcell2_0.S0 cm2_pcell_0.cm2_pcell2_0.S2 1.24591f
C7 cm2_pcell_0.cm2_pcell2_0.S1 cm2_pcell_0.cm2_pcell2_0.S2 0.7893f
C8 cm2_pcell_0.cm2_pcell2_0.S4 VBNLV 0.06438f
C9 cm2_pcell_0.cm2_pcell2_0.S4 VBNDEC 0.29277f
C10 VBPDEC VBPLV 0.32439f
C11 VDDA a_7717_n1120# 0.39996f
C12 VBPDEC a_6960_n2188# 0.02655f
C13 VBPDEC cm2_pcell_0.cm2_pcell2_0.S2 0.21449f
C14 a_6960_n2188# a_6960_n1912# 0.02286f
C15 cm2_pcell_0.cm2_pcell2_0.S4 cm2_pcell_0.cm2_pcell2_0.S3 1.13576f
C16 a_7053_n81# VDDA 1.41184f
C17 VBNDEC a_4929_n3098# 0.02764f
C18 VDDA cm2_pcell_0.cm2_pcell2_0.S4 3.17848f
C19 cm2_pcell_0.cm2_pcell2_0.S1 cm2_pcell_0.cm2_pcell2_0.S0 0.80785f
C20 VBPLV VBNLV 0.11339f
C21 cm2_pcell_0.cm2_pcell2_0.S1 ROUT 0.01357f
C22 a_11259_n81# ROUT 0.08397f
C23 a_5776_n2188# a_5776_n1912# 0.02286f
C24 VBPLV VBNDEC 0.08863f
C25 VBNLV cm2_pcell_0.cm2_pcell2_0.S2 0.03773f
C26 VBPLV a_7053_n1120# 0.06598f
C27 VBNDEC cm2_pcell_0.cm2_pcell2_0.S2 0.07818f
C28 VBPDEC cm2_pcell_0.cm2_pcell2_0.S0 0.35106f
C29 cm2_pcell_0.cm2_pcell2_0.S1 VBPDEC 0.05993f
C30 VBPLV a_9099_n520# 0.02974f
C31 a_5776_n2188# VBNDEC 0.02882f
C32 VBPLV cm2_pcell_0.cm2_pcell2_0.S3 0.09782f
C33 VBPLV a_7053_n520# 0.03219f
C34 VDDA VBPLV 6.09482f
C35 cm2_pcell_0.cm2_pcell2_0.S2 cm2_pcell_0.cm2_pcell2_0.S3 1.05222f
C36 VDDA cm2_pcell_0.cm2_pcell2_0.S2 2.42731f
C37 VBPDEC a_5776_n1912# 0.02697f
C38 VBNLV cm2_pcell_0.cm2_pcell2_0.S0 0.08581f
C39 cm2_pcell_0.cm2_pcell2_0.S1 VBNLV 0.0921f
C40 a_4996_n1864# VBPLV 0.02063f
C41 a_4005_n2817# a_4005_n3115# 0.015f
C42 cm2_pcell_0.cm2_pcell2_0.S0 VBNDEC 0.04477f
C43 cm2_pcell_0.cm2_pcell2_0.S1 VBNDEC 0.10137f
C44 VBPLV a_7717_n1120# 0.0755f
C45 a_5809_n2723# VBNLV 0.02804f
C46 a_5809_n2723# VBNDEC 0.01035f
C47 VBPDEC VBNLV 0.80363f
C48 a_4929_n3098# a_4787_n3115# 0.04234f
C49 VBPDEC VBNDEC 2.5778f
C50 cm2_pcell_0.cm2_pcell2_0.S0 cm2_pcell_0.cm2_pcell2_0.S3 0.65201f
C51 cm2_pcell_0.cm2_pcell2_0.S1 cm2_pcell_0.cm2_pcell2_0.S3 3.83598f
C52 cm2_pcell_0.cm2_pcell2_0.S3 ROUT 0.04838f
C53 VDDA cm2_pcell_0.cm2_pcell2_0.S0 6.06684f
C54 cm2_pcell_0.cm2_pcell2_0.S1 VDDA 2.24135f
C55 VDDA a_11259_n81# 1.21922f
C56 a_6960_n1912# VBNDEC 0.02781f
C57 a_5776_n1912# VBNDEC 0.01092f
C58 VDDA ROUT 8.46658f
C59 VBPLV cm2_pcell_0.cm2_pcell2_0.S4 0.24016f
C60 VBPLV a_4214_n2282# 0.01119f
C61 VBPDEC cm2_pcell_0.cm2_pcell2_0.S3 0.04279f
C62 cm2_pcell_0.cm2_pcell2_0.S4 cm2_pcell_0.cm2_pcell2_0.S2 3.55677f
C63 VBPDEC VDDA 0.17653f
C64 a_7075_n2723# VBNLV 0.02789f
C65 VBNLV VBNDEC 2.31944f
C66 VBNLV cm2_pcell_0.cm2_pcell2_0.S3 0.26736f
C67 VBNDEC cm2_pcell_0.cm2_pcell2_0.S3 0.12549f
C68 VDDA VBNLV 0.74221f
C69 cm2_pcell_0.cm2_pcell2_0.S4 cm2_pcell_0.cm2_pcell2_0.S0 0.80349f
C70 a_7053_n81# ROUT 0.14001f
C71 cm2_pcell_0.cm2_pcell2_0.S1 cm2_pcell_0.cm2_pcell2_0.S4 0.17741f
C72 VDDA VBNDEC 0.55365f
C73 a_4787_n3115# a_4787_n2817# 0.015f
C74 VDDA a_7053_n1120# 0.4519f
C75 VDDA a_9099_n520# 0.28979f
C76 VBPLV GNDA 3.73927f
C77 ROUT GNDA 11.76964f
C78 VBNLV GNDA 4.11963f
C79 VBPDEC GNDA 2.2221f
C80 VBNDEC GNDA 7.13538f
C81 VDDA GNDA 70.87076f
C82 a_7075_n3479# GNDA 0.24801f $ **FLOATING
C83 a_4469_n3479# GNDA 0.27572f $ **FLOATING
C84 a_7075_n3098# GNDA 0.23625f $ **FLOATING
C85 a_4929_n3098# GNDA 0.2216f $ **FLOATING
C86 a_4787_n3115# GNDA 0.18327f $ **FLOATING
C87 a_4005_n3115# GNDA 0.22622f $ **FLOATING
C88 a_7075_n2723# GNDA 0.23867f $ **FLOATING
C89 a_5809_n2723# GNDA 0.24765f $ **FLOATING
C90 a_4787_n2817# GNDA 0.21832f $ **FLOATING
C91 a_4005_n2817# GNDA 0.22368f $ **FLOATING
C92 a_6960_n2188# GNDA 0.18027f $ **FLOATING
C93 a_5776_n2188# GNDA 0.17916f $ **FLOATING
C94 a_6960_n1912# GNDA 0.18226f $ **FLOATING
C95 a_5776_n1912# GNDA 0.18241f $ **FLOATING
C96 a_4996_n2282# GNDA 0.18717f $ **FLOATING
C97 a_4214_n2282# GNDA 0.18294f $ **FLOATING
C98 a_4996_n1864# GNDA 0.18848f $ **FLOATING
C99 a_4214_n1864# GNDA 0.18388f $ **FLOATING
C100 a_7717_n1120# GNDA 0.05347f $ **FLOATING
C101 a_7053_n1120# GNDA 0.01074f $ **FLOATING
C102 a_9099_n520# GNDA 0.03847f $ **FLOATING
C103 a_11259_n81# GNDA 0.18138f $ **FLOATING
C104 a_7053_n81# GNDA 0.03843f $ **FLOATING
C105 cm2_pcell_0.cm2_pcell2_0.S3 GNDA 0.26788f
C106 cm2_pcell_0.cm2_pcell2_0.S1 GNDA 0.2916f
C107 cm2_pcell_0.cm2_pcell2_0.S2 GNDA 2.99356f
C108 cm2_pcell_0.cm2_pcell2_0.S4 GNDA 3.27416f
C109 cm2_pcell_0.cm2_pcell2_0.S0 GNDA 2.30752f
C110 cm2_pcell_0.cm2_pcell2_0.S1.t0 GNDA 0.39374f
C111 cm2_pcell_0.cm2_pcell2_0.S1.t2 GNDA 0.19462f
C112 cm2_pcell_0.cm2_pcell2_0.S1.t3 GNDA 0.21619f
C113 cm2_pcell_0.cm2_pcell2_0.S1.n0 GNDA 1.60492f
C114 cm2_pcell_0.cm2_pcell2_0.S1.t1 GNDA 0.20263f
C115 cm2_pcell_0.cm2_pcell2_0.S1.n1 GNDA 3.37677f
C116 cm2_pcell_0.cm2_pcell2_0.S3.t0 GNDA 0.38205f
C117 cm2_pcell_0.cm2_pcell2_0.S3.t2 GNDA 0.19864f
C118 cm2_pcell_0.cm2_pcell2_0.S3.t3 GNDA 0.2028f
C119 cm2_pcell_0.cm2_pcell2_0.S3.n0 GNDA 1.78846f
C120 cm2_pcell_0.cm2_pcell2_0.S3.n1 GNDA 2.76369f
C121 cm2_pcell_0.cm2_pcell2_0.S3.t1 GNDA 0.19467f
C122 cm2_pcell_0.cm2_pcell2_0.S3.n2 GNDA 0.35783f
C123 VBNLV.t6 GNDA 0.53779f
C124 VBNLV.n0 GNDA 0.1895f
C125 VBNLV.t2 GNDA 0.09539f
C126 VBNLV.t1 GNDA 0.01931f
C127 VBNLV.t3 GNDA 0.01931f
C128 VBNLV.n1 GNDA 0.07175f
C129 VBNLV.n2 GNDA 0.09138f
C130 VBNLV.t0 GNDA 0.09524f
C131 VBNLV.n3 GNDA 0.05563f
C132 VBNLV.n4 GNDA 0.40112f
C133 VBNLV.t4 GNDA 0.06249f
C134 VBNLV.n5 GNDA 0.3608f
C135 VBNLV.t5 GNDA 0.06035f
C136 VBNLV.n6 GNDA 0.23279f
C137 VBPLV.t6 GNDA 2.32652f
C138 VBPLV.t3 GNDA 0.0924f
C139 VBPLV.t2 GNDA 0.34803f
C140 VBPLV.n0 GNDA 0.30808f
C141 VBPLV.t4 GNDA 0.34803f
C142 VBPLV.n1 GNDA 0.14391f
C143 VBPLV.t5 GNDA 0.09171f
C144 VBPLV.n2 GNDA 0.17226f
C145 VBPLV.n3 GNDA 0.78347f
C146 VBPLV.t1 GNDA 0.03087f
C147 VBPLV.t0 GNDA 0.03937f
C148 VBPLV.n4 GNDA 0.67262f
C149 a_4080_n3027.t2 GNDA 0.05539f
C150 a_4080_n3027.t3 GNDA 0.05331f
C151 a_4080_n3027.n0 GNDA 0.5884f
C152 a_4080_n3027.t1 GNDA 0.09815f
C153 a_4080_n3027.n1 GNDA 1.64869f
C154 a_4080_n3027.t0 GNDA 0.05605f
C155 ROUT.t3 GNDA 0.02283f
C156 ROUT.t0 GNDA 1.30025f
C157 ROUT.t5 GNDA 1.87382f
C158 ROUT.t4 GNDA 2.13764f
C159 ROUT.t2 GNDA 1.56407f
C160 ROUT.n0 GNDA 1.3493f
C161 ROUT.n1 GNDA 0.19702f
C162 ROUT.t1 GNDA 0.02268f
C163 ROUT.n2 GNDA 0.02664f
C164 a_4080_n2791.t2 GNDA 0.03016f
C165 a_4080_n2791.t1 GNDA 0.14825f
C166 a_4080_n2791.n0 GNDA 0.16973f
C167 a_4080_n2791.t7 GNDA 0.15058f
C168 a_4080_n2791.n1 GNDA 0.279f
C169 a_4080_n2791.t6 GNDA 0.15058f
C170 a_4080_n2791.t3 GNDA 0.14825f
C171 a_4080_n2791.t4 GNDA 0.03016f
C172 a_4080_n2791.n2 GNDA 0.16973f
C173 a_4080_n2791.n3 GNDA 0.29912f
C174 a_4080_n2791.t5 GNDA 0.05237f
C175 a_4080_n2791.n4 GNDA 0.83928f
C176 a_4080_n2791.t0 GNDA 0.03278f
C177 VBNDEC.t5 GNDA 0.08977f
C178 VBNDEC.t6 GNDA 1.43368f
C179 VBNDEC.n0 GNDA 0.2112f
C180 VBNDEC.t0 GNDA 0.14211f
C181 VBNDEC.n1 GNDA 0.09571f
C182 VBNDEC.t2 GNDA 0.14211f
C183 VBNDEC.t1 GNDA 0.02878f
C184 VBNDEC.n2 GNDA 0.16872f
C185 VBNDEC.t3 GNDA 0.02878f
C186 VBNDEC.n3 GNDA 0.23193f
C187 VBNDEC.n4 GNDA 0.44337f
C188 VBNDEC.n5 GNDA 0.27955f
C189 VBNDEC.n6 GNDA 0.65817f
C190 VBNDEC.n7 GNDA 0.44043f
C191 VBNDEC.t4 GNDA 0.09426f
C192 VBNDEC.n8 GNDA 0.40081f
C193 cm2_pcell_0.cm2_pcell2_0.S2.t2 GNDA 0.20734f
C194 cm2_pcell_0.cm2_pcell2_0.S2.t3 GNDA 0.19458f
C195 cm2_pcell_0.cm2_pcell2_0.S2.n0 GNDA 1.54108f
C196 cm2_pcell_0.cm2_pcell2_0.S2.t0 GNDA 0.20013f
C197 cm2_pcell_0.cm2_pcell2_0.S2.n1 GNDA 0.76408f
C198 cm2_pcell_0.cm2_pcell2_0.S2.t1 GNDA 0.39974f
C199 VBPDEC.t2 GNDA 0.1401f
C200 VBPDEC.n0 GNDA 0.2903f
C201 VBPDEC.t3 GNDA 0.02838f
C202 VBPDEC.n1 GNDA 0.09142f
C203 VBPDEC.n2 GNDA 0.17301f
C204 VBPDEC.t1 GNDA 0.02838f
C205 VBPDEC.n3 GNDA 0.08096f
C206 VBPDEC.t0 GNDA 0.1401f
C207 VBPDEC.n4 GNDA 0.10554f
C208 VBPDEC.n5 GNDA 0.62142f
C209 VBPDEC.t4 GNDA 0.09192f
C210 VBPDEC.n6 GNDA 0.49433f
C211 VBPDEC.t5 GNDA 0.08878f
C212 VBPDEC.n7 GNDA 0.13349f
C213 cm2_pcell_0.D0.t4 GNDA 0.04207f
C214 cm2_pcell_0.D0.t2 GNDA 0.04207f
C215 cm2_pcell_0.D0.t3 GNDA 0.15904f
C216 cm2_pcell_0.D0.t7 GNDA 0.16048f
C217 cm2_pcell_0.D0.t6 GNDA 0.15996f
C218 cm2_pcell_0.D0.n0 GNDA 0.19996f
C219 cm2_pcell_0.D0.t12 GNDA 0.16046f
C220 cm2_pcell_0.D0.t13 GNDA 0.15996f
C221 cm2_pcell_0.D0.n1 GNDA 0.19556f
C222 cm2_pcell_0.D0.n2 GNDA 0.04891f
C223 cm2_pcell_0.D0.n3 GNDA 0.08386f
C224 cm2_pcell_0.D0.t1 GNDA 0.15904f
C225 cm2_pcell_0.D0.t5 GNDA 0.0423f
C226 cm2_pcell_0.D0.t0 GNDA 0.04183f
C227 cm2_pcell_0.D0.n4 GNDA 0.16659f
C228 cm2_pcell_0.D0.t11 GNDA 0.15996f
C229 cm2_pcell_0.D0.n5 GNDA 0.18631f
C230 cm2_pcell_0.D0.t10 GNDA 0.15996f
C231 cm2_pcell_0.D0.n6 GNDA 0.10596f
C232 cm2_pcell_0.D0.t8 GNDA 0.16046f
C233 cm2_pcell_0.D0.t9 GNDA 0.15996f
C234 cm2_pcell_0.D0.n7 GNDA 0.19556f
C235 cm2_pcell_0.D0.n8 GNDA 0.04891f
C236 cm2_pcell_0.D0.n9 GNDA 0.08386f
C237 cm2_pcell_0.D0.n10 GNDA 0.06653f
C238 cm2_pcell_0.D0.n11 GNDA 0.14113f
C239 cm2_pcell_0.cm2_pcell2_0.S4.t0 GNDA 0.21475f
C240 cm2_pcell_0.cm2_pcell2_0.S4.t3 GNDA 0.22412f
C241 cm2_pcell_0.cm2_pcell2_0.S4.t2 GNDA 0.22155f
C242 cm2_pcell_0.cm2_pcell2_0.S4.n0 GNDA 2.08687f
C243 cm2_pcell_0.cm2_pcell2_0.S4.n1 GNDA 0.6997f
C244 cm2_pcell_0.cm2_pcell2_0.S4.t1 GNDA 0.44343f
C245 VDDA.n0 GNDA 0.15386f
C246 VDDA.n1 GNDA 0.15982f
C247 VDDA.n2 GNDA 0.12808f
C248 VDDA.n3 GNDA 0.32686f
C249 VDDA.n4 GNDA 0.30044f
C250 VDDA.n5 GNDA 0.06685f
C251 VDDA.n6 GNDA 0.23204f
C252 VDDA.n7 GNDA 0.59648f
C253 VDDA.n9 GNDA 0.41636f
C254 VDDA.t3 GNDA 4.43225f
C255 VDDA.t19 GNDA 0.02323f
C256 VDDA.t16 GNDA 0.02323f
C257 VDDA.t15 GNDA 0.02323f
C258 VDDA.n10 GNDA 0.0771f
C259 VDDA.t13 GNDA 0.08773f
C260 VDDA.n11 GNDA 0.10203f
C261 VDDA.t42 GNDA 0.02309f
C262 VDDA.t18 GNDA 0.02309f
C263 VDDA.n12 GNDA 0.08243f
C264 VDDA.t44 GNDA 0.02309f
C265 VDDA.t38 GNDA 0.02309f
C266 VDDA.n13 GNDA 0.09361f
C267 VDDA.t45 GNDA 0.02309f
C268 VDDA.t39 GNDA 0.02309f
C269 VDDA.n14 GNDA 0.09318f
C270 VDDA.t21 GNDA 0.02323f
C271 VDDA.t22 GNDA 0.02323f
C272 VDDA.n15 GNDA 0.0771f
C273 VDDA.t20 GNDA 0.08773f
C274 VDDA.n16 GNDA 0.04422f
C275 VDDA.t12 GNDA 0.02323f
C276 VDDA.t11 GNDA 0.02323f
C277 VDDA.n17 GNDA 0.0771f
C278 VDDA.t9 GNDA 0.08773f
C279 VDDA.n18 GNDA 0.1093f
C280 VDDA.n19 GNDA 0.11826f
C281 VDDA.n20 GNDA 0.08462f
C282 VDDA.n21 GNDA 0.09937f
C283 VDDA.n22 GNDA 0.07981f
C284 VDDA.t17 GNDA 0.08773f
C285 VDDA.n23 GNDA 0.12704f
C286 VDDA.n24 GNDA 0.05573f
C287 VDDA.t34 GNDA 0.02323f
C288 VDDA.t33 GNDA 0.02323f
C289 VDDA.t41 GNDA 0.02309f
C290 VDDA.t40 GNDA 0.02309f
C291 VDDA.n25 GNDA 0.09361f
C292 VDDA.t36 GNDA 0.02309f
C293 VDDA.t43 GNDA 0.02309f
C294 VDDA.n26 GNDA 0.09361f
C295 VDDA.t31 GNDA 0.02309f
C296 VDDA.t37 GNDA 0.02309f
C297 VDDA.n27 GNDA 0.08998f
C298 VDDA.t30 GNDA 0.02323f
C299 VDDA.n28 GNDA 0.10972f
C300 VDDA.t29 GNDA 0.08773f
C301 VDDA.n29 GNDA 0.04514f
C302 VDDA.n30 GNDA 0.08104f
C303 VDDA.n31 GNDA 0.09814f
C304 VDDA.n32 GNDA 0.08524f
C305 VDDA.n33 GNDA 0.06774f
C306 VDDA.t32 GNDA 0.08773f
C307 VDDA.n34 GNDA 0.04725f
C308 VDDA.n35 GNDA 0.10972f
C309 VDDA.t24 GNDA 0.02323f
C310 VDDA.t25 GNDA 0.02323f
C311 VDDA.n36 GNDA 0.0771f
C312 VDDA.t23 GNDA 0.08773f
C313 VDDA.n37 GNDA 0.1093f
C314 VDDA.n38 GNDA 0.2536f
C315 VDDA.t27 GNDA 0.02323f
C316 VDDA.t28 GNDA 0.02323f
C317 VDDA.n39 GNDA 0.0771f
C318 VDDA.t26 GNDA 0.08773f
C319 VDDA.n40 GNDA 0.1093f
C320 VDDA.n41 GNDA 0.28878f
C321 VDDA.n42 GNDA 0.10452f
C322 VDDA.n43 GNDA 0.06293f
C323 VDDA.n45 GNDA 0.05571f
C324 VDDA.n46 GNDA 0.7077f
C325 VDDA.t14 GNDA 1.41176f
C326 VDDA.t2 GNDA 1.41876f
C327 VDDA.t8 GNDA 1.41876f
C328 VDDA.t7 GNDA 1.41526f
C329 VDDA.t35 GNDA 1.41876f
C330 VDDA.t4 GNDA 1.41876f
C331 VDDA.t10 GNDA 1.4565f
C332 VDDA.n47 GNDA 1.26406f
C333 VDDA.t0 GNDA 1.0037f
C334 VDDA.t1 GNDA 1.18482f
C335 VDDA.n48 GNDA 1.46359f
C336 VDDA.t5 GNDA 3.07335f
C337 VDDA.n49 GNDA 0.0254f
C338 VDDA.n50 GNDA 0.87935f
C339 VDDA.n51 GNDA 0.94956f
C340 VDDA.n52 GNDA 0.12865f
C341 VDDA.n53 GNDA 0.30362f
C342 VDDA.n54 GNDA 0.15053f
C343 VDDA.t6 GNDA 0.01281f
C344 VDDA.n55 GNDA 0.14901f
C345 VDDA.n56 GNDA 0.13017f
C346 VDDA.n57 GNDA 0.18598f
C347 VDDA.n58 GNDA 0.05147f
C348 VDDA.n59 GNDA 0.15755f
C349 VDDA.n60 GNDA 0.06723f
C350 VDDA.n61 GNDA 0.18857f
C351 VDDA.n62 GNDA 0.23399f
C352 VDDA.n63 GNDA 0.12432f
C353 cm2_pcell_0.cm2_pcell2_0.S0.t0 GNDA 0.07426f
C354 cm2_pcell_0.cm2_pcell2_0.S0.t4 GNDA 0.07421f
C355 cm2_pcell_0.cm2_pcell2_0.S0.n0 GNDA 0.13951f
C356 cm2_pcell_0.cm2_pcell2_0.S0.t2 GNDA 0.07421f
C357 cm2_pcell_0.cm2_pcell2_0.S0.t1 GNDA 0.28052f
C358 cm2_pcell_0.cm2_pcell2_0.S0.t12 GNDA 0.28306f
C359 cm2_pcell_0.cm2_pcell2_0.S0.t13 GNDA 0.28214f
C360 cm2_pcell_0.cm2_pcell2_0.S0.n1 GNDA 0.35268f
C361 cm2_pcell_0.cm2_pcell2_0.S0.t9 GNDA 0.28302f
C362 cm2_pcell_0.cm2_pcell2_0.S0.t8 GNDA 0.28214f
C363 cm2_pcell_0.cm2_pcell2_0.S0.n2 GNDA 0.34492f
C364 cm2_pcell_0.cm2_pcell2_0.S0.n3 GNDA 0.08627f
C365 cm2_pcell_0.cm2_pcell2_0.S0.n4 GNDA 0.1486f
C366 cm2_pcell_0.cm2_pcell2_0.S0.t3 GNDA 0.28052f
C367 cm2_pcell_0.cm2_pcell2_0.S0.t6 GNDA 0.28302f
C368 cm2_pcell_0.cm2_pcell2_0.S0.t10 GNDA 0.28214f
C369 cm2_pcell_0.cm2_pcell2_0.S0.n5 GNDA 0.34492f
C370 cm2_pcell_0.cm2_pcell2_0.S0.t7 GNDA 0.28306f
C371 cm2_pcell_0.cm2_pcell2_0.S0.t11 GNDA 0.28214f
C372 cm2_pcell_0.cm2_pcell2_0.S0.n6 GNDA 0.35268f
C373 cm2_pcell_0.cm2_pcell2_0.S0.n7 GNDA 0.08627f
C374 cm2_pcell_0.cm2_pcell2_0.S0.n8 GNDA 0.1486f
C375 cm2_pcell_0.cm2_pcell2_0.S0.n9 GNDA 0.1223f
C376 cm2_pcell_0.cm2_pcell2_0.S0.n10 GNDA 0.13547f
C377 cm2_pcell_0.cm2_pcell2_0.S0.n11 GNDA 0.34481f
C378 cm2_pcell_0.cm2_pcell2_0.S0.n12 GNDA 0.25812f
C379 cm2_pcell_0.cm2_pcell2_0.S0.t5 GNDA 0.07421f
.ends

