magic
tech sky130A
magscale 1 2
timestamp 1750133197
<< metal3 >>
rect -1904 1652 -1132 1680
rect -1904 1228 -1216 1652
rect -1152 1228 -1132 1652
rect -1904 1200 -1132 1228
rect -892 1652 -120 1680
rect -892 1228 -204 1652
rect -140 1228 -120 1652
rect -892 1200 -120 1228
rect 120 1652 892 1680
rect 120 1228 808 1652
rect 872 1228 892 1652
rect 120 1200 892 1228
rect 1132 1652 1904 1680
rect 1132 1228 1820 1652
rect 1884 1228 1904 1652
rect 1132 1200 1904 1228
rect -1904 932 -1132 960
rect -1904 508 -1216 932
rect -1152 508 -1132 932
rect -1904 480 -1132 508
rect -892 932 -120 960
rect -892 508 -204 932
rect -140 508 -120 932
rect -892 480 -120 508
rect 120 932 892 960
rect 120 508 808 932
rect 872 508 892 932
rect 120 480 892 508
rect 1132 932 1904 960
rect 1132 508 1820 932
rect 1884 508 1904 932
rect 1132 480 1904 508
rect -1904 212 -1132 240
rect -1904 -212 -1216 212
rect -1152 -212 -1132 212
rect -1904 -240 -1132 -212
rect -892 212 -120 240
rect -892 -212 -204 212
rect -140 -212 -120 212
rect -892 -240 -120 -212
rect 120 212 892 240
rect 120 -212 808 212
rect 872 -212 892 212
rect 120 -240 892 -212
rect 1132 212 1904 240
rect 1132 -212 1820 212
rect 1884 -212 1904 212
rect 1132 -240 1904 -212
rect -1904 -508 -1132 -480
rect -1904 -932 -1216 -508
rect -1152 -932 -1132 -508
rect -1904 -960 -1132 -932
rect -892 -508 -120 -480
rect -892 -932 -204 -508
rect -140 -932 -120 -508
rect -892 -960 -120 -932
rect 120 -508 892 -480
rect 120 -932 808 -508
rect 872 -932 892 -508
rect 120 -960 892 -932
rect 1132 -508 1904 -480
rect 1132 -932 1820 -508
rect 1884 -932 1904 -508
rect 1132 -960 1904 -932
rect -1904 -1228 -1132 -1200
rect -1904 -1652 -1216 -1228
rect -1152 -1652 -1132 -1228
rect -1904 -1680 -1132 -1652
rect -892 -1228 -120 -1200
rect -892 -1652 -204 -1228
rect -140 -1652 -120 -1228
rect -892 -1680 -120 -1652
rect 120 -1228 892 -1200
rect 120 -1652 808 -1228
rect 872 -1652 892 -1228
rect 120 -1680 892 -1652
rect 1132 -1228 1904 -1200
rect 1132 -1652 1820 -1228
rect 1884 -1652 1904 -1228
rect 1132 -1680 1904 -1652
<< via3 >>
rect -1216 1228 -1152 1652
rect -204 1228 -140 1652
rect 808 1228 872 1652
rect 1820 1228 1884 1652
rect -1216 508 -1152 932
rect -204 508 -140 932
rect 808 508 872 932
rect 1820 508 1884 932
rect -1216 -212 -1152 212
rect -204 -212 -140 212
rect 808 -212 872 212
rect 1820 -212 1884 212
rect -1216 -932 -1152 -508
rect -204 -932 -140 -508
rect 808 -932 872 -508
rect 1820 -932 1884 -508
rect -1216 -1652 -1152 -1228
rect -204 -1652 -140 -1228
rect 808 -1652 872 -1228
rect 1820 -1652 1884 -1228
<< mimcap >>
rect -1864 1600 -1464 1640
rect -1864 1280 -1824 1600
rect -1504 1280 -1464 1600
rect -1864 1240 -1464 1280
rect -852 1600 -452 1640
rect -852 1280 -812 1600
rect -492 1280 -452 1600
rect -852 1240 -452 1280
rect 160 1600 560 1640
rect 160 1280 200 1600
rect 520 1280 560 1600
rect 160 1240 560 1280
rect 1172 1600 1572 1640
rect 1172 1280 1212 1600
rect 1532 1280 1572 1600
rect 1172 1240 1572 1280
rect -1864 880 -1464 920
rect -1864 560 -1824 880
rect -1504 560 -1464 880
rect -1864 520 -1464 560
rect -852 880 -452 920
rect -852 560 -812 880
rect -492 560 -452 880
rect -852 520 -452 560
rect 160 880 560 920
rect 160 560 200 880
rect 520 560 560 880
rect 160 520 560 560
rect 1172 880 1572 920
rect 1172 560 1212 880
rect 1532 560 1572 880
rect 1172 520 1572 560
rect -1864 160 -1464 200
rect -1864 -160 -1824 160
rect -1504 -160 -1464 160
rect -1864 -200 -1464 -160
rect -852 160 -452 200
rect -852 -160 -812 160
rect -492 -160 -452 160
rect -852 -200 -452 -160
rect 160 160 560 200
rect 160 -160 200 160
rect 520 -160 560 160
rect 160 -200 560 -160
rect 1172 160 1572 200
rect 1172 -160 1212 160
rect 1532 -160 1572 160
rect 1172 -200 1572 -160
rect -1864 -560 -1464 -520
rect -1864 -880 -1824 -560
rect -1504 -880 -1464 -560
rect -1864 -920 -1464 -880
rect -852 -560 -452 -520
rect -852 -880 -812 -560
rect -492 -880 -452 -560
rect -852 -920 -452 -880
rect 160 -560 560 -520
rect 160 -880 200 -560
rect 520 -880 560 -560
rect 160 -920 560 -880
rect 1172 -560 1572 -520
rect 1172 -880 1212 -560
rect 1532 -880 1572 -560
rect 1172 -920 1572 -880
rect -1864 -1280 -1464 -1240
rect -1864 -1600 -1824 -1280
rect -1504 -1600 -1464 -1280
rect -1864 -1640 -1464 -1600
rect -852 -1280 -452 -1240
rect -852 -1600 -812 -1280
rect -492 -1600 -452 -1280
rect -852 -1640 -452 -1600
rect 160 -1280 560 -1240
rect 160 -1600 200 -1280
rect 520 -1600 560 -1280
rect 160 -1640 560 -1600
rect 1172 -1280 1572 -1240
rect 1172 -1600 1212 -1280
rect 1532 -1600 1572 -1280
rect 1172 -1640 1572 -1600
<< mimcapcontact >>
rect -1824 1280 -1504 1600
rect -812 1280 -492 1600
rect 200 1280 520 1600
rect 1212 1280 1532 1600
rect -1824 560 -1504 880
rect -812 560 -492 880
rect 200 560 520 880
rect 1212 560 1532 880
rect -1824 -160 -1504 160
rect -812 -160 -492 160
rect 200 -160 520 160
rect 1212 -160 1532 160
rect -1824 -880 -1504 -560
rect -812 -880 -492 -560
rect 200 -880 520 -560
rect 1212 -880 1532 -560
rect -1824 -1600 -1504 -1280
rect -812 -1600 -492 -1280
rect 200 -1600 520 -1280
rect 1212 -1600 1532 -1280
<< metal4 >>
rect -1716 1601 -1612 1800
rect -1236 1652 -1132 1800
rect -1825 1600 -1503 1601
rect -1825 1280 -1824 1600
rect -1504 1280 -1503 1600
rect -1825 1279 -1503 1280
rect -1716 881 -1612 1279
rect -1236 1228 -1216 1652
rect -1152 1228 -1132 1652
rect -704 1601 -600 1800
rect -224 1652 -120 1800
rect -813 1600 -491 1601
rect -813 1280 -812 1600
rect -492 1280 -491 1600
rect -813 1279 -491 1280
rect -1236 932 -1132 1228
rect -1825 880 -1503 881
rect -1825 560 -1824 880
rect -1504 560 -1503 880
rect -1825 559 -1503 560
rect -1716 161 -1612 559
rect -1236 508 -1216 932
rect -1152 508 -1132 932
rect -704 881 -600 1279
rect -224 1228 -204 1652
rect -140 1228 -120 1652
rect 308 1601 412 1800
rect 788 1652 892 1800
rect 199 1600 521 1601
rect 199 1280 200 1600
rect 520 1280 521 1600
rect 199 1279 521 1280
rect -224 932 -120 1228
rect -813 880 -491 881
rect -813 560 -812 880
rect -492 560 -491 880
rect -813 559 -491 560
rect -1236 212 -1132 508
rect -1825 160 -1503 161
rect -1825 -160 -1824 160
rect -1504 -160 -1503 160
rect -1825 -161 -1503 -160
rect -1716 -559 -1612 -161
rect -1236 -212 -1216 212
rect -1152 -212 -1132 212
rect -704 161 -600 559
rect -224 508 -204 932
rect -140 508 -120 932
rect 308 881 412 1279
rect 788 1228 808 1652
rect 872 1228 892 1652
rect 1320 1601 1424 1800
rect 1800 1652 1904 1800
rect 1211 1600 1533 1601
rect 1211 1280 1212 1600
rect 1532 1280 1533 1600
rect 1211 1279 1533 1280
rect 788 932 892 1228
rect 199 880 521 881
rect 199 560 200 880
rect 520 560 521 880
rect 199 559 521 560
rect -224 212 -120 508
rect -813 160 -491 161
rect -813 -160 -812 160
rect -492 -160 -491 160
rect -813 -161 -491 -160
rect -1236 -508 -1132 -212
rect -1825 -560 -1503 -559
rect -1825 -880 -1824 -560
rect -1504 -880 -1503 -560
rect -1825 -881 -1503 -880
rect -1716 -1279 -1612 -881
rect -1236 -932 -1216 -508
rect -1152 -932 -1132 -508
rect -704 -559 -600 -161
rect -224 -212 -204 212
rect -140 -212 -120 212
rect 308 161 412 559
rect 788 508 808 932
rect 872 508 892 932
rect 1320 881 1424 1279
rect 1800 1228 1820 1652
rect 1884 1228 1904 1652
rect 1800 932 1904 1228
rect 1211 880 1533 881
rect 1211 560 1212 880
rect 1532 560 1533 880
rect 1211 559 1533 560
rect 788 212 892 508
rect 199 160 521 161
rect 199 -160 200 160
rect 520 -160 521 160
rect 199 -161 521 -160
rect -224 -508 -120 -212
rect -813 -560 -491 -559
rect -813 -880 -812 -560
rect -492 -880 -491 -560
rect -813 -881 -491 -880
rect -1236 -1228 -1132 -932
rect -1825 -1280 -1503 -1279
rect -1825 -1600 -1824 -1280
rect -1504 -1600 -1503 -1280
rect -1825 -1601 -1503 -1600
rect -1716 -1800 -1612 -1601
rect -1236 -1652 -1216 -1228
rect -1152 -1652 -1132 -1228
rect -704 -1279 -600 -881
rect -224 -932 -204 -508
rect -140 -932 -120 -508
rect 308 -559 412 -161
rect 788 -212 808 212
rect 872 -212 892 212
rect 1320 161 1424 559
rect 1800 508 1820 932
rect 1884 508 1904 932
rect 1800 212 1904 508
rect 1211 160 1533 161
rect 1211 -160 1212 160
rect 1532 -160 1533 160
rect 1211 -161 1533 -160
rect 788 -508 892 -212
rect 199 -560 521 -559
rect 199 -880 200 -560
rect 520 -880 521 -560
rect 199 -881 521 -880
rect -224 -1228 -120 -932
rect -813 -1280 -491 -1279
rect -813 -1600 -812 -1280
rect -492 -1600 -491 -1280
rect -813 -1601 -491 -1600
rect -1236 -1800 -1132 -1652
rect -704 -1800 -600 -1601
rect -224 -1652 -204 -1228
rect -140 -1652 -120 -1228
rect 308 -1279 412 -881
rect 788 -932 808 -508
rect 872 -932 892 -508
rect 1320 -559 1424 -161
rect 1800 -212 1820 212
rect 1884 -212 1904 212
rect 1800 -508 1904 -212
rect 1211 -560 1533 -559
rect 1211 -880 1212 -560
rect 1532 -880 1533 -560
rect 1211 -881 1533 -880
rect 788 -1228 892 -932
rect 199 -1280 521 -1279
rect 199 -1600 200 -1280
rect 520 -1600 521 -1280
rect 199 -1601 521 -1600
rect -224 -1800 -120 -1652
rect 308 -1800 412 -1601
rect 788 -1652 808 -1228
rect 872 -1652 892 -1228
rect 1320 -1279 1424 -881
rect 1800 -932 1820 -508
rect 1884 -932 1904 -508
rect 1800 -1228 1904 -932
rect 1211 -1280 1533 -1279
rect 1211 -1600 1212 -1280
rect 1532 -1600 1533 -1280
rect 1211 -1601 1533 -1600
rect 788 -1800 892 -1652
rect 1320 -1800 1424 -1601
rect 1800 -1652 1820 -1228
rect 1884 -1652 1904 -1228
rect 1800 -1800 1904 -1652
<< properties >>
string FIXED_BBOX 1132 1200 1612 1680
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 4 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
