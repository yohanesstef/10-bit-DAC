magic
tech sky130A
magscale 1 2
timestamp 1749922348
<< pwell >>
rect -715 -327 715 327
<< mvnmos >>
rect -487 -131 -287 69
rect -229 -131 -29 69
rect 29 -131 229 69
rect 287 -131 487 69
<< mvndiff >>
rect -545 57 -487 69
rect -545 -119 -533 57
rect -499 -119 -487 57
rect -545 -131 -487 -119
rect -287 57 -229 69
rect -287 -119 -275 57
rect -241 -119 -229 57
rect -287 -131 -229 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 229 57 287 69
rect 229 -119 241 57
rect 275 -119 287 57
rect 229 -131 287 -119
rect 487 57 545 69
rect 487 -119 499 57
rect 533 -119 545 57
rect 487 -131 545 -119
<< mvndiffc >>
rect -533 -119 -499 57
rect -275 -119 -241 57
rect -17 -119 17 57
rect 241 -119 275 57
rect 499 -119 533 57
<< mvpsubdiff >>
rect -679 279 679 291
rect -679 245 -571 279
rect 571 245 679 279
rect -679 233 679 245
rect -679 183 -621 233
rect -679 -183 -667 183
rect -633 -183 -621 183
rect 621 183 679 233
rect -679 -233 -621 -183
rect 621 -183 633 183
rect 667 -183 679 183
rect 621 -233 679 -183
rect -679 -245 679 -233
rect -679 -279 -571 -245
rect 571 -279 679 -245
rect -679 -291 679 -279
<< mvpsubdiffcont >>
rect -571 245 571 279
rect -667 -183 -633 183
rect 633 -183 667 183
rect -571 -279 571 -245
<< poly >>
rect -487 141 -287 157
rect -487 107 -471 141
rect -303 107 -287 141
rect -487 69 -287 107
rect -229 141 -29 157
rect -229 107 -213 141
rect -45 107 -29 141
rect -229 69 -29 107
rect 29 141 229 157
rect 29 107 45 141
rect 213 107 229 141
rect 29 69 229 107
rect 287 141 487 157
rect 287 107 303 141
rect 471 107 487 141
rect 287 69 487 107
rect -487 -157 -287 -131
rect -229 -157 -29 -131
rect 29 -157 229 -131
rect 287 -157 487 -131
<< polycont >>
rect -471 107 -303 141
rect -213 107 -45 141
rect 45 107 213 141
rect 303 107 471 141
<< locali >>
rect -667 245 -571 279
rect 571 245 667 279
rect -667 183 -633 245
rect 633 183 667 245
rect -487 107 -471 141
rect -303 107 -287 141
rect -229 107 -213 141
rect -45 107 -29 141
rect 29 107 45 141
rect 213 107 229 141
rect 287 107 303 141
rect 471 107 487 141
rect -533 57 -499 73
rect -533 -135 -499 -119
rect -275 57 -241 73
rect -275 -135 -241 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 241 57 275 73
rect 241 -135 275 -119
rect 499 57 533 73
rect 499 -135 533 -119
rect -667 -245 -633 -183
rect 633 -245 667 -183
rect -667 -279 -571 -245
rect 571 -279 667 -245
<< viali >>
rect -450 107 -324 141
rect -192 107 -66 141
rect 66 107 192 141
rect 324 107 450 141
rect -533 -119 -499 57
rect -275 -119 -241 57
rect -17 -119 17 57
rect 241 -119 275 57
rect 499 -119 533 57
<< metal1 >>
rect -462 141 -312 147
rect -462 107 -450 141
rect -324 107 -312 141
rect -462 101 -312 107
rect -204 141 -54 147
rect -204 107 -192 141
rect -66 107 -54 141
rect -204 101 -54 107
rect 54 141 204 147
rect 54 107 66 141
rect 192 107 204 141
rect 54 101 204 107
rect 312 141 462 147
rect 312 107 324 141
rect 450 107 462 141
rect 312 101 462 107
rect -539 57 -493 69
rect -539 -119 -533 57
rect -499 -119 -493 57
rect -539 -131 -493 -119
rect -281 57 -235 69
rect -281 -119 -275 57
rect -241 -119 -235 57
rect -281 -131 -235 -119
rect -23 57 23 69
rect -23 -119 -17 57
rect 17 -119 23 57
rect -23 -131 23 -119
rect 235 57 281 69
rect 235 -119 241 57
rect 275 -119 281 57
rect 235 -131 281 -119
rect 493 57 539 69
rect 493 -119 499 57
rect 533 -119 539 57
rect 493 -131 539 -119
<< properties >>
string FIXED_BBOX -650 -262 650 262
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
