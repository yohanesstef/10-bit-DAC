magic
tech sky130A
magscale 1 2
timestamp 1749007001
<< xpolycontact >>
rect -141 593 141 1025
rect -141 -1025 141 -593
<< xpolyres >>
rect -141 -593 141 593
<< viali >>
rect -125 610 125 1007
rect -125 -1007 125 -610
<< metal1 >>
rect -131 1007 131 1019
rect -131 610 -125 1007
rect 125 610 131 1007
rect -131 598 131 610
rect -131 -610 131 -598
rect -131 -1007 -125 -610
rect 125 -1007 131 -610
rect -131 -1019 131 -1007
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 6.089 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 8.903k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
