magic
tech sky130A
magscale 1 2
timestamp 1749007001
<< xpolycontact >>
rect -141 449 141 881
rect -141 -881 141 -449
<< xpolyres >>
rect -141 -449 141 449
<< viali >>
rect -125 466 125 863
rect -125 -863 125 -466
<< metal1 >>
rect -131 863 131 875
rect -131 466 -125 863
rect 125 466 131 863
rect -131 454 131 466
rect -131 -466 131 -454
rect -131 -863 -125 -466
rect 125 -863 131 -466
rect -131 -875 131 -863
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 4.654 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 6.868k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
