magic
tech sky130A
magscale 1 2
timestamp 1750150351
<< nwell >>
rect 35082 4 37002 2128
<< mvnsubdiff >>
rect 35148 948 35161 1184
rect 35195 948 35208 1184
rect 36876 945 36889 1188
rect 36923 945 36936 1188
<< mvnsubdiffcont >>
rect 35221 2015 36863 2049
rect 35161 143 35195 1989
rect 36889 143 36923 1989
rect 35221 83 36863 117
<< metal1 >>
rect 35246 948 35306 1184
rect 35334 948 35394 1184
rect 35503 1156 35549 1184
rect 36019 1156 36065 1184
rect 36535 1156 36581 1184
rect 35503 1096 35509 1156
rect 35569 1096 35640 1156
rect 35929 1096 36156 1156
rect 36373 1096 36515 1156
rect 36575 1096 36581 1156
rect 35503 976 35509 1036
rect 35569 976 35640 1036
rect 35929 976 36156 1036
rect 36373 976 36515 1036
rect 36575 976 36581 1036
rect 35503 948 35549 976
rect 36019 948 36065 976
rect 36535 948 36581 976
<< via1 >>
rect 35246 1898 35306 1958
rect 35334 1810 35394 1870
rect 35509 1096 35569 1156
rect 36515 1096 36575 1156
rect 35509 976 35569 1036
rect 36515 976 36575 1036
rect 35246 262 35306 322
rect 35334 174 35394 234
<< metal2 >>
rect 35503 1096 35509 1156
rect 35569 1096 35575 1156
rect 35503 976 35509 1036
rect 35569 976 35575 1036
rect 36012 860 36072 1272
rect 36509 1096 36515 1156
rect 36575 1096 36936 1156
rect 36509 976 36515 1036
rect 36575 976 36936 1036
use cross_pair  cross_pair_0
timestamp 1750150351
transform 1 0 -474 0 1 -879
box 36114 1855 36403 2035
use cross_pair  cross_pair_1
timestamp 1750150351
transform 1 0 42 0 1 -879
box 36114 1855 36403 2035
use dp_pmos_4  dp_pmos_4_0
timestamp 1749915489
transform 1 0 35637 0 1 1105
box -555 13 1365 1023
use dp_pmos_4  dp_pmos_4_1
timestamp 1749915489
transform 1 0 35637 0 -1 1027
box -555 13 1365 1023
<< labels >>
flabel metal1 s 35246 1041 35246 1041 4 FreeSans 320 90 0 0 P_IN
port 0 se
flabel metal1 s 35334 1041 35334 1041 4 FreeSans 320 90 0 0 N_IN
port 1 se
flabel metal2 s 35966 1298 35966 1298 3 FreeSans 320 0 0 0 I_HEAD
port 4 e
flabel locali s 35161 2049 35161 2049 4 FreeSans 320 0 0 0 VPB
port 5 se
flabel metal1 s 36455 1126 36455 1126 7 FreeSans 320 0 0 0 I_OPA
port 2 w
flabel metal1 s 36455 1005 36455 1005 7 FreeSans 320 0 0 0 I_OPB
port 3 w
<< end >>
