** sch_path: /home/yohanes/10-bit-DAC/xschem/cm_pcell1.sch
.subckt cm_pcell1 G1 io0 io1 io2 ho0 ho1 ho2 ho3 ho4 VDDA
*.PININFO G1:I io[0..2]:O VDDA:I ho[0..4]:O
XM1 io0 G1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1.8 nf=1 m=20
XM2 io1 G1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1.8 nf=1 m=20
XM3 io2 G1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1.8 nf=1 m=8
XM4 ho0 G1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1.8 nf=1 m=2
XM6 ho2 G1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1.8 nf=1 m=4
XM7 ho3 G1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1.8 nf=1 m=8
XM8 ho4 G1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1.8 nf=1 m=16
XM5 ho1 G1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1.8 nf=1 m=2
XM9 VDDA VDDA VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1.8 nf=1 m=16
.ends
