magic
tech sky130A
magscale 1 2
timestamp 1750060524
<< metal2 >>
rect -34 153 718 213
use cm_ncell_1  cm_ncell_1_0
timestamp 1750060524
transform 1 0 19 0 1 -4
box -23 -7 293 227
use cm_ncell_1  cm_ncell_1_1
timestamp 1750060524
transform 1 0 395 0 1 -4
box -23 -7 293 227
<< end >>
