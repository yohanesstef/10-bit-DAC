magic
tech sky130A
magscale 1 2
timestamp 1749624948
<< error_p >>
rect -204 198 204 202
rect -204 -130 -174 198
rect -138 132 138 136
rect -138 -64 -108 132
rect 108 -64 138 132
rect 174 -130 204 198
<< nwell >>
rect -174 -164 174 198
<< mvpmos >>
rect -80 -64 80 136
<< mvpdiff >>
rect -138 124 -80 136
rect -138 -52 -126 124
rect -92 -52 -80 124
rect -138 -64 -80 -52
rect 80 124 138 136
rect 80 -52 92 124
rect 126 -52 138 124
rect 80 -64 138 -52
<< mvpdiffc >>
rect -126 -52 -92 124
rect 92 -52 126 124
<< poly >>
rect -80 136 80 162
rect -80 -111 80 -64
rect -80 -145 -64 -111
rect 64 -145 80 -111
rect -80 -161 80 -145
<< polycont >>
rect -64 -145 64 -111
<< locali >>
rect -126 124 -92 140
rect -126 -68 -92 -52
rect 92 124 126 140
rect 92 -68 126 -52
rect -80 -145 -64 -111
rect 64 -145 80 -111
<< viali >>
rect -126 -52 -92 124
rect 92 -52 126 124
rect -64 -145 64 -111
<< metal1 >>
rect -132 124 -86 136
rect -132 -52 -126 124
rect -92 -52 -86 124
rect -132 -64 -86 -52
rect 86 124 132 136
rect 86 -52 92 124
rect 126 -52 132 124
rect 86 -64 132 -52
rect -76 -111 76 -105
rect -76 -145 -64 -111
rect 64 -145 76 -111
rect -76 -151 76 -145
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
