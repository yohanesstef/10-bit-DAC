magic
tech sky130A
magscale 1 2
timestamp 1750060524
<< error_s >>
rect -1843 859 -1837 865
rect -1789 859 -1783 865
rect -339 859 -333 865
rect -285 859 -279 865
rect -1849 853 -1843 859
rect -1783 853 -1777 859
rect -345 853 -339 859
rect -279 853 -273 859
rect -1849 799 -1843 805
rect -1783 799 -1777 805
rect -345 799 -339 805
rect -279 799 -273 805
rect -1843 793 -1837 799
rect -1789 793 -1783 799
rect -339 793 -333 799
rect -285 793 -279 799
rect -2595 683 -2589 689
rect -2541 683 -2535 689
rect -1091 683 -1085 689
rect -1037 683 -1031 689
rect -2601 677 -2595 683
rect -2535 677 -2529 683
rect -1097 677 -1091 683
rect -1031 677 -1025 683
rect -2601 623 -2595 629
rect -2535 623 -2529 629
rect -1097 623 -1091 629
rect -1031 623 -1025 629
rect -2595 617 -2589 623
rect -2541 617 -2535 623
rect -1091 617 -1085 623
rect -1037 617 -1031 623
rect -527 595 -521 601
rect -473 595 -467 601
rect -533 589 -527 595
rect -467 589 -461 595
rect -533 535 -527 541
rect -467 535 -461 541
rect -527 529 -521 535
rect -473 529 -467 535
rect -1467 507 -1461 513
rect -1413 507 -1407 513
rect -1473 501 -1467 507
rect -1407 501 -1401 507
rect -1473 447 -1467 453
rect -1407 447 -1401 453
rect -1467 441 -1461 447
rect -1413 441 -1407 447
rect -2219 419 -2213 425
rect -2165 419 -2159 425
rect -2225 413 -2219 419
rect -2159 413 -2153 419
rect -2225 359 -2219 365
rect -2159 359 -2153 365
rect -2219 353 -2213 359
rect -2165 353 -2159 359
<< metal1 >>
rect -1849 799 -1843 859
rect -1783 799 -1777 859
rect -345 799 -339 859
rect -279 799 -273 859
rect -1843 573 -1783 799
rect -527 595 -467 601
rect -339 573 -279 799
rect -1473 447 -1467 507
rect -1407 447 -1401 507
rect -527 469 -467 535
rect -604 409 -467 469
<< via1 >>
rect -1843 799 -1783 859
rect -339 799 -279 859
rect -2595 623 -2535 683
rect -1091 623 -1031 683
rect -527 535 -467 595
rect -1467 447 -1407 507
rect -2219 359 -2159 419
use cm_ncell1_cell  cm_ncell1_cell_0
timestamp 1750060524
transform -1 0 137 0 1 -9
box -12 -4 3580 1064
<< end >>
