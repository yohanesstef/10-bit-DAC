magic
tech sky130A
magscale 1 2
timestamp 1749890363
<< error_s >>
rect 1156 983 1162 989
rect 1210 983 1216 989
rect 2660 983 2666 989
rect 2714 983 2720 989
rect 4164 983 4170 989
rect 4218 983 4224 989
rect 1150 977 1156 983
rect 1216 977 1222 983
rect 2654 977 2660 983
rect 2720 977 2726 983
rect 4158 977 4164 983
rect 4224 977 4230 983
rect 1150 923 1156 929
rect 1216 923 1222 929
rect 2654 923 2660 929
rect 2720 923 2726 929
rect 4158 923 4164 929
rect 4224 923 4230 929
rect 1156 917 1162 923
rect 1210 917 1216 923
rect 2660 917 2666 923
rect 2714 917 2720 923
rect 4164 917 4170 923
rect 4218 917 4224 923
rect 1908 895 1914 901
rect 1962 895 1968 901
rect 3412 895 3418 901
rect 3466 895 3472 901
rect 1902 889 1908 895
rect 1968 889 1974 895
rect 3406 889 3412 895
rect 3472 889 3478 895
rect 1902 835 1908 841
rect 1968 835 1974 841
rect 3406 835 3412 841
rect 3472 835 3478 841
rect 1908 829 1914 835
rect 1962 829 1968 835
rect 3412 829 3418 835
rect 3466 829 3472 835
rect 2284 631 2290 637
rect 2338 631 2344 637
rect 2278 625 2284 631
rect 2344 625 2350 631
rect 2278 571 2284 577
rect 2344 571 2350 577
rect 2284 565 2290 571
rect 2338 565 2344 571
rect 839 543 845 549
rect 893 543 899 549
rect 1532 543 1538 549
rect 1586 543 1592 549
rect 3036 543 3042 549
rect 3090 543 3096 549
rect 833 537 839 543
rect 899 537 905 543
rect 1526 537 1532 543
rect 1592 537 1598 543
rect 3030 537 3036 543
rect 3096 537 3102 543
rect 833 483 839 489
rect 899 483 905 489
rect 1526 483 1532 489
rect 1592 483 1598 489
rect 3030 483 3036 489
rect 3096 483 3102 489
rect 839 477 845 483
rect 893 477 899 483
rect 1532 477 1538 483
rect 1586 477 1592 483
rect 3036 477 3042 483
rect 3090 477 3096 483
rect 3788 455 3794 461
rect 3842 455 3848 461
rect 3782 449 3788 455
rect 3848 449 3854 455
rect 3782 395 3788 401
rect 3848 395 3854 401
rect 3788 389 3794 395
rect 3842 389 3848 395
<< metal1 >>
rect 839 543 899 549
rect 839 477 899 483
<< via1 >>
rect 1156 923 1216 983
rect 2660 923 2720 983
rect 4164 923 4224 983
rect 1908 835 1968 895
rect 3412 835 3472 895
rect 2284 571 2344 631
rect 839 483 899 543
rect 1532 483 1592 543
rect 3036 483 3096 543
rect 3788 395 3848 455
use cm_pcell1_cell  cm_pcell1_cell_0
timestamp 1749890363
transform -1 0 4617 0 1 -4
box -35 -10 4729 1308
<< end >>
