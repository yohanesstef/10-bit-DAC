magic
tech sky130A
magscale 1 2
timestamp 1750207421
<< metal2 >>
rect 1933 804 1943 860
rect 1999 804 2009 860
rect 928 772 1503 774
rect 923 716 933 772
rect 989 716 1503 772
rect 928 714 1503 716
rect 1298 628 1308 684
rect 1364 628 1374 684
rect 2059 540 2069 596
rect 2125 540 2135 596
rect 923 -214 933 -158
rect 989 -214 999 -158
rect 1933 -214 1943 -158
rect 1999 -214 2009 -158
rect 797 -302 807 -246
rect 863 -302 873 -246
rect 2059 -302 2069 -246
rect 2125 -302 2135 -246
rect 1298 -854 1308 -798
rect 1364 -854 1374 -798
<< via2 >>
rect 1943 804 1999 860
rect 933 716 989 772
rect 1308 628 1364 684
rect 2069 540 2125 596
rect 807 452 863 508
rect 933 -214 989 -158
rect 1943 -214 1999 -158
rect 807 -302 863 -246
rect 2069 -302 2125 -246
rect 1308 -854 1364 -798
<< metal3 >>
rect 1938 860 2004 870
rect 1938 804 1943 860
rect 1999 804 2004 860
rect 928 772 994 782
rect 928 716 933 772
rect 989 716 994 772
rect 802 508 868 514
rect 802 452 807 508
rect 863 452 868 508
rect 802 -246 868 452
rect 928 -158 994 716
rect 928 -214 933 -158
rect 989 -214 994 -158
rect 928 -224 994 -214
rect 1303 684 1369 694
rect 1303 628 1308 684
rect 1364 628 1369 684
rect 802 -302 807 -246
rect 863 -302 868 -246
rect 802 -312 868 -302
rect 1303 -798 1369 628
rect 1938 -158 2004 804
rect 1938 -214 1943 -158
rect 1999 -214 2004 -158
rect 1938 -224 2004 -214
rect 2064 596 2130 606
rect 2064 540 2069 596
rect 2125 540 2130 596
rect 2064 -246 2130 540
rect 2064 -302 2069 -246
rect 2125 -302 2130 -246
rect 2064 -312 2130 -302
rect 1303 -854 1308 -798
rect 1364 -854 1369 -798
rect 1303 -864 1369 -854
use cm2_pcell1  cm2_pcell1_0
timestamp 1750206734
transform 1 0 -1957 0 1 -1663
box 1957 1661 4889 2977
use cm2_pcell2  cm2_pcell2_0
timestamp 1750166469
transform 1 0 -1957 0 1 -3145
box 1803 1303 5043 3335
<< labels >>
flabel metal2 s 1565 -856 1625 -796 0 FreeSans 320 0 0 0 D0
port 0 nsew
flabel metal2 s 1060 -680 1120 -620 0 FreeSans 320 0 0 0 D1
port 1 nsew
flabel metal2 s 555 -944 615 -884 0 FreeSans 320 0 0 0 D3
port 3 nsew
flabel metal2 s 684 -1032 744 -972 0 FreeSans 320 0 0 0 D4
port 4 nsew
flabel metal2 s 1258 -757 1299 -723 0 FreeSans 320 0 0 0 D2
port 2 nsew
flabel locali s -75 -1763 -41 -1729 0 FreeSans 320 0 0 0 VDDA
port 5 nsew
<< end >>
