* PEX produced on Thu Jun 26 04:02:24 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from top_digital_cell.ext - technology: sky130A

.subckt top_digital_posim DIN0 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 DIN9 VBPLV VBNLV
+ VBPDEC VBNDEC b[0] b[1] b[2] b[3] b[4] b[5] b[6] bb[0] bb[1] bb[2] bb[3] bb[4] bb[5]
+ bb[6] dec0[0] dec0[1] dec0[2] dec0[3] dec1[0] dec1[1] dec1[2] dec1[3] dec2[0] dec2[1]
+ dec2[2] dec2[3] dec2b[0] dec2b[1] dec2b[2] dec2b[3] SH[1] SH[2] SH[3] SH[4] VDD
+ VDDH GND
X0 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t4 GND.t273 GND.t272 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_24840_n1428.t1 decoder_3_0/decoder_2to4_2.bb[0].t2 GND.t36 GND.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_16484_n199.t1 VBPLV.t0 VDDH.t127 VDDH.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X3 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t1 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t4 GND.t110 GND.t109 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 VDDH.t12 VBPDEC.t0 a_22706_943.t0 VDDH.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X5 a_13908_n296.t1 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t2 a_14504_n199.t0 VDDH.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X6 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t5 VDD.t161 VDD.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t3 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t5 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 GND.t69 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t4 a_20048_n709.t0 GND.t68 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X9 a_17344_n1619.t0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t4 GND.t94 GND.t93 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X10 dcell_lv_0.b[8].t3 dcell_lv_0.bb[8].t4 GND.t91 GND.t90 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VDD.t169 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t4 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 VDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 VDDH.t125 VBPLV.t1 a_17038_n199.t1 VDDH.t124 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X13 dcell_lv_0.b[8].t1 dcell_lv_0.bb[8].t5 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t4 VDD.t57 VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t3 decoder_3_0/decoder_2to4_1.bb[1].t4 a_7030_204.t1 GND.t18 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X16 VDDH.t13 VBPDEC.t1 a_23732_943.t1 VDDH.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X17 GND.t338 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t4 a_16088_n709.t0 GND.t337 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X18 a_23732_943.t0 dec1[0].t2 a_23732_685.t0 VDDH.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X19 dcell_lv_0.logic_shift_seg2_0.x7.Y.t2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t4 a_6682_n1748.t1 GND.t201 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_18858_n296.t0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t2 a_19454_n199.t0 VDDH.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X21 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t2 dcell_lv_0.seg_selector_logic_0.x2/x4.A.t3 a_7766_n660.t1 GND.t86 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X22 a_16048_n199.t0 a_15888_n296.t2 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t0 VDDH.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X23 a_24472_685.t0 dec0[2].t2 a_24472_427.t1 VDDH.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X24 a_13118_n709.t1 VBNLV.t0 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t1 GND.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X25 VDD.t119 dcell_lv_0.seg_selector_logic_0.x2/x4.A.t4 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t1 VDD.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X26 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t0 dcell_lv_0.seg_selector_logic_0.x1/x3.B.t3 GND.t169 GND.t168 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 a_25156_427.t1 dec0[2].t3 dec0[3].t1 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X28 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t4 VDD.t181 VDD.t180 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X29 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t1 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t3 GND.t8 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X30 dcell_lv_0.seg_selector_logic_0.x1/x3.A.t2 decoder_3_0/decoder_2to4_1.bb[1].t5 a_7510_428.t1 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 b[2].t1 bb[2].t2 VDDH.t59 VDDH.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X32 a_13908_n296.t0 VBNLV.t1 a_14374_n1619.t0 GND.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X33 SH[1].t1 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t2 VDDH.t80 VDDH.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X34 a_7786_428.t0 dcell_lv_0.bb[8].t6 GND.t154 GND.t153 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X35 bb[3].t1 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t2 VDDH.t72 VDDH.t71 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X36 decoder_3_0/decoder_2to4_2.bb[0].t1 decoder_3_0/decoder_2to4_2.b[0].t4 VDD.t199 VDD.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X37 b[3].t1 bb[3].t2 VDDH.t131 VDDH.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X38 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t1 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t3 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X39 a_7130_n1748.t0 dcell_lv_0.logic_shift_seg2_0.x6.Y.t3 a_7046_n1748.t1 GND.t333 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X40 GND.t320 DIN6.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t2 GND.t319 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X41 dcell_lv_0.logic_shift_seg2_0.x7.Y.t0 dcell_lv_0.b[8].t4 VDD.t120 VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X42 bb[4].t1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t2 VDDH.t42 VDDH.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X43 b[4].t1 bb[4].t2 VDDH.t16 VDDH.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X44 VDD.t201 decoder_3_0/decoder_2to4_2.b[0].t5 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 VDD.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X45 VDD.t213 DIN6.t1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t3 VDD.t212 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X46 decoder_3_0/decoder_2to4_2.b[0].t1 dcell_lv_0.logic_shift_seg2_0.x8.Y.t4 a_7130_n1748.t1 GND.t218 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X47 a_19324_n1619.t0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t5 GND.t107 GND.t106 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X48 bb[5].t1 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t3 VDDH.t64 VDDH.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X49 b[5].t1 bb[5].t2 VDDH.t33 VDDH.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X50 a_6866_n660.t1 dcell_lv_0.bb[9].t4 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X51 dcell_lv_0.logic_shift_seg2_0.x4.B.t2 dcell_lv_0.b[9].t4 VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X52 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 decoder_3_0/decoder_2to4_2.bb[1].t2 a_24288_n1428.t0 GND.t221 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X53 a_21282_685.t1 dec2[2].t2 a_21282_427.t0 VDDH.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X54 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t0 DIN2.t0 GND.t34 GND.t33 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X55 a_13384_n1619.t1 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t3 GND.t172 GND.t171 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X56 GND.t313 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 a_22669_n395.t1 GND.t312 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X57 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t2 dcell_lv_0.bb[9].t5 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X58 GND.t230 decoder_3_0/decoder_2to4_1.bb[1].t6 decoder_3_0/decoder_2to4_1.b[1].t3 GND.t229 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X59 SH[1].t0 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t3 GND.t25 GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X60 a_7322_n884.t1 dcell_lv_0.logic_shift_seg2_0.x4.C.t3 GND.t59 GND.t58 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X61 a_17078_n709.t1 VBNLV.t2 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t1 GND.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X62 a_19848_n296.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t2 a_20444_n199.t0 VDDH.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X63 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t1 DIN2.t1 VDD.t117 VDD.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X64 a_7046_n1748.t0 dcell_lv_0.logic_shift_seg2_0.x7.Y.t3 GND.t174 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X65 a_22706_685.t0 dec1[2].t2 a_22706_427.t0 VDDH.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X66 VDD.t137 decoder_3_0/decoder_2to4_1.bb[1].t7 decoder_3_0/decoder_2to4_1.b[1].t1 VDD.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X67 a_7510_428.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t5 GND.t71 GND.t70 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X68 SH[2].t0 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t2 GND.t21 GND.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X69 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t1 DIN6.t2 GND.t96 GND.t95 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X70 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 decoder_3_0/decoder_2to4_2.b[0].t6 a_25116_n1428.t1 GND.t297 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X71 VDDH.t123 VBPLV.t2 a_14068_n199.t1 VDDH.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X72 dcell_lv_0.logic_shift_seg2_0.x4.A.t2 dcell_lv_0.b[9].t5 a_6406_n884.t1 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X73 a_21992_n1428.t1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t6 GND.t271 GND.t270 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X74 GND.t234 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t2 a_12128_n709.t0 GND.t233 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X75 a_12524_n199.t1 VBPLV.t3 VDDH.t121 VDDH.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X76 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t0 DIN6.t3 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X77 b[2].t0 bb[2].t3 GND.t181 GND.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X78 VDD.t43 decoder_3_0/decoder_2to4_1.b[1].t4 dcell_lv_0.logic_shift_seg2_0.x4.C.t0 VDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X79 a_17868_n296.t1 VBNLV.t3 a_18334_n1619.t0 GND.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X80 a_24288_n1428.t1 decoder_3_0/decoder_2to4_2.bb[0].t3 GND.t38 GND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X81 VDD.t35 decoder_3_0/decoder_2to4_2.b[1].t4 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 VDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X82 a_13078_n199.t0 a_12918_n296.t2 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t0 VDDH.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X83 bb[3].t0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t3 GND.t261 GND.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X84 a_7690_n1748.t0 dcell_lv_0.bb[8].t7 GND.t156 GND.t155 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X85 b[3].t0 bb[3].t3 GND.t203 GND.t202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X86 decoder_3_0/decoder_2to4_1.b[1].t2 decoder_3_0/decoder_2to4_1.bb[1].t8 GND.t73 GND.t72 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X87 a_25142_n983.t1 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 GND.t263 GND.t262 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X88 a_24472_427.t0 dec0[3].t2 dec0[1].t1 VDDH.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X89 bb[4].t0 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t3 GND.t134 GND.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X90 GND.t269 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t7 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t0 GND.t268 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X91 b[4].t0 bb[4].t3 GND.t12 GND.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X92 decoder_3_0/decoder_2to4_1.b[1].t0 decoder_3_0/decoder_2to4_1.bb[1].t9 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X93 a_17474_n199.t1 VBPLV.t4 VDDH.t119 VDDH.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X94 a_25116_n1428.t0 decoder_3_0/decoder_2to4_2.b[1].t5 GND.t57 GND.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X95 bb[5].t0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t4 GND.t239 GND.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X96 VDD.t159 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t8 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t2 VDD.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X97 b[5].t0 bb[5].t3 GND.t329 GND.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X98 VDDH.t7 dec2[0].t2 dec2b[0].t1 VDDH.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X99 a_22294_n983.t0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 GND.t82 GND.t81 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X100 GND.t158 dcell_lv_0.bb[8].t8 dcell_lv_0.b[8].t2 GND.t157 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X101 a_14898_n296.t1 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t2 a_15494_n199.t1 VDDH.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X102 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t1 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t5 GND.t125 GND.t124 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X103 VDD.t86 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t6 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t1 VDD.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X104 VDD.t222 dcell_lv_0.bb[8].t9 dcell_lv_0.b[8].t0 VDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X105 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t0 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t6 VDD.t170 VDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X106 a_18334_n1619.t1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t5 GND.t183 GND.t182 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X107 a_7050_n884.t1 dcell_lv_0.b[9].t6 GND.t243 GND.t242 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X108 dec1[1].t0 VBNDEC.t0 a_23006_n983.t0 GND.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X109 VDDH.t117 VBPLV.t5 a_18028_n199.t1 VDDH.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X110 VDD.t103 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t5 dcell_lv_0.seg_selector_logic_0.x4/x3.B.t1 VDD.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X111 a_24130_943.t0 dec0[1].t2 a_24130_685.t0 VDDH.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X112 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t6 a_21992_n1428.t0 GND.t170 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X113 VDD.t45 decoder_3_0/decoder_2to4_1.b[1].t5 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 VDD.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X114 VDDH.t30 VBPDEC.t2 a_21624_943.t1 VDDH.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X115 decoder_3_0/decoder_2to4_2.b[1].t3 dcell_lv_0.logic_shift_seg2_0.x4.A.t3 a_7406_n884.t1 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X116 a_9948_n296.t1 VBNLV.t4 a_10414_n1619.t1 GND.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X117 a_21966_685.t0 dec2[1].t2 a_21966_427.t1 VDDH.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X118 GND.t67 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t4 a_17078_n709.t0 GND.t66 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X119 a_17038_n199.t0 a_16878_n296.t2 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t0 VDDH.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X120 a_21282_427.t1 dec2[3].t2 dec2[0].t0 VDDH.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X121 a_7030_204.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t6 a_6946_204.t1 GND.t195 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X122 a_14108_n709.t1 VBNLV.t5 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t1 GND.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X123 GND.t225 DIN5.t0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t2 GND.t224 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X124 a_7766_n660.t0 dcell_lv_0.seg_selector_logic_0.x2/x4.B.t3 a_7682_n660.t0 GND.t276 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X125 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t3 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t5 GND.t179 GND.t178 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X126 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t7 a_7314_n660.t0 GND.t167 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X127 VDD.t237 DIN5.t1 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t3 VDD.t236 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X128 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t0 dcell_lv_0.seg_selector_logic_0.x2/x4.B.t4 VDD.t115 VDD.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X129 a_22706_427.t1 dec1[3].t2 dec1[0].t1 VDDH.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X130 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t5 a_21440_n1428.t0 GND.t296 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X131 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t6 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X132 a_14898_n296.t0 VBNLV.t6 a_15364_n1619.t0 GND.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X133 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t8 VDD.t163 VDD.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X134 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t9 VDD.t165 VDD.t164 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X135 VDD.t99 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t7 dcell_lv_0.logic_shift_seg2_0.x7.Y.t1 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X136 bb[0].t1 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t3 VDDH.t51 VDDH.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X137 b[0].t1 bb[0].t2 VDDH.t66 VDDH.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X138 dcell_lv_0.seg_selector_logic_0.x4/x3.B.t0 decoder_3_0/decoder_2to4_1.b[1].t6 VDD.t215 VDD.t214 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X139 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 decoder_3_0/decoder_2to4_2.bb[0].t4 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X140 VDDH.t115 VBPLV.t6 a_10108_n199.t1 VDDH.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X141 VDD.t41 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t8 dcell_lv_0.logic_shift_seg2_0.x4.B.t1 VDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X142 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t1 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t5 a_7326_204.t0 GND.t316 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X143 a_22308_943.t0 dec2[0].t3 a_22308_685.t1 VDDH.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X144 bb[1].t1 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t3 VDDH.t78 VDDH.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X145 b[1].t1 bb[1].t2 VDDH.t56 VDDH.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X146 GND.t251 DIN2.t2 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t2 GND.t250 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X147 a_23048_685.t1 dec1[2].t3 a_23048_427.t0 VDDH.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X148 dec2[0].t1 VBNDEC.t1 a_21245_n395.t1 GND.t258 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X149 VDD.t141 dcell_lv_0.b[9].t7 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t3 VDD.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X150 bb[2].t1 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t2 VDDH.t68 VDDH.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X151 VDD.t122 dcell_lv_0.b[8].t5 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t1 VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X152 VDD.t147 DIN2.t3 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t3 VDD.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X153 VDD.t228 dcell_lv_0.logic_shift_seg2_0.x6.Y.t4 decoder_3_0/decoder_2to4_2.b[0].t3 VDD.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X154 a_7598_n660.t0 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t4 GND.t209 GND.t208 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X155 a_23390_943.t0 dec1[0].t3 a_23390_685.t0 VDDH.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X156 a_14374_n1619.t1 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t4 GND.t197 GND.t196 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X157 a_18068_n709.t0 VBNLV.t7 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t1 GND.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X158 a_22864_n1428.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t10 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X159 VDDH.t113 VBPLV.t7 a_15058_n199.t1 VDDH.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X160 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t4 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t5 VDD.t217 VDD.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X161 a_24430_n983.t0 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 GND.t115 GND.t114 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X162 VDD.t5 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t3 a_6862_678.t1 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X163 GND.t84 DIN1.t0 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t3 GND.t83 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X164 decoder_3_0/decoder_2to4_2.b[0].t2 dcell_lv_0.logic_shift_seg2_0.x8.Y.t5 VDD.t124 VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X165 a_24814_943.t1 dec0[0].t2 a_24814_685.t1 VDDH.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X166 a_13514_n199.t1 VBPLV.t8 VDDH.t111 VDDH.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X167 VDD.t139 DIN1.t1 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t1 VDD.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X168 a_18858_n296.t1 VBNLV.t8 a_19324_n1619.t1 GND.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X169 a_7774_n1748.t1 decoder_3_0/decoder_2to4_1.bb[1].t10 a_7690_n1748.t1 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X170 GND.t75 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t2 a_13118_n709.t0 GND.t74 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X171 a_10938_n296.t0 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t3 a_11534_n199.t0 VDDH.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X172 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t0 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t4 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X173 dcell_lv_0.logic_shift_seg2_0.x6.Y.t0 dcell_lv_0.b[8].t6 a_6406_n1748.t0 GND.t53 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X174 a_21582_n983.t1 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 GND.t282 GND.t281 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X175 a_14068_n199.t0 a_13908_n296.t2 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t0 VDDH.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X176 a_23692_n1428.t0 decoder_3_0/decoder_2to4_1.b[1].t7 GND.t325 GND.t324 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X177 a_21966_427.t0 dec2[3].t3 dec2[2].t1 VDDH.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X178 GND.t340 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t5 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t3 GND.t339 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X179 decoder_3_0/decoder_2to4_2.b[0].t0 dcell_lv_0.logic_shift_seg2_0.x7.Y.t4 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X180 bb[0].t0 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t4 GND.t247 GND.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X181 GND.t40 dec2[0].t4 dec2b[0].t0 GND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X182 b[0].t0 bb[0].t3 GND.t241 GND.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X183 dec2[3].t1 VBNDEC.t2 a_22294_n983.t1 GND.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X184 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t2 dcell_lv_0.b[9].t8 VDD.t143 VDD.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X185 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t0 DIN5.t2 GND.t52 GND.t51 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X186 a_18464_n199.t1 VBPLV.t9 VDDH.t109 VDDH.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X187 bb[1].t0 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t4 GND.t142 GND.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X188 VDD.t130 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t6 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t1 VDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X189 b[1].t0 bb[1].t3 GND.t213 GND.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X190 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t4 dcell_lv_0.b[9].t9 VDD.t185 VDD.t184 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X191 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t2 DIN1.t2 GND.t50 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X192 a_15888_n296.t1 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t3 a_16484_n199.t0 VDDH.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X193 VDDH.t44 dec2[2].t3 dec2b[2].t1 VDDH.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X194 a_23732_685.t1 dec1[1].t2 a_23732_427.t1 VDDH.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X195 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t1 DIN5.t3 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X196 bb[2].t0 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t4 GND.t284 GND.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X197 a_21440_n1428.t1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t9 GND.t267 GND.t266 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X198 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t0 DIN1.t3 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X199 dcell_lv_0.bb[9].t2 DIN9.t0 GND.t205 GND.t204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X200 dcell_lv_0.logic_shift_seg2_0.x8.Y.t2 dcell_lv_0.bb[8].t10 VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X201 a_7326_204.t1 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t5 GND.t140 GND.t139 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X202 a_6406_n1748.t1 decoder_3_0/decoder_2to4_1.b[1].t8 GND.t327 GND.t326 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X203 a_21624_943.t0 dec2[0].t5 a_21624_685.t1 VDDH.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X204 VDDH.t107 VBPLV.t10 a_19018_n199.t1 VDDH.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X205 VDD.t195 decoder_3_0/decoder_2to4_2.bb[1].t3 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 VDD.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X206 dcell_lv_0.bb[9].t3 DIN9.t1 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X207 VDD.t49 decoder_3_0/decoder_2to4_1.bb[1].t11 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t2 VDD.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X208 VDDH.t48 dec2[3].t4 dec2b[3].t1 VDDH.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X209 a_6682_n884.t1 dcell_lv_0.b[9].t10 GND.t300 GND.t299 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X210 a_10938_n296.t1 VBNLV.t9 a_11404_n1619.t1 GND.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X211 VDDH.t31 VBPDEC.t3 a_22308_943.t1 VDDH.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X212 bb[6].t1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t3 VDDH.t20 VDDH.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X213 a_10414_n1619.t0 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t2 GND.t275 GND.t274 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X214 a_18028_n199.t0 a_17868_n296.t2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t0 VDDH.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X215 a_23048_427.t1 dec1[3].t3 dec1[1].t1 VDDH.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X216 b[6].t1 bb[6].t2 VDDH.t133 VDDH.t132 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X217 a_7406_n884.t0 dcell_lv_0.logic_shift_seg2_0.x4.B.t3 a_7322_n884.t0 GND.t323 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X218 a_19848_n296.t1 VBNLV.t10 a_20314_n1619.t1 GND.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X219 VDD.t183 decoder_3_0/decoder_2to4_2.b[0].t7 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 VDD.t182 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X220 VDDH.t60 VBPDEC.t4 a_24472_943.t0 VDDH.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X221 GND.t89 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t7 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t1 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X222 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t10 VDD.t157 VDD.t156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X223 GND.t265 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t11 a_18068_n709.t1 GND.t264 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X224 dcell_lv_0.logic_shift_seg2_0.x8.Y.t1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t11 a_7774_n1748.t0 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X225 a_6590_n660.t0 decoder_3_0/decoder_2to4_1.b[1].t9 GND.t291 GND.t290 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X226 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t0 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t4 VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X227 VDD.t67 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t8 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t2 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X228 decoder_3_0/decoder_2to4_2.b[1].t1 dcell_lv_0.logic_shift_seg2_0.x4.C.t4 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X229 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 decoder_3_0/decoder_2to4_2.bb[0].t5 VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X230 dcell_lv_0.seg_selector_logic_0.x2/x4.B.t0 decoder_3_0/decoder_2to4_1.b[1].t10 VDD.t173 VDD.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X231 a_15888_n296.t0 VBNLV.t11 a_16354_n1619.t0 GND.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X232 a_7314_n660.t1 decoder_3_0/decoder_2to4_1.bb[1].t12 a_7230_n660.t1 GND.t42 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X233 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t9 a_23140_n1428.t0 GND.t80 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X234 VDD.t19 decoder_3_0/decoder_2to4_1.bb[1].t13 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t3 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X235 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 decoder_3_0/decoder_2to4_2.b[1].t6 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X236 a_23718_n983.t0 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 GND.t211 GND.t210 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X237 VDDH.t105 VBPLV.t11 a_11098_n199.t0 VDDH.t104 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X238 dcell_lv_0.seg_selector_logic_0.x4/x3.B.t2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t10 a_6590_428.t1 GND.t102 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X239 VDDH.t103 VBPLV.t12 a_20008_n199.t1 VDDH.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X240 a_6862_678.t0 dcell_lv_0.seg_selector_logic_0.x4/x3.B.t3 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t2 VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X241 dec0[1].t0 VBNDEC.t3 a_24430_n983.t1 GND.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X242 GND.t44 DIN8.t0 dcell_lv_0.bb[8].t0 GND.t43 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X243 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t0 dcell_lv_0.b[8].t7 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X244 a_25156_943.t1 dec0[0].t3 a_25156_685.t1 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X245 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 decoder_3_0/decoder_2to4_1.bb[1].t14 a_22864_n1428.t1 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X246 VDD.t231 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t6 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t2 VDD.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X247 VDD.t149 dcell_lv_0.seg_selector_logic_0.x1/x3.A.t3 a_8058_678.t0 VDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X248 bb[6].t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t4 GND.t23 GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X249 b[6].t0 bb[6].t3 GND.t346 GND.t345 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X250 a_19058_n709.t1 VBNLV.t12 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t1 GND.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X251 a_23732_427.t0 dec1[2].t4 dec1[3].t1 VDDH.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X252 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t3 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t12 GND.t138 GND.t137 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X253 a_6406_n884.t0 dcell_lv_0.b[8].t8 GND.t55 GND.t54 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X254 dec0[0].t1 VBNDEC.t4 a_24093_n395.t1 GND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X255 dcell_lv_0.logic_shift_seg2_0.x4.C.t1 decoder_3_0/decoder_2to4_1.b[1].t11 a_7050_n884.t0 GND.t285 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X256 VDD.t21 DIN8.t1 dcell_lv_0.bb[8].t1 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X257 VDD.t88 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t7 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 VDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X258 VDDH.t101 VBPLV.t13 a_16048_n199.t1 VDDH.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X259 a_15364_n1619.t1 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t4 GND.t253 GND.t252 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X260 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t13 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X261 a_14504_n199.t1 VBPLV.t14 VDDH.t99 VDDH.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X262 dec2[1].t0 VBNDEC.t5 a_21582_n983.t0 GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X263 a_24564_n1428.t0 decoder_3_0/decoder_2to4_2.bb[1].t4 GND.t309 GND.t60 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X264 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t11 a_23692_n1428.t1 GND.t103 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X265 GND.t315 dcell_lv_0.bb[9].t6 dcell_lv_0.b[9].t3 GND.t314 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X266 a_11928_n296.t0 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t2 a_12524_n199.t0 VDDH.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X267 a_6314_n660.t1 dcell_lv_0.b[9].t11 GND.t302 GND.t301 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X268 GND.t144 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t6 a_14108_n709.t0 GND.t143 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X269 a_6590_428.t0 decoder_3_0/decoder_2to4_1.b[1].t12 GND.t287 GND.t286 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X270 VDD.t203 dcell_lv_0.bb[9].t7 dcell_lv_0.b[9].t1 VDD.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X271 dcell_lv_0.bb[8].t2 DIN8.t2 GND.t215 GND.t214 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X272 dcell_lv_0.seg_selector_logic_0.x2/x4.A.t0 dcell_lv_0.b[9].t12 VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X273 VDD.t235 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t6 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 VDD.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X274 dcell_lv_0.bb[8].t3 DIN8.t3 VDD.t113 VDD.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X275 a_24130_685.t1 dec0[2].t4 a_24130_427.t1 VDDH.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X276 GND.t27 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 a_24805_n395.t0 GND.t26 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X277 a_10148_n709.t1 VBNLV.t13 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t1 GND.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X278 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t0 dcell_lv_0.b[8].t9 a_6314_428.t0 GND.t76 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X279 a_6946_204.t0 dcell_lv_0.b[8].t10 a_6862_204.t0 GND.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X280 GND.t191 DIN9.t2 dcell_lv_0.bb[9].t0 GND.t190 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X281 a_16878_n296.t0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t4 a_17474_n199.t0 VDDH.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X282 VDD.t90 decoder_3_0/decoder_2to4_1.bb[1].t15 dcell_lv_0.logic_shift_seg2_0.x8.Y.t3 VDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X283 dec0[3].t0 VBNDEC.t6 a_25142_n983.t0 GND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X284 VDD.t39 dcell_lv_0.b[8].t11 dcell_lv_0.logic_shift_seg2_0.x6.Y.t1 VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X285 a_11138_n709.t0 VBNLV.t14 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t1 GND.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X286 VDD.t96 DIN9.t3 dcell_lv_0.bb[9].t1 VDD.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X287 GND.t280 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 a_21957_n395.t0 GND.t279 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X288 GND.t200 dec2[3].t5 dec2b[3].t0 GND.t199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X289 GND.t117 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t14 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t2 GND.t116 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X290 dec1[0].t0 VBNDEC.t7 a_22669_n395.t0 GND.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X291 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t6 a_22268_n1428.t1 GND.t248 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X292 a_23140_n1428.t1 decoder_3_0/decoder_2to4_1.bb[1].t16 GND.t220 GND.t219 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X293 VDD.t133 dcell_lv_0.b[9].t13 dcell_lv_0.logic_shift_seg2_0.x4.A.t1 VDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X294 VDD.t65 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t15 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t0 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X295 a_11928_n296.t1 VBNLV.t15 a_12394_n1619.t1 GND.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X296 decoder_3_0/decoder_2to4_2.bb[1].t0 decoder_3_0/decoder_2to4_2.b[1].t7 GND.t98 GND.t97 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X297 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t1 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t5 GND.t245 GND.t244 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X298 a_24472_943.t1 dec0[0].t4 a_24472_685.t1 VDDH.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X299 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t0 DIN0.t0 GND.t123 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X300 a_19018_n199.t0 a_18858_n296.t2 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t0 VDDH.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X301 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t16 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X302 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t12 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X303 GND.t344 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t7 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t3 GND.t343 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X304 VDD.t205 dcell_lv_0.bb[9].t8 dcell_lv_0.seg_selector_logic_0.x1/x3.B.t1 VDD.t204 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X305 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t3 DIN0.t1 VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X306 a_11404_n1619.t0 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t2 GND.t342 GND.t341 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X307 VDD.t211 dcell_lv_0.logic_shift_seg2_0.x4.B.t4 decoder_3_0/decoder_2to4_2.b[1].t0 VDD.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X308 VDDH.t61 VBPDEC.t5 a_25156_943.t0 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X309 dcell_lv_0.logic_shift_seg2_0.x6.Y.t2 decoder_3_0/decoder_2to4_1.b[1].t13 VDD.t218 VDD.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X310 VDD.t175 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t8 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t0 VDD.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X311 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t7 a_21716_n1428.t1 GND.t249 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X312 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t3 DIN4.t0 GND.t318 GND.t317 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X313 a_23006_n983.t1 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 GND.t232 GND.t231 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X314 a_22308_685.t0 dec2[1].t3 a_22308_427.t1 VDDH.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X315 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t4 dcell_lv_0.b[9].t14 a_6478_204.t1 GND.t226 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X316 a_6314_428.t1 dcell_lv_0.b[9].t15 GND.t304 GND.t303 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X317 GND.t295 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t9 a_19058_n709.t0 GND.t294 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X318 a_6862_204.t1 dcell_lv_0.b[9].t16 GND.t305 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X319 a_22268_n1428.t0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t8 GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X320 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 decoder_3_0/decoder_2to4_1.b[1].t14 VDD.t220 VDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X321 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t2 DIN4.t1 VDD.t187 VDD.t186 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X322 dcell_lv_0.logic_shift_seg2_0.x4.A.t0 dcell_lv_0.b[8].t12 VDD.t191 VDD.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X323 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t13 a_6866_n660.t0 GND.t48 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X324 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t3 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t4 GND.t308 GND.t307 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X325 a_6478_204.t0 dcell_lv_0.b[8].t13 a_6394_204.t0 GND.t306 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X326 GND.t228 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t5 a_10148_n709.t0 GND.t227 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X327 dec1[3].t0 VBNDEC.t8 a_23718_n983.t1 GND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X328 VDD.t153 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t14 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t1 VDD.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X329 VDDH.t36 VBPDEC.t6 a_23390_943.t1 VDDH.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X330 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t1 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t5 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X331 GND.t32 DIN7.t0 decoder_3_0/decoder_2to4_1.bb[1].t0 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X332 a_15098_n709.t0 VBNLV.t16 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t0 GND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X333 a_23390_685.t1 dec1[1].t3 a_23390_427.t0 VDDH.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X334 dcell_lv_0.b[9].t2 dcell_lv_0.bb[9].t9 GND.t185 GND.t184 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X335 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t1 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t10 GND.t322 GND.t321 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X336 dec1[2].t0 VBNDEC.t9 a_23381_n395.t1 GND.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X337 VDDH.t97 VBPLV.t15 a_12088_n199.t1 VDDH.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X338 decoder_3_0/decoder_2to4_2.bb[1].t1 decoder_3_0/decoder_2to4_2.b[1].t8 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X339 VDD.t15 DIN7.t1 decoder_3_0/decoder_2to4_1.bb[1].t1 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X340 dcell_lv_0.logic_shift_seg2_0.x8.Y.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t17 VDD.t61 VDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X341 a_10108_n199.t0 a_9948_n296.t2 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t0 VDDH.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X342 dcell_lv_0.b[9].t0 dcell_lv_0.bb[9].t10 VDD.t94 VDD.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X343 a_10544_n199.t1 VBPLV.t16 VDDH.t95 VDDH.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X344 a_21282_943.t0 dec2[1].t4 a_21282_685.t0 VDDH.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X345 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t2 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t11 VDD.t209 VDD.t208 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X346 VDD.t193 dcell_lv_0.b[8].t14 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t0 VDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X347 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t12 VDD.t155 VDD.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X348 a_21716_n1428.t0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t12 GND.t87 GND.t62 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X349 a_24814_685.t0 dec0[1].t3 a_24814_427.t0 VDDH.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X350 a_24130_427.t0 dec0[3].t3 dec0[0].t0 VDDH.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X351 GND.t85 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t4 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t1 GND.t77 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X352 a_11098_n199.t1 a_10938_n296.t2 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t0 VDDH.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X353 a_20314_n1619.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t15 GND.t257 GND.t256 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X354 a_20048_n709.t1 VBNLV.t17 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t1 GND.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X355 a_22706_943.t1 dec1[1].t4 a_22706_685.t1 VDDH.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X356 VDDH.t24 dec2[1].t5 dec2b[1].t1 VDDH.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X357 a_8058_678.t1 dcell_lv_0.seg_selector_logic_0.x1/x3.B.t4 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t1 VDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X358 VDD.t128 decoder_3_0/decoder_2to4_1.bb[1].t17 dcell_lv_0.seg_selector_logic_0.x1/x3.A.t1 VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X359 GND.t129 DIN4.t2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t1 GND.t128 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X360 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 decoder_3_0/decoder_2to4_2.b[0].t8 a_24564_n1428.t1 GND.t298 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X361 dcell_lv_0.logic_shift_seg2_0.x4.B.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t16 a_6682_n884.t0 GND.t147 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X362 a_15494_n199.t0 VBPLV.t17 VDDH.t93 VDDH.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X363 a_6394_204.t1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t18 a_6310_204.t0 GND.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X364 VDDH.t37 VBPDEC.t7 a_24814_943.t0 VDDH.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X365 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t2 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t7 GND.t223 GND.t222 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X366 a_16354_n1619.t1 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t4 GND.t47 GND.t46 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X367 decoder_3_0/decoder_2to4_2.b[1].t2 dcell_lv_0.logic_shift_seg2_0.x4.A.t4 VDD.t233 VDD.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X368 GND.t105 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 a_24093_n395.t0 GND.t104 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X369 VDD.t33 DIN4.t3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t0 VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X370 dcell_lv_0.seg_selector_logic_0.x1/x3.B.t0 dcell_lv_0.bb[8].t11 VDD.t226 VDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X371 dec0[2].t0 VBNDEC.t10 a_24805_n395.t1 GND.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X372 a_12918_n296.t0 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t2 a_13514_n199.t0 VDDH.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X373 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t0 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t8 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X374 VDDH.t45 VBPDEC.t8 a_21966_943.t1 VDDH.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X375 GND.t311 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 a_21245_n395.t0 GND.t310 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X376 GND.t121 DIN3.t0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t0 GND.t120 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X377 dcell_lv_0.seg_selector_logic_0.x2/x4.B.t2 dcell_lv_0.bb[9].t11 a_6590_n660.t1 GND.t186 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X378 GND.t278 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t6 a_15098_n709.t1 GND.t277 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X379 a_21624_685.t0 dec2[2].t4 a_21624_427.t0 VDDH.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X380 dec2[2].t0 VBNDEC.t11 a_21957_n395.t1 GND.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X381 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t0 dcell_lv_0.seg_selector_logic_0.x4/x3.B.t4 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X382 VDD.t239 DIN3.t1 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t3 VDD.t238 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X383 VDD.t230 dcell_lv_0.bb[9].t12 dcell_lv_0.seg_selector_logic_0.x2/x4.B.t1 VDD.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X384 VDD.t77 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t17 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X385 a_22308_427.t0 dec2[2].t5 dec2[3].t0 VDDH.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X386 decoder_3_0/decoder_2to4_2.bb[0].t0 decoder_3_0/decoder_2to4_2.b[0].t9 GND.t29 GND.t28 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X387 a_17868_n296.t0 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t4 a_18464_n199.t0 VDDH.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X388 SH[2].t1 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t4 VDDH.t75 VDDH.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X389 a_15058_n199.t0 a_14898_n296.t2 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t1 VDDH.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X390 a_6682_n1748.t0 dcell_lv_0.b[8].t15 GND.t164 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X391 a_12128_n709.t1 VBNLV.t18 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t1 GND.t330 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X392 SH[3].t1 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t3 VDDH.t54 VDDH.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X393 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 decoder_3_0/decoder_2to4_2.b[1].t9 a_24840_n1428.t0 GND.t130 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X394 dcell_lv_0.seg_selector_logic_0.x1/x3.A.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t19 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X395 a_6310_204.t1 decoder_3_0/decoder_2to4_1.b[1].t15 GND.t207 GND.t206 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X396 a_23390_427.t1 dec1[3].t4 dec1[2].t1 VDDH.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X397 decoder_3_0/decoder_2to4_1.bb[1].t2 DIN7.t2 GND.t255 GND.t254 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X398 SH[4].t1 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t3 VDDH.t129 VDDH.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X399 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t1 DIN3.t2 GND.t152 GND.t151 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X400 a_19454_n199.t1 VBPLV.t18 VDDH.t91 VDDH.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X401 GND.t293 dec2[2].t6 dec2b[2].t0 GND.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X402 GND.t127 DIN0.t2 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t1 GND.t126 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X403 a_12918_n296.t1 VBNLV.t19 a_13384_n1619.t0 GND.t331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X404 a_21966_943.t0 dec2[0].t6 a_21966_685.t1 VDDH.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X405 VDD.t177 decoder_3_0/decoder_2to4_1.bb[1].t18 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 VDD.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X406 decoder_3_0/decoder_2to4_1.bb[1].t3 DIN7.t3 VDD.t151 VDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X407 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t2 DIN3.t3 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X408 a_20008_n199.t0 a_19848_n296.t2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t0 VDDH.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X409 a_24814_427.t1 dec0[3].t4 dec0[2].t1 VDDH.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X410 VDD.t73 DIN0.t3 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t2 VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X411 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t2 decoder_3_0/decoder_2to4_1.b[1].t16 VDD.t107 VDD.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X412 VDDH.t46 VBPDEC.t9 a_23048_943.t1 VDDH.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X413 SH[3].t0 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t4 GND.t217 GND.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X414 VDD.t82 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t18 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 VDD.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X415 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 decoder_3_0/decoder_2to4_2.bb[1].t5 VDD.t197 VDD.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X416 a_12394_n1619.t0 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t4 GND.t193 GND.t192 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X417 GND.t119 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t7 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t2 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X418 VDDH.t81 VBPDEC.t10 a_24130_943.t1 VDDH.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X419 SH[4].t0 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t4 GND.t335 GND.t334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X420 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t0 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t5 VDD.t98 VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X421 a_7230_n660.t0 dcell_lv_0.b[8].t16 GND.t166 GND.t165 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X422 a_9948_n296.t0 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t4 a_10544_n199.t0 VDDH.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X423 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 decoder_3_0/decoder_2to4_1.b[1].t17 a_23416_n1428.t1 GND.t45 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X424 VDD.t92 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t8 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t0 VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X425 dcell_lv_0.seg_selector_logic_0.x2/x4.A.t2 dcell_lv_0.bb[8].t12 a_6314_n660.t0 GND.t198 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X426 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t0 dcell_lv_0.b[8].t17 VDD.t84 VDD.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X427 a_25156_685.t0 dec0[1].t4 a_25156_427.t0 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X428 a_16088_n709.t1 VBNLV.t20 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t1 GND.t332 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X429 VDDH.t82 VBPDEC.t11 a_21282_943.t1 VDDH.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X430 VDD.t101 dcell_lv_0.bb[8].t13 dcell_lv_0.seg_selector_logic_0.x2/x4.A.t1 VDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X431 GND.t289 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t7 a_11138_n709.t1 GND.t288 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X432 a_7682_n660.t1 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t3 a_7598_n660.t1 GND.t194 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X433 VDDH.t89 VBPLV.t19 a_13078_n199.t1 VDDH.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X434 GND.t146 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t7 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t0 GND.t145 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X435 GND.t132 dcell_lv_0.seg_selector_logic_0.x1/x3.A.t4 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t2 GND.t131 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X436 VDD.t207 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t4 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t3 VDD.t206 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X437 a_23048_943.t0 dec1[0].t4 a_23048_685.t0 VDDH.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X438 a_11534_n199.t1 VBPLV.t20 VDDH.t87 VDDH.t86 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X439 a_21624_427.t1 dec2[3].t6 dec2[1].t1 VDDH.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X440 VDD.t1 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t8 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t2 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X441 a_16878_n296.t1 VBNLV.t21 a_17344_n1619.t1 GND.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X442 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t0 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t6 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X443 GND.t79 dec2[1].t6 dec2b[1].t0 GND.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X444 GND.t136 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 a_23381_n395.t0 GND.t135 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X445 a_20444_n199.t1 VBPLV.t21 VDDH.t85 VDDH.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X446 a_12088_n199.t0 a_11928_n296.t2 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t0 VDDH.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X447 dcell_lv_0.logic_shift_seg2_0.x4.C.t2 dcell_lv_0.b[9].t17 VDD.t189 VDD.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X448 dcell_lv_0.seg_selector_logic_0.x1/x3.B.t2 dcell_lv_0.bb[9].t13 a_7786_428.t1 GND.t336 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X449 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 decoder_3_0/decoder_2to4_1.bb[1].t19 VDD.t179 VDD.t178 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X450 VDD.t167 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t8 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 VDD.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X451 a_23416_n1428.t0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t20 GND.t176 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t11 732.773
R1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t10 229.369
R2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t12 229.369
R3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t8 212.081
R4 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t5 212.081
R5 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 208.964
R6 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 186.001
R7 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t6 157.07
R8 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t9 157.07
R9 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 152.712
R10 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 152.475
R11 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t7 139.78
R12 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t4 139.78
R13 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 96.8352
R14 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 61.346
R15 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t0 26.5955
R16 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t2 26.5955
R17 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t1 24.9236
R18 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t3 24.9236
R19 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 15.8609
R20 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 13.6401
R21 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 12.5445
R22 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 11.2645
R23 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 10.2234
R24 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 9.77342
R25 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 9.65467
R26 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 9.30258
R27 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 6.86092
R28 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 6.1445
R29 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 5.45235
R30 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 5.21532
R31 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 5.04425
R32 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 4.8645
R33 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 4.65505
R34 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 3.0725
R35 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 2.0485
R36 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 1.55202
R37 GND.t236 GND.n530 29070.7
R38 GND.n530 GND.n419 21705.6
R39 GND.n693 GND.n57 14701.8
R40 GND.n692 GND.n691 13398.7
R41 GND.n419 GND.n94 11266
R42 GND.n693 GND.n692 6790.35
R43 GND.n461 GND.n431 4533.07
R44 GND.n505 GND.n431 4533.07
R45 GND.n533 GND.n88 3250.5
R46 GND.n544 GND.n88 3250.5
R47 GND.n544 GND.n82 3250.5
R48 GND.n548 GND.n82 3250.5
R49 GND.n548 GND.n74 3250.5
R50 GND.n559 GND.n74 3250.5
R51 GND.n559 GND.n68 3250.5
R52 GND.n563 GND.n68 3250.5
R53 GND.n566 GND.n563 3250.5
R54 GND.n566 GND.n62 3250.5
R55 GND.n536 GND.n90 3151.5
R56 GND.n542 GND.n90 3151.5
R57 GND.n542 GND.n81 3151.5
R58 GND.n551 GND.n81 3151.5
R59 GND.n551 GND.n77 3151.5
R60 GND.n557 GND.n77 3151.5
R61 GND.n557 GND.n67 3151.5
R62 GND.n569 GND.n67 3151.5
R63 GND.n569 GND.n63 3151.5
R64 GND.n574 GND.n63 3151.5
R65 GND.n691 GND.n690 2730.51
R66 GND.n298 GND.n297 2179.52
R67 GND.n265 GND.n264 2179.52
R68 GND.n284 GND.n283 2179.52
R69 GND.n690 GND.n689 2079.22
R70 GND.n309 GND.n244 1783.49
R71 GND.n122 GND.n106 1644.76
R72 GND.n687 GND.t124 1576.25
R73 GND.n128 GND.n127 1571.43
R74 GND.n145 GND.n144 1571.43
R75 GND.n838 GND.t145 1512.83
R76 GND.n837 GND.t118 1512.83
R77 GND.t339 GND.n12 1512.83
R78 GND.t88 GND.n16 1512.83
R79 GND.t268 GND.n20 1512.83
R80 GND.t343 GND.n24 1512.83
R81 GND.t116 GND.n28 1512.83
R82 GND.t229 GND.n32 1512.83
R83 GND.t157 GND.n36 1512.83
R84 GND.t314 GND.n40 1512.83
R85 GND.n405 GND.n160 1392.92
R86 GND.n387 GND.n386 1392.92
R87 GND.n373 GND.n188 1392.92
R88 GND.n355 GND.n354 1392.92
R89 GND.n341 GND.n216 1392.92
R90 GND.n323 GND.n322 1392.92
R91 GND GND.t63 1360.92
R92 GND GND.t126 1331.72
R93 GND.t83 GND 1331.72
R94 GND.t250 GND 1331.72
R95 GND.t120 GND 1331.72
R96 GND.t128 GND 1331.72
R97 GND.t224 GND 1331.72
R98 GND.t319 GND 1331.72
R99 GND.t31 GND 1331.72
R100 GND.t43 GND 1331.72
R101 GND.t190 GND 1331.72
R102 GND.t131 GND.n61 1213.79
R103 GND.n748 GND.n40 1198.25
R104 GND.n759 GND.n36 1198.25
R105 GND.n770 GND.n32 1198.25
R106 GND.n781 GND.n28 1198.25
R107 GND.n792 GND.n24 1198.25
R108 GND.n803 GND.n20 1198.25
R109 GND.n814 GND.n16 1198.25
R110 GND.n825 GND.n12 1198.25
R111 GND.n837 GND.n836 1198.25
R112 GND.n839 GND.n838 1198.25
R113 GND.n701 GND.n55 1198.25
R114 GND.n700 GND.n57 1198.25
R115 GND.n664 GND.n663 1198.25
R116 GND.n687 GND.n686 1198.25
R117 GND.n662 GND.n661 1198.25
R118 GND.n674 GND.n641 1198.25
R119 GND.n587 GND.n582 1198.25
R120 GND.n604 GND.n588 1198.25
R121 GND.n586 GND.n579 1198.25
R122 GND.n627 GND.n580 1198.25
R123 GND.n712 GND.n52 1198.25
R124 GND.n645 GND.n58 1198.01
R125 GND GND.n430 1173.31
R126 GND.n529 GND 1173.31
R127 GND GND.n507 1173.31
R128 GND GND.n489 1173.31
R129 GND.n487 GND 1173.31
R130 GND.t86 GND 1104.21
R131 GND.n691 GND.n60 1063.62
R132 GND.n689 GND.t188 1007.9
R133 GND.n123 GND.n122 1005.71
R134 GND.n127 GND.n124 1005.71
R135 GND.n146 GND.n145 1005.71
R136 GND.n419 GND.n418 942.273
R137 GND.t199 GND.n106 932.381
R138 GND.n128 GND.t292 932.381
R139 GND.n144 GND.t78 932.381
R140 GND.t39 GND.n94 932.381
R141 GND.n111 GND.n110 900.971
R142 GND.n838 GND.n5 894.915
R143 GND.t145 GND.t109 894.915
R144 GND.t126 GND.t122 894.915
R145 GND.t307 GND.t118 894.915
R146 GND.t49 GND.t83 894.915
R147 GND.t222 GND.t339 894.915
R148 GND.t33 GND.t250 894.915
R149 GND.t178 GND.t88 894.915
R150 GND.t151 GND.t120 894.915
R151 GND.t272 GND.t268 894.915
R152 GND.t317 GND.t128 894.915
R153 GND.t321 GND.t343 894.915
R154 GND.t51 GND.t224 894.915
R155 GND.t137 GND.t116 894.915
R156 GND.t95 GND.t319 894.915
R157 GND.t72 GND.t229 894.915
R158 GND.t254 GND.t31 894.915
R159 GND.t90 GND.t157 894.915
R160 GND.t214 GND.t43 894.915
R161 GND.t184 GND.t314 894.915
R162 GND.t204 GND.t190 894.915
R163 GND GND.t124 842.913
R164 GND GND.n837 799.032
R165 GND.n12 GND 799.032
R166 GND.n16 GND 799.032
R167 GND.n20 GND 799.032
R168 GND.n24 GND 799.032
R169 GND.n28 GND 799.032
R170 GND.n32 GND 799.032
R171 GND.n36 GND 799.032
R172 GND.n40 GND 799.032
R173 GND.t167 GND.t30 775.48
R174 GND.n689 GND.n688 744.027
R175 GND.t109 GND 713.802
R176 GND.t122 GND 713.802
R177 GND GND.t307 713.802
R178 GND GND.t49 713.802
R179 GND GND.t222 713.802
R180 GND GND.t33 713.802
R181 GND GND.t178 713.802
R182 GND GND.t151 713.802
R183 GND GND.t272 713.802
R184 GND GND.t317 713.802
R185 GND GND.t321 713.802
R186 GND GND.t51 713.802
R187 GND GND.t137 713.802
R188 GND GND.t95 713.802
R189 GND GND.t72 713.802
R190 GND GND.t254 713.802
R191 GND GND.t90 713.802
R192 GND GND.t214 713.802
R193 GND GND.t184 713.802
R194 GND GND.t204 713.802
R195 GND.n75 GND 713.802
R196 GND.n688 GND.n687 708.047
R197 GND.t58 GND.t323 708.047
R198 GND.t147 GND.t299 708.047
R199 GND.t108 GND.t54 708.047
R200 GND.n694 GND.n693 708.047
R201 GND.n690 GND.n61 708.047
R202 GND.t77 GND.t195 708.047
R203 GND.t2 GND.t77 708.047
R204 GND.t102 GND.t286 708.047
R205 GND.n692 GND.n59 708.047
R206 GND.t306 GND.t76 674.331
R207 GND.t41 GND.t303 674.331
R208 GND.n489 GND.n487 668.355
R209 GND.n507 GND.n430 668.355
R210 GND.t7 GND 649.043
R211 GND.t244 GND 649.043
R212 GND.n588 GND 640.614
R213 GND.n580 GND 632.184
R214 GND.n694 GND 623.755
R215 GND GND.n59 623.755
R216 GND.n530 GND.n529 618.521
R217 GND.n695 GND.n694 599.125
R218 GND.n634 GND.n61 599.125
R219 GND.n594 GND.n59 599.125
R220 GND GND.t6 590.654
R221 GND.t242 GND 590.038
R222 GND.t16 GND 590.038
R223 GND.t290 GND 590.038
R224 GND GND.t153 590.038
R225 GND GND.t70 590.038
R226 GND GND.t139 590.038
R227 GND.n112 GND.n108 585
R228 GND.n114 GND.n113 585
R229 GND.n113 GND.n106 585
R230 GND.n121 GND.n120 585
R231 GND.n122 GND.n121 585
R232 GND.n105 GND.n104 585
R233 GND.n123 GND.n105 585
R234 GND.n130 GND.n129 585
R235 GND.n129 GND.n128 585
R236 GND.n126 GND.n125 585
R237 GND.n127 GND.n126 585
R238 GND.n101 GND.n100 585
R239 GND.n124 GND.n100 585
R240 GND.n143 GND.n142 585
R241 GND.n144 GND.n143 585
R242 GND.n136 GND.n99 585
R243 GND.n145 GND.n99 585
R244 GND.n147 GND.n98 585
R245 GND.n147 GND.n146 585
R246 GND.n149 GND.n148 585
R247 GND.n148 GND.n94 585
R248 GND.n417 GND.n416 585
R249 GND.n418 GND.n417 585
R250 GND.n96 GND.n95 585
R251 GND.n158 GND.n95 585
R252 GND.n156 GND.n154 585
R253 GND.n159 GND.n156 585
R254 GND.n409 GND.n408 585
R255 GND.n408 GND.n407 585
R256 GND.n157 GND.n155 585
R257 GND.n406 GND.n157 585
R258 GND.n404 GND.n403 585
R259 GND.n405 GND.n404 585
R260 GND.n398 GND.n163 585
R261 GND.n163 GND.n160 585
R262 GND.n397 GND.n396 585
R263 GND.n396 GND.n395 585
R264 GND.n165 GND.n164 585
R265 GND.n394 GND.n165 585
R266 GND.n392 GND.n391 585
R267 GND.n393 GND.n392 585
R268 GND.n390 GND.n166 585
R269 GND.n174 GND.n166 585
R270 GND.n389 GND.n388 585
R271 GND.n388 GND.n387 585
R272 GND.n385 GND.n384 585
R273 GND.n386 GND.n385 585
R274 GND.n176 GND.n175 585
R275 GND.n186 GND.n175 585
R276 GND.n184 GND.n182 585
R277 GND.n187 GND.n184 585
R278 GND.n377 GND.n376 585
R279 GND.n376 GND.n375 585
R280 GND.n185 GND.n183 585
R281 GND.n374 GND.n185 585
R282 GND.n372 GND.n371 585
R283 GND.n373 GND.n372 585
R284 GND.n366 GND.n191 585
R285 GND.n191 GND.n188 585
R286 GND.n365 GND.n364 585
R287 GND.n364 GND.n363 585
R288 GND.n193 GND.n192 585
R289 GND.n362 GND.n193 585
R290 GND.n360 GND.n359 585
R291 GND.n361 GND.n360 585
R292 GND.n358 GND.n194 585
R293 GND.n202 GND.n194 585
R294 GND.n357 GND.n356 585
R295 GND.n356 GND.n355 585
R296 GND.n353 GND.n352 585
R297 GND.n354 GND.n353 585
R298 GND.n204 GND.n203 585
R299 GND.n214 GND.n203 585
R300 GND.n212 GND.n210 585
R301 GND.n215 GND.n212 585
R302 GND.n345 GND.n344 585
R303 GND.n344 GND.n343 585
R304 GND.n213 GND.n211 585
R305 GND.n342 GND.n213 585
R306 GND.n340 GND.n339 585
R307 GND.n341 GND.n340 585
R308 GND.n334 GND.n219 585
R309 GND.n219 GND.n216 585
R310 GND.n333 GND.n332 585
R311 GND.n332 GND.n331 585
R312 GND.n221 GND.n220 585
R313 GND.n330 GND.n221 585
R314 GND.n328 GND.n327 585
R315 GND.n329 GND.n328 585
R316 GND.n326 GND.n222 585
R317 GND.n230 GND.n222 585
R318 GND.n325 GND.n324 585
R319 GND.n324 GND.n323 585
R320 GND.n321 GND.n320 585
R321 GND.n322 GND.n321 585
R322 GND.n232 GND.n231 585
R323 GND.n242 GND.n231 585
R324 GND.n240 GND.n238 585
R325 GND.n243 GND.n240 585
R326 GND.n313 GND.n312 585
R327 GND.n312 GND.n311 585
R328 GND.n241 GND.n239 585
R329 GND.n310 GND.n241 585
R330 GND.n308 GND.n307 585
R331 GND.n309 GND.n308 585
R332 GND.n302 GND.n247 585
R333 GND.n247 GND.n244 585
R334 GND.n301 GND.n300 585
R335 GND.n300 GND.n299 585
R336 GND.n249 GND.n248 585
R337 GND.n298 GND.n249 585
R338 GND.n296 GND.n295 585
R339 GND.n297 GND.n296 585
R340 GND.n251 GND.n250 585
R341 GND.n261 GND.n250 585
R342 GND.n263 GND.n262 585
R343 GND.n264 GND.n263 585
R344 GND.n288 GND.n258 585
R345 GND.n265 GND.n258 585
R346 GND.n287 GND.n286 585
R347 GND.n286 GND.n285 585
R348 GND.n260 GND.n259 585
R349 GND.n284 GND.n260 585
R350 GND.n282 GND.n281 585
R351 GND.n283 GND.n282 585
R352 GND.n268 GND.n267 585
R353 GND.n267 GND.n266 585
R354 GND.n274 GND.n273 585
R355 GND.n273 GND.n60 585
R356 GND GND.t208 539.465
R357 GND GND.t165 539.465
R358 GND GND.t168 539.465
R359 GND GND.t2 539.465
R360 GND.t206 GND 539.465
R361 GND.n282 GND.n267 539.294
R362 GND.n273 GND.n267 539.294
R363 GND.n286 GND.n258 539.294
R364 GND.n286 GND.n260 539.294
R365 GND.n296 GND.n250 539.294
R366 GND.n263 GND.n250 539.294
R367 GND.n300 GND.n247 539.294
R368 GND.n300 GND.n249 539.294
R369 GND.n321 GND.n231 539.294
R370 GND.n240 GND.n231 539.294
R371 GND.n312 GND.n240 539.294
R372 GND.n312 GND.n241 539.294
R373 GND.n308 GND.n241 539.294
R374 GND.n332 GND.n219 539.294
R375 GND.n332 GND.n221 539.294
R376 GND.n328 GND.n221 539.294
R377 GND.n328 GND.n222 539.294
R378 GND.n324 GND.n222 539.294
R379 GND.n353 GND.n203 539.294
R380 GND.n212 GND.n203 539.294
R381 GND.n344 GND.n212 539.294
R382 GND.n344 GND.n213 539.294
R383 GND.n340 GND.n213 539.294
R384 GND.n364 GND.n191 539.294
R385 GND.n364 GND.n193 539.294
R386 GND.n360 GND.n193 539.294
R387 GND.n360 GND.n194 539.294
R388 GND.n356 GND.n194 539.294
R389 GND.n385 GND.n175 539.294
R390 GND.n184 GND.n175 539.294
R391 GND.n376 GND.n184 539.294
R392 GND.n376 GND.n185 539.294
R393 GND.n372 GND.n185 539.294
R394 GND.n396 GND.n163 539.294
R395 GND.n396 GND.n165 539.294
R396 GND.n392 GND.n165 539.294
R397 GND.n392 GND.n166 539.294
R398 GND.n388 GND.n166 539.294
R399 GND.n417 GND.n95 539.294
R400 GND.n156 GND.n95 539.294
R401 GND.n408 GND.n156 539.294
R402 GND.n408 GND.n157 539.294
R403 GND.n404 GND.n157 539.294
R404 GND.n147 GND.n99 539.294
R405 GND.n148 GND.n147 539.294
R406 GND.n126 GND.n100 539.294
R407 GND.n143 GND.n100 539.294
R408 GND.n121 GND.n105 539.294
R409 GND.n129 GND.n105 539.294
R410 GND.n113 GND.n112 539.294
R411 GND.n502 GND.n432 525.178
R412 GND.n504 GND.n503 525.178
R413 GND.t186 GND 522.606
R414 GND.t198 GND 522.606
R415 GND GND.t19 514.177
R416 GND.t276 GND.t97 480.461
R417 GND GND.t42 472.031
R418 GND.t99 GND.t187 470.267
R419 GND.t149 GND.t159 470.267
R420 GND.t162 GND.t237 470.267
R421 GND.t332 GND.t148 470.267
R422 GND.t14 GND.t161 470.267
R423 GND.t101 GND.t331 470.267
R424 GND.t160 GND.t13 470.267
R425 GND.t226 GND 455.173
R426 GND.t18 GND.t244 446.743
R427 GND GND.t18 446.743
R428 GND.t301 GND.n645 438.315
R429 GND.n111 GND.t199 416.084
R430 GND GND.t276 413.027
R431 GND.t336 GND.n580 404.599
R432 GND.n588 GND.t102 404.599
R433 GND.t330 GND.t235 389.087
R434 GND.t189 GND.t100 389.087
R435 GND.t15 GND.t150 389.087
R436 GND.t19 GND.t7 379.31
R437 GND.t208 GND.n641 370.882
R438 GND.n663 GND.t285 370.882
R439 GND.t48 GND.n662 370.882
R440 GND.n586 GND.t336 370.882
R441 GND.n587 GND.t316 370.882
R442 GND.t0 GND.t131 362.452
R443 GND.t195 GND 362.452
R444 GND GND.t130 357.628
R445 GND GND.t45 357.628
R446 GND GND.t170 357.628
R447 GND GND.t306 354.024
R448 GND.t168 GND.t0 345.594
R449 GND.n641 GND.t194 337.166
R450 GND.n663 GND.t242 337.166
R451 GND.n662 GND.t16 337.166
R452 GND.t153 GND.n586 337.166
R453 GND.t139 GND.n587 337.166
R454 GND.t182 GND.t99 328.938
R455 GND.t264 GND.t149 328.938
R456 GND.t159 GND.t93 328.938
R457 GND.t66 GND.t162 328.938
R458 GND.t237 GND.t46 328.938
R459 GND.t337 GND.t332 328.938
R460 GND.t148 GND.t252 328.938
R461 GND.t277 GND.t14 328.938
R462 GND.t161 GND.t196 328.938
R463 GND.t143 GND.t101 328.938
R464 GND.t331 GND.t171 328.938
R465 GND.t74 GND.t160 328.938
R466 GND.t97 GND.t86 328.736
R467 GND.t194 GND 295.019
R468 GND.n713 GND.t174 274.812
R469 GND.n724 GND.t156 274.812
R470 GND.n643 GND.t166 274.812
R471 GND.n668 GND.t59 274.812
R472 GND.t233 GND.t330 272.154
R473 GND.t235 GND.t341 272.154
R474 GND.t288 GND.t189 272.154
R475 GND.t100 GND.t274 272.154
R476 GND.t188 GND.t227 272.154
R477 GND.t256 GND.t236 272.154
R478 GND.t68 GND.t15 272.154
R479 GND.t150 GND.t106 272.154
R480 GND.t30 GND 269.733
R481 GND.t285 GND 269.733
R482 GND.n159 GND.n158 262.197
R483 GND.n407 GND.n159 262.197
R484 GND.n406 GND.n405 262.197
R485 GND.n395 GND.n394 262.197
R486 GND.n394 GND.n393 262.197
R487 GND.n387 GND.n174 262.197
R488 GND.n187 GND.n186 262.197
R489 GND.n375 GND.n187 262.197
R490 GND.n374 GND.n373 262.197
R491 GND.n363 GND.n362 262.197
R492 GND.n362 GND.n361 262.197
R493 GND.n355 GND.n202 262.197
R494 GND.n215 GND.n214 262.197
R495 GND.n343 GND.n215 262.197
R496 GND.n342 GND.n341 262.197
R497 GND.n331 GND.n330 262.197
R498 GND.n330 GND.n329 262.197
R499 GND.n323 GND.n230 262.197
R500 GND.n243 GND.n242 262.197
R501 GND.n311 GND.n243 262.197
R502 GND.n310 GND.n309 262.197
R503 GND.n299 GND.n298 262.197
R504 GND.n264 GND.n261 262.197
R505 GND.n285 GND.n284 262.197
R506 GND.n266 GND.n60 262.197
R507 GND GND.t48 252.875
R508 GND GND.t147 252.875
R509 GND GND.t108 252.875
R510 GND.t316 GND 252.875
R511 GND GND.t28 249.387
R512 GND.t298 GND.t60 246.237
R513 GND.t80 GND.t219 246.237
R514 GND.t249 GND.t62 246.237
R515 GND.n418 GND.t345 243.079
R516 GND.n407 GND.t22 243.079
R517 GND.t328 GND.n160 243.079
R518 GND.n393 GND.t238 243.079
R519 GND.n386 GND.t11 243.079
R520 GND.n375 GND.t133 243.079
R521 GND.t202 GND.n188 243.079
R522 GND.n361 GND.t260 243.079
R523 GND.n354 GND.t180 243.079
R524 GND.n343 GND.t283 243.079
R525 GND.t212 GND.n216 243.079
R526 GND.n329 GND.t141 243.079
R527 GND.n322 GND.t240 243.079
R528 GND.n311 GND.t246 243.079
R529 GND.t334 GND.n244 243.079
R530 GND.n297 GND.t216 243.079
R531 GND.t20 GND.n265 243.079
R532 GND.n283 GND.t24 243.079
R533 GND.t165 GND 236.016
R534 GND.n75 GND.t192 234.901
R535 GND.t112 GND.t35 234.511
R536 GND.t111 GND.t175 234.511
R537 GND.t113 GND.t270 234.511
R538 GND.t63 GND.t297 222.786
R539 GND.t65 GND.t103 222.786
R540 GND.t259 GND.t248 222.786
R541 GND.t35 GND 205.197
R542 GND.t60 GND 205.197
R543 GND.t37 GND 205.197
R544 GND.t175 GND 205.197
R545 GND.t219 GND 205.197
R546 GND.t4 GND 205.197
R547 GND.t270 GND 205.197
R548 GND.t62 GND 205.197
R549 GND.t266 GND 205.197
R550 GND.t187 GND.n5 205.118
R551 GND.t201 GND.n52 204.177
R552 GND.n574 GND.n573 196.319
R553 GND.t70 GND 193.87
R554 GND GND.t114 187.608
R555 GND.n487 GND.t61 187.608
R556 GND.n489 GND.t65 187.608
R557 GND GND.t231 187.608
R558 GND.t64 GND.n430 187.608
R559 GND.n507 GND.t259 187.608
R560 GND GND.t281 187.608
R561 GND.n529 GND.t258 187.608
R562 GND GND.t290 185.441
R563 GND GND.t301 185.441
R564 GND.n462 GND.t298 184.678
R565 GND.n488 GND.t80 184.678
R566 GND.n506 GND.t249 184.678
R567 GND.t56 GND.t26 181.745
R568 GND.t324 GND.t135 181.745
R569 GND.t9 GND.t279 181.745
R570 GND GND.t218 179.383
R571 GND.t53 GND 177.925
R572 GND GND.n462 172.952
R573 GND GND.n488 172.952
R574 GND GND.n506 172.952
R575 GND.t297 GND.t262 170.02
R576 GND.t114 GND.t221 170.02
R577 GND.t103 GND.t210 170.02
R578 GND.t231 GND.t177 170.02
R579 GND.t248 GND.t81 170.02
R580 GND.t281 GND.t296 170.02
R581 GND.n753 GND.t44 162.471
R582 GND.n35 GND.t158 162.471
R583 GND.n764 GND.t32 162.471
R584 GND.n31 GND.t230 162.471
R585 GND.n775 GND.t320 162.471
R586 GND.n27 GND.t117 162.471
R587 GND.n786 GND.t225 162.471
R588 GND.n23 GND.t344 162.471
R589 GND.n797 GND.t129 162.471
R590 GND.n19 GND.t269 162.471
R591 GND.n808 GND.t121 162.471
R592 GND.n15 GND.t89 162.471
R593 GND.n819 GND.t251 162.471
R594 GND.n11 GND.t340 162.471
R595 GND.n830 GND.t84 162.471
R596 GND.n6 GND.t119 162.471
R597 GND.n845 GND.t127 162.471
R598 GND.n3 GND.t146 162.471
R599 GND.n39 GND.t315 162.471
R600 GND.n742 GND.t191 162.471
R601 GND.n749 GND.t215 160.017
R602 GND.n754 GND.t91 160.017
R603 GND.n760 GND.t255 160.017
R604 GND.n765 GND.t73 160.017
R605 GND.n771 GND.t96 160.017
R606 GND.n776 GND.t138 160.017
R607 GND.n782 GND.t52 160.017
R608 GND.n787 GND.t322 160.017
R609 GND.n793 GND.t318 160.017
R610 GND.n798 GND.t273 160.017
R611 GND.n804 GND.t152 160.017
R612 GND.n809 GND.t179 160.017
R613 GND.n815 GND.t34 160.017
R614 GND.n820 GND.t223 160.017
R615 GND.n826 GND.t50 160.017
R616 GND.n831 GND.t308 160.017
R617 GND.n7 GND.t123 160.017
R618 GND.n844 GND.t110 160.017
R619 GND.n743 GND.t185 160.017
R620 GND.n43 GND.t205 160.017
R621 GND.n48 GND.t29 158.361
R622 GND.n639 GND.t98 158.361
R623 GND.n681 GND.t125 158.361
R624 GND.n583 GND.t245 158.361
R625 GND.n581 GND.t8 158.361
R626 GND.t104 GND.t37 158.294
R627 GND.t312 GND.t4 158.294
R628 GND.t310 GND.t266 158.294
R629 GND.n605 GND.t3 155.63
R630 GND.t28 GND 154.591
R631 GND.n609 GND.t85 154.131
R632 GND.n633 GND.t132 154.131
R633 GND.n109 GND.t200 153.707
R634 GND.n578 GND.t1 153.631
R635 GND.n537 GND.n93 153.276
R636 GND.n628 GND.t169 152.381
R637 GND.n645 GND 151.725
R638 GND.n539 GND.n538 151.319
R639 GND.n540 GND.n539 151.319
R640 GND.n572 GND.n571 151.319
R641 GND.n573 GND.n572 151.319
R642 GND.n570 GND.n66 151.319
R643 GND.n571 GND.n570 151.319
R644 GND.n72 GND.n71 151.319
R645 GND.n71 GND.n66 151.319
R646 GND.n556 GND.n555 151.319
R647 GND.n556 GND.n72 151.319
R648 GND.n554 GND.n553 151.319
R649 GND.n555 GND.n554 151.319
R650 GND.n552 GND.n80 151.319
R651 GND.n553 GND.n552 151.319
R652 GND.n86 GND.n85 151.319
R653 GND.n85 GND.n80 151.319
R654 GND.n541 GND.n540 151.319
R655 GND.n541 GND.n86 151.319
R656 GND.n538 GND.n537 151.319
R657 GND.n452 GND.t38 150.922
R658 GND.n455 GND.t309 150.922
R659 GND.n445 GND.t220 150.922
R660 GND.n439 GND.t5 150.922
R661 GND.n521 GND.t87 150.922
R662 GND.n527 GND.t267 150.922
R663 GND.n513 GND.t10 150.922
R664 GND.n518 GND.t271 150.922
R665 GND.n496 GND.t325 150.922
R666 GND.n498 GND.t176 150.922
R667 GND.n707 GND.t164 150.922
R668 GND.n702 GND.t327 150.922
R669 GND.n651 GND.t55 150.922
R670 GND.n655 GND.t291 150.922
R671 GND.n656 GND.t300 150.922
R672 GND.n646 GND.t17 150.922
R673 GND.n644 GND.t243 150.922
R674 GND.n58 GND.t302 150.922
R675 GND.n614 GND.t140 150.922
R676 GND.n618 GND.t71 150.922
R677 GND.n623 GND.t154 150.922
R678 GND.n600 GND.t287 150.922
R679 GND.n470 GND.t57 150.922
R680 GND.n475 GND.t36 150.922
R681 GND.n605 GND.t305 149.493
R682 GND.n640 GND.t209 149.493
R683 GND.n139 GND.t40 149.067
R684 GND.n133 GND.t79 149.067
R685 GND.n117 GND.t293 149.067
R686 GND.n277 GND.t25 149.067
R687 GND.n271 GND.t21 149.067
R688 GND.n291 GND.t217 149.067
R689 GND.n254 GND.t335 149.067
R690 GND.n304 GND.t247 149.067
R691 GND.n316 GND.t241 149.067
R692 GND.n234 GND.t142 149.067
R693 GND.n225 GND.t213 149.067
R694 GND.n336 GND.t284 149.067
R695 GND.n348 GND.t181 149.067
R696 GND.n206 GND.t261 149.067
R697 GND.n197 GND.t203 149.067
R698 GND.n368 GND.t134 149.067
R699 GND.n380 GND.t12 149.067
R700 GND.n178 GND.t239 149.067
R701 GND.n169 GND.t329 149.067
R702 GND.n400 GND.t23 149.067
R703 GND.n412 GND.t346 149.067
R704 GND.n591 GND.t304 147.411
R705 GND.n590 GND.t207 146.245
R706 GND.t6 GND.t92 140.007
R707 GND.t218 GND.t333 140.007
R708 GND.n688 GND 138.548
R709 GND.t286 GND.t226 134.867
R710 GND.n57 GND.n55 134.173
R711 GND.t92 GND.t155 122.507
R712 GND.t333 GND.t173 122.507
R713 GND.t163 GND.t201 122.507
R714 GND.t326 GND.t53 122.507
R715 GND.n112 GND.n111 116.203
R716 GND GND.n52 110.84
R717 GND.n55 GND 107.922
R718 GND.t294 GND.n5 102.447
R719 GND GND.t163 102.088
R720 GND GND.t326 102.088
R721 GND.t155 GND 93.3383
R722 GND.t173 GND 93.3383
R723 GND.t221 GND.t104 87.9419
R724 GND.t177 GND.t312 87.9419
R725 GND.t296 GND.t310 87.9419
R726 GND.t262 GND.t56 76.2164
R727 GND.t210 GND.t324 76.2164
R728 GND.t81 GND.t9 76.2164
R729 GND.t292 GND.n123 73.3338
R730 GND.n124 GND.t78 73.3338
R731 GND.n146 GND.t39 73.3338
R732 GND.t42 GND.t58 67.4335
R733 GND.t299 GND.t186 67.4335
R734 GND.t54 GND.t198 67.4335
R735 GND.n543 GND.t182 55.0318
R736 GND.n543 GND.t264 55.0318
R737 GND.t93 GND.n89 55.0318
R738 GND.n89 GND.t66 55.0318
R739 GND.n550 GND.t46 55.0318
R740 GND.n550 GND.t337 55.0318
R741 GND.t252 GND.n549 55.0318
R742 GND.n549 GND.t277 55.0318
R743 GND.n558 GND.t196 55.0318
R744 GND.n558 GND.t143 55.0318
R745 GND.t171 GND.n76 55.0318
R746 GND.n76 GND.t74 55.0318
R747 GND.n65 GND.n62 45.7159
R748 GND.n566 GND.n565 45.7159
R749 GND.n563 GND.n562 45.7159
R750 GND.n561 GND.n68 45.7159
R751 GND.n560 GND.n559 45.7159
R752 GND.n79 GND.n74 45.7159
R753 GND.n548 GND.n547 45.7159
R754 GND.n546 GND.n82 45.7159
R755 GND.n545 GND.n544 45.7159
R756 GND.n92 GND.n88 45.7159
R757 GND.n533 GND.n532 45.7159
R758 GND.n568 GND.t192 45.532
R759 GND.n568 GND.t233 45.532
R760 GND.t341 GND.n567 45.532
R761 GND.n567 GND.t288 45.532
R762 GND.n575 GND.t274 45.532
R763 GND.t227 GND.n575 45.532
R764 GND.n535 GND.t256 45.532
R765 GND.n535 GND.t68 45.532
R766 GND.t106 GND.n534 45.532
R767 GND.n534 GND.t294 45.532
R768 GND.n575 GND.n62 45.0005
R769 GND.n567 GND.n566 45.0005
R770 GND.n568 GND.n563 45.0005
R771 GND.n76 GND.n68 45.0005
R772 GND.n559 GND.n558 45.0005
R773 GND.n549 GND.n74 45.0005
R774 GND.n550 GND.n548 45.0005
R775 GND.n89 GND.n82 45.0005
R776 GND.n544 GND.n543 45.0005
R777 GND.n534 GND.n88 45.0005
R778 GND.n535 GND.n533 45.0005
R779 GND.n539 GND.n90 45.0005
R780 GND.n534 GND.n90 45.0005
R781 GND.n575 GND.n574 45.0005
R782 GND.n572 GND.n63 45.0005
R783 GND.n567 GND.n63 45.0005
R784 GND.n570 GND.n569 45.0005
R785 GND.n569 GND.n568 45.0005
R786 GND.n71 GND.n67 45.0005
R787 GND.n76 GND.n67 45.0005
R788 GND.n557 GND.n556 45.0005
R789 GND.n558 GND.n557 45.0005
R790 GND.n554 GND.n77 45.0005
R791 GND.n549 GND.n77 45.0005
R792 GND.n552 GND.n551 45.0005
R793 GND.n551 GND.n550 45.0005
R794 GND.n85 GND.n81 45.0005
R795 GND.n89 GND.n81 45.0005
R796 GND.n542 GND.n541 45.0005
R797 GND.n543 GND.n542 45.0005
R798 GND.n537 GND.n536 45.0005
R799 GND.n536 GND.n535 45.0005
R800 GND.n735 GND.n734 43.9358
R801 GND.n505 GND.n504 41.7076
R802 GND.n520 GND.n519 39.8486
R803 GND.n447 GND.n446 39.8486
R804 GND.n477 GND.n476 39.8486
R805 GND.n136 GND.n98 36.1417
R806 GND.n149 GND.n98 36.1417
R807 GND.n125 GND.n101 36.1417
R808 GND.n142 GND.n101 36.1417
R809 GND.n120 GND.n104 36.1417
R810 GND.n130 GND.n104 36.1417
R811 GND.n281 GND.n268 36.1417
R812 GND.n274 GND.n268 36.1417
R813 GND.n288 GND.n287 36.1417
R814 GND.n287 GND.n259 36.1417
R815 GND.n295 GND.n251 36.1417
R816 GND.n262 GND.n251 36.1417
R817 GND.n302 GND.n301 36.1417
R818 GND.n301 GND.n248 36.1417
R819 GND.n320 GND.n232 36.1417
R820 GND.n238 GND.n232 36.1417
R821 GND.n313 GND.n238 36.1417
R822 GND.n313 GND.n239 36.1417
R823 GND.n307 GND.n239 36.1417
R824 GND.n334 GND.n333 36.1417
R825 GND.n333 GND.n220 36.1417
R826 GND.n327 GND.n220 36.1417
R827 GND.n327 GND.n326 36.1417
R828 GND.n326 GND.n325 36.1417
R829 GND.n352 GND.n204 36.1417
R830 GND.n210 GND.n204 36.1417
R831 GND.n345 GND.n210 36.1417
R832 GND.n345 GND.n211 36.1417
R833 GND.n339 GND.n211 36.1417
R834 GND.n366 GND.n365 36.1417
R835 GND.n365 GND.n192 36.1417
R836 GND.n359 GND.n192 36.1417
R837 GND.n359 GND.n358 36.1417
R838 GND.n358 GND.n357 36.1417
R839 GND.n384 GND.n176 36.1417
R840 GND.n182 GND.n176 36.1417
R841 GND.n377 GND.n182 36.1417
R842 GND.n377 GND.n183 36.1417
R843 GND.n371 GND.n183 36.1417
R844 GND.n398 GND.n397 36.1417
R845 GND.n397 GND.n164 36.1417
R846 GND.n391 GND.n164 36.1417
R847 GND.n391 GND.n390 36.1417
R848 GND.n390 GND.n389 36.1417
R849 GND.n416 GND.n96 36.1417
R850 GND.n154 GND.n96 36.1417
R851 GND.n409 GND.n154 36.1417
R852 GND.n409 GND.n155 36.1417
R853 GND.n403 GND.n155 36.1417
R854 GND.n110 GND.n108 36.1417
R855 GND.n114 GND.n108 36.1417
R856 GND.n482 GND.n481 34.6358
R857 GND.n440 GND.n434 34.6358
R858 GND.n526 GND.n422 34.6358
R859 GND.n512 GND.n429 34.6358
R860 GND.n517 GND.n426 34.6358
R861 GND.n491 GND.n449 34.6358
R862 GND.n499 GND.n497 34.6358
R863 GND.n719 GND.n718 34.6358
R864 GND.n718 GND.n49 34.6358
R865 GND.n714 GND.n49 34.6358
R866 GND.n723 GND.n47 34.6358
R867 GND.n734 GND.n44 34.6358
R868 GND.n730 GND.n44 34.6358
R869 GND.n730 GND.n729 34.6358
R870 GND.n729 GND.n728 34.6358
R871 GND.n728 GND.n46 34.6358
R872 GND.n708 GND.n51 34.6358
R873 GND.n706 GND.n54 34.6358
R874 GND.n670 GND.n669 34.6358
R875 GND.n680 GND.n679 34.6358
R876 GND.n679 GND.n638 34.6358
R877 GND.n682 GND.n576 34.6358
R878 GND.n599 GND.n589 34.6358
R879 GND.n469 GND.n460 34.6358
R880 GND.n474 GND.n457 34.6358
R881 GND.t323 GND.t167 33.717
R882 GND.t76 GND.t41 33.717
R883 GND.t303 GND.t206 33.717
R884 GND.n524 GND.n423 33.5688
R885 GND.n442 GND.n435 33.5688
R886 GND.n428 GND.n427 33.5688
R887 GND.n454 GND.n453 33.5688
R888 GND.n494 GND.n450 33.5688
R889 GND.n459 GND.n458 33.5688
R890 GND.n590 GND.n589 32.7534
R891 GND.n506 GND.n505 30.79
R892 GND.n503 GND.n431 30.79
R893 GND.n488 GND.n431 30.79
R894 GND.n461 GND.n432 30.79
R895 GND.n462 GND.n461 30.79
R896 GND GND.t61 29.3143
R897 GND GND.t64 29.3143
R898 GND GND.t258 29.3143
R899 GND.n714 GND.n713 25.977
R900 GND.n724 GND.n46 25.977
R901 GND.n669 GND.n668 25.977
R902 GND.n753 GND.n38 25.224
R903 GND.n749 GND.n38 25.224
R904 GND.n755 GND.n35 25.224
R905 GND.n755 GND.n754 25.224
R906 GND.n764 GND.n34 25.224
R907 GND.n760 GND.n34 25.224
R908 GND.n766 GND.n31 25.224
R909 GND.n766 GND.n765 25.224
R910 GND.n775 GND.n30 25.224
R911 GND.n771 GND.n30 25.224
R912 GND.n777 GND.n27 25.224
R913 GND.n777 GND.n776 25.224
R914 GND.n786 GND.n26 25.224
R915 GND.n782 GND.n26 25.224
R916 GND.n788 GND.n23 25.224
R917 GND.n788 GND.n787 25.224
R918 GND.n797 GND.n22 25.224
R919 GND.n793 GND.n22 25.224
R920 GND.n799 GND.n19 25.224
R921 GND.n799 GND.n798 25.224
R922 GND.n808 GND.n18 25.224
R923 GND.n804 GND.n18 25.224
R924 GND.n810 GND.n15 25.224
R925 GND.n810 GND.n809 25.224
R926 GND.n819 GND.n14 25.224
R927 GND.n815 GND.n14 25.224
R928 GND.n821 GND.n11 25.224
R929 GND.n821 GND.n820 25.224
R930 GND.n830 GND.n10 25.224
R931 GND.n826 GND.n10 25.224
R932 GND.n832 GND.n6 25.224
R933 GND.n832 GND.n831 25.224
R934 GND.n845 GND.n1 25.224
R935 GND.n7 GND.n1 25.224
R936 GND.n843 GND.n3 25.224
R937 GND.n844 GND.n843 25.224
R938 GND.n744 GND.n39 25.224
R939 GND.n744 GND.n743 25.224
R940 GND.n742 GND.n741 25.224
R941 GND.n741 GND.n43 25.224
R942 GND.n532 GND.n531 25.1797
R943 GND.n92 GND.n91 25.1797
R944 GND.n545 GND.n87 25.1797
R945 GND.n546 GND.n84 25.1797
R946 GND.n547 GND.n83 25.1797
R947 GND.n79 GND.n78 25.1797
R948 GND.n560 GND.n73 25.1797
R949 GND.n561 GND.n70 25.1797
R950 GND.n562 GND.n69 25.1797
R951 GND.n565 GND.n564 25.1797
R952 GND.n65 GND.n64 25.1797
R953 GND.n438 GND 24.9384
R954 GND GND.n528 24.9384
R955 GND.n508 GND 24.9384
R956 GND.n490 GND 24.9384
R957 GND GND.n486 24.9384
R958 GND.n463 GND 24.9384
R959 GND.n609 GND.n584 24.4711
R960 GND.n610 GND.n609 24.4711
R961 GND.n633 GND.n577 24.4711
R962 GND.n724 GND.n723 24.0946
R963 GND.n670 GND.n640 24.0946
R964 GND.n595 GND.n594 23.7181
R965 GND.n481 GND.n455 23.7181
R966 GND.n445 GND.n434 23.7181
R967 GND.n521 GND.n422 23.7181
R968 GND.n508 GND.n429 23.7181
R969 GND.n513 GND.n426 23.7181
R970 GND.n491 GND.n490 23.7181
R971 GND.n497 GND.n496 23.7181
R972 GND.n712 GND.n51 23.7181
R973 GND.n707 GND.n706 23.7181
R974 GND.n655 GND.n649 23.7181
R975 GND.n657 GND.n646 23.7181
R976 GND.n675 GND.n674 23.7181
R977 GND.n686 GND.n576 23.7181
R978 GND.n614 GND.n613 23.7181
R979 GND.n623 GND.n622 23.7181
R980 GND.n604 GND.n585 23.7181
R981 GND.n600 GND.n599 23.7181
R982 GND.n463 GND.n460 23.7181
R983 GND.n470 GND.n457 23.7181
R984 GND.t26 GND 23.4515
R985 GND.t135 GND 23.4515
R986 GND.t279 GND 23.4515
R987 GND.n628 GND.n627 23.3417
R988 GND.n482 GND.n452 22.2123
R989 GND.n440 GND.n439 22.2123
R990 GND.n527 GND.n526 22.2123
R991 GND.n513 GND.n512 22.2123
R992 GND.n518 GND.n517 22.2123
R993 GND.n521 GND.n520 22.2123
R994 GND.n496 GND.n449 22.2123
R995 GND.n499 GND.n498 22.2123
R996 GND.n446 GND.n445 22.2123
R997 GND.n708 GND.n707 22.2123
R998 GND.n702 GND.n54 22.2123
R999 GND.n651 GND.n649 22.2123
R1000 GND.n657 GND.n656 22.2123
R1001 GND.n619 GND.n618 22.2123
R1002 GND.n600 GND.n585 22.2123
R1003 GND.n470 GND.n469 22.2123
R1004 GND.n475 GND.n474 22.2123
R1005 GND.n477 GND.n455 22.2123
R1006 GND.n456 GND.n432 21.0574
R1007 GND.t13 GND.n75 20.3866
R1008 GND.n754 GND.n753 20.3299
R1009 GND.n765 GND.n764 20.3299
R1010 GND.n776 GND.n775 20.3299
R1011 GND.n787 GND.n786 20.3299
R1012 GND.n798 GND.n797 20.3299
R1013 GND.n809 GND.n808 20.3299
R1014 GND.n820 GND.n819 20.3299
R1015 GND.n831 GND.n830 20.3299
R1016 GND.n845 GND.n844 20.3299
R1017 GND.n743 GND.n742 20.3299
R1018 GND.n605 GND.n584 19.9534
R1019 GND.n578 GND.n577 19.2005
R1020 GND.n158 GND.t345 19.1191
R1021 GND.t22 GND.n406 19.1191
R1022 GND.n395 GND.t328 19.1191
R1023 GND.n174 GND.t238 19.1191
R1024 GND.n186 GND.t11 19.1191
R1025 GND.t133 GND.n374 19.1191
R1026 GND.n363 GND.t202 19.1191
R1027 GND.n202 GND.t260 19.1191
R1028 GND.n214 GND.t180 19.1191
R1029 GND.t283 GND.n342 19.1191
R1030 GND.n331 GND.t212 19.1191
R1031 GND.n230 GND.t141 19.1191
R1032 GND.n242 GND.t240 19.1191
R1033 GND.t246 GND.n310 19.1191
R1034 GND.n299 GND.t334 19.1191
R1035 GND.n261 GND.t216 19.1191
R1036 GND.n285 GND.t20 19.1191
R1037 GND.n266 GND.t24 19.1191
R1038 GND.n759 GND.n35 17.3181
R1039 GND.n770 GND.n31 17.3181
R1040 GND.n781 GND.n27 17.3181
R1041 GND.n792 GND.n23 17.3181
R1042 GND.n803 GND.n19 17.3181
R1043 GND.n814 GND.n15 17.3181
R1044 GND.n825 GND.n11 17.3181
R1045 GND.n836 GND.n6 17.3181
R1046 GND.n839 GND.n3 17.3181
R1047 GND.n748 GND.n39 17.3181
R1048 GND.n749 GND.n748 15.8123
R1049 GND.n760 GND.n759 15.8123
R1050 GND.n771 GND.n770 15.8123
R1051 GND.n782 GND.n781 15.8123
R1052 GND.n793 GND.n792 15.8123
R1053 GND.n804 GND.n803 15.8123
R1054 GND.n815 GND.n814 15.8123
R1055 GND.n826 GND.n825 15.8123
R1056 GND.n836 GND.n7 15.8123
R1057 GND.n466 GND.n465 15.6245
R1058 GND.n668 GND.n643 15.4358
R1059 GND.n629 GND.n578 15.4358
R1060 GND.n634 GND.n633 13.5534
R1061 GND.n713 GND.n712 13.177
R1062 GND.n664 GND.n643 13.177
R1063 GND.n605 GND.n604 13.177
R1064 GND.n465 GND.n464 13.0995
R1065 GND.n486 GND.n452 12.8005
R1066 GND.n439 GND.n438 12.8005
R1067 GND.n528 GND.n527 12.8005
R1068 GND.n702 GND.n701 12.8005
R1069 GND.n701 GND.n700 12.8005
R1070 GND.n661 GND.n644 12.8005
R1071 GND.n695 GND.n58 12.8005
R1072 GND.n618 GND.n582 12.8005
R1073 GND.n627 GND.n579 12.8005
R1074 GND.t130 GND.t112 11.726
R1075 GND.t45 GND.t111 11.726
R1076 GND.t170 GND.t113 11.726
R1077 GND.n651 GND.n58 11.2946
R1078 GND.n656 GND.n655 11.2946
R1079 GND.n661 GND.n646 11.2946
R1080 GND.n664 GND.n644 11.2946
R1081 GND.n614 GND.n582 11.2946
R1082 GND.n623 GND.n579 11.2946
R1083 GND.n503 GND.n502 10.9181
R1084 GND.n48 GND.n47 10.5417
R1085 GND.n639 GND.n638 10.5417
R1086 GND.n682 GND.n681 10.5417
R1087 GND.n613 GND.n583 10.5417
R1088 GND.n622 GND.n581 10.5417
R1089 GND.n504 GND.n425 10.1398
R1090 GND.n502 GND.n501 10.1398
R1091 GND.n110 GND.n109 9.32838
R1092 GND.n466 GND.n463 9.3031
R1093 GND.n523 GND.n422 9.3005
R1094 GND.n526 GND.n525 9.3005
R1095 GND.n527 GND.n421 9.3005
R1096 GND.n528 GND.n420 9.3005
R1097 GND.n522 GND.n521 9.3005
R1098 GND.n520 GND.n424 9.3005
R1099 GND.n443 GND.n434 9.3005
R1100 GND.n441 GND.n440 9.3005
R1101 GND.n439 GND.n436 9.3005
R1102 GND.n438 GND.n437 9.3005
R1103 GND.n509 GND.n508 9.3005
R1104 GND.n510 GND.n429 9.3005
R1105 GND.n512 GND.n511 9.3005
R1106 GND.n514 GND.n513 9.3005
R1107 GND.n515 GND.n426 9.3005
R1108 GND.n517 GND.n516 9.3005
R1109 GND.n445 GND.n444 9.3005
R1110 GND.n446 GND.n433 9.3005
R1111 GND.n479 GND.n455 9.3005
R1112 GND.n481 GND.n480 9.3005
R1113 GND.n483 GND.n482 9.3005
R1114 GND.n484 GND.n452 9.3005
R1115 GND.n490 GND.n451 9.3005
R1116 GND.n492 GND.n491 9.3005
R1117 GND.n493 GND.n449 9.3005
R1118 GND.n496 GND.n495 9.3005
R1119 GND.n497 GND.n448 9.3005
R1120 GND.n500 GND.n499 9.3005
R1121 GND.n486 GND.n485 9.3005
R1122 GND.n412 GND.n411 9.3005
R1123 GND.n413 GND.n412 9.3005
R1124 GND.n401 GND.n400 9.3005
R1125 GND.n400 GND.n161 9.3005
R1126 GND.n170 GND.n169 9.3005
R1127 GND.n169 GND.n168 9.3005
R1128 GND.n179 GND.n178 9.3005
R1129 GND.n178 GND.n177 9.3005
R1130 GND.n380 GND.n379 9.3005
R1131 GND.n381 GND.n380 9.3005
R1132 GND.n369 GND.n368 9.3005
R1133 GND.n368 GND.n189 9.3005
R1134 GND.n198 GND.n197 9.3005
R1135 GND.n197 GND.n196 9.3005
R1136 GND.n207 GND.n206 9.3005
R1137 GND.n206 GND.n205 9.3005
R1138 GND.n348 GND.n347 9.3005
R1139 GND.n349 GND.n348 9.3005
R1140 GND.n337 GND.n336 9.3005
R1141 GND.n336 GND.n217 9.3005
R1142 GND.n226 GND.n225 9.3005
R1143 GND.n225 GND.n224 9.3005
R1144 GND.n235 GND.n234 9.3005
R1145 GND.n234 GND.n233 9.3005
R1146 GND.n316 GND.n315 9.3005
R1147 GND.n317 GND.n316 9.3005
R1148 GND.n305 GND.n304 9.3005
R1149 GND.n304 GND.n245 9.3005
R1150 GND.n255 GND.n254 9.3005
R1151 GND.n254 GND.n253 9.3005
R1152 GND.n291 GND.n290 9.3005
R1153 GND.n292 GND.n291 9.3005
R1154 GND.n272 GND.n271 9.3005
R1155 GND.n271 GND.n270 9.3005
R1156 GND.n277 GND.n276 9.3005
R1157 GND.n278 GND.n277 9.3005
R1158 GND.n416 GND.n415 9.3005
R1159 GND.n414 GND.n96 9.3005
R1160 GND.n154 GND.n152 9.3005
R1161 GND.n410 GND.n409 9.3005
R1162 GND.n155 GND.n153 9.3005
R1163 GND.n403 GND.n402 9.3005
R1164 GND.n399 GND.n398 9.3005
R1165 GND.n397 GND.n162 9.3005
R1166 GND.n167 GND.n164 9.3005
R1167 GND.n391 GND.n171 9.3005
R1168 GND.n390 GND.n172 9.3005
R1169 GND.n389 GND.n173 9.3005
R1170 GND.n384 GND.n383 9.3005
R1171 GND.n382 GND.n176 9.3005
R1172 GND.n182 GND.n180 9.3005
R1173 GND.n378 GND.n377 9.3005
R1174 GND.n183 GND.n181 9.3005
R1175 GND.n371 GND.n370 9.3005
R1176 GND.n367 GND.n366 9.3005
R1177 GND.n365 GND.n190 9.3005
R1178 GND.n195 GND.n192 9.3005
R1179 GND.n359 GND.n199 9.3005
R1180 GND.n358 GND.n200 9.3005
R1181 GND.n357 GND.n201 9.3005
R1182 GND.n352 GND.n351 9.3005
R1183 GND.n350 GND.n204 9.3005
R1184 GND.n210 GND.n208 9.3005
R1185 GND.n346 GND.n345 9.3005
R1186 GND.n211 GND.n209 9.3005
R1187 GND.n339 GND.n338 9.3005
R1188 GND.n335 GND.n334 9.3005
R1189 GND.n333 GND.n218 9.3005
R1190 GND.n223 GND.n220 9.3005
R1191 GND.n327 GND.n227 9.3005
R1192 GND.n326 GND.n228 9.3005
R1193 GND.n325 GND.n229 9.3005
R1194 GND.n320 GND.n319 9.3005
R1195 GND.n318 GND.n232 9.3005
R1196 GND.n238 GND.n236 9.3005
R1197 GND.n314 GND.n313 9.3005
R1198 GND.n239 GND.n237 9.3005
R1199 GND.n307 GND.n306 9.3005
R1200 GND.n303 GND.n302 9.3005
R1201 GND.n301 GND.n246 9.3005
R1202 GND.n252 GND.n248 9.3005
R1203 GND.n295 GND.n294 9.3005
R1204 GND.n293 GND.n251 9.3005
R1205 GND.n262 GND.n256 9.3005
R1206 GND.n289 GND.n288 9.3005
R1207 GND.n287 GND.n257 9.3005
R1208 GND.n269 GND.n259 9.3005
R1209 GND.n281 GND.n280 9.3005
R1210 GND.n279 GND.n268 9.3005
R1211 GND.n275 GND.n274 9.3005
R1212 GND.n594 GND.n593 9.3005
R1213 GND.n635 GND.n634 9.3005
R1214 GND.n633 GND.n632 9.3005
R1215 GND.n631 GND.n577 9.3005
R1216 GND.n630 GND.n629 9.3005
R1217 GND.n627 GND.n626 9.3005
R1218 GND.n625 GND.n579 9.3005
R1219 GND.n624 GND.n623 9.3005
R1220 GND.n622 GND.n621 9.3005
R1221 GND.n620 GND.n619 9.3005
R1222 GND.n618 GND.n617 9.3005
R1223 GND.n616 GND.n582 9.3005
R1224 GND.n615 GND.n614 9.3005
R1225 GND.n613 GND.n612 9.3005
R1226 GND.n611 GND.n610 9.3005
R1227 GND.n609 GND.n608 9.3005
R1228 GND.n607 GND.n584 9.3005
R1229 GND.n606 GND.n605 9.3005
R1230 GND.n604 GND.n603 9.3005
R1231 GND.n602 GND.n585 9.3005
R1232 GND.n601 GND.n600 9.3005
R1233 GND.n599 GND.n598 9.3005
R1234 GND.n597 GND.n589 9.3005
R1235 GND.n596 GND.n595 9.3005
R1236 GND.n696 GND.n695 9.3005
R1237 GND.n686 GND.n685 9.3005
R1238 GND.n684 GND.n576 9.3005
R1239 GND.n683 GND.n682 9.3005
R1240 GND.n680 GND.n637 9.3005
R1241 GND.n679 GND.n678 9.3005
R1242 GND.n677 GND.n638 9.3005
R1243 GND.n676 GND.n675 9.3005
R1244 GND.n674 GND.n673 9.3005
R1245 GND.n672 GND.n640 9.3005
R1246 GND.n671 GND.n670 9.3005
R1247 GND.n669 GND.n642 9.3005
R1248 GND.n668 GND.n667 9.3005
R1249 GND.n666 GND.n643 9.3005
R1250 GND.n665 GND.n664 9.3005
R1251 GND.n647 GND.n644 9.3005
R1252 GND.n661 GND.n660 9.3005
R1253 GND.n659 GND.n646 9.3005
R1254 GND.n658 GND.n657 9.3005
R1255 GND.n656 GND.n648 9.3005
R1256 GND.n655 GND.n654 9.3005
R1257 GND.n653 GND.n649 9.3005
R1258 GND.n652 GND.n651 9.3005
R1259 GND.n650 GND.n58 9.3005
R1260 GND.n700 GND.n699 9.3005
R1261 GND.n734 GND.n733 9.3005
R1262 GND.n732 GND.n44 9.3005
R1263 GND.n731 GND.n730 9.3005
R1264 GND.n729 GND.n45 9.3005
R1265 GND.n728 GND.n727 9.3005
R1266 GND.n726 GND.n46 9.3005
R1267 GND.n725 GND.n724 9.3005
R1268 GND.n723 GND.n722 9.3005
R1269 GND.n721 GND.n47 9.3005
R1270 GND.n720 GND.n719 9.3005
R1271 GND.n718 GND.n717 9.3005
R1272 GND.n716 GND.n49 9.3005
R1273 GND.n715 GND.n714 9.3005
R1274 GND.n713 GND.n50 9.3005
R1275 GND.n710 GND.n51 9.3005
R1276 GND.n709 GND.n708 9.3005
R1277 GND.n707 GND.n53 9.3005
R1278 GND.n706 GND.n705 9.3005
R1279 GND.n704 GND.n54 9.3005
R1280 GND.n703 GND.n702 9.3005
R1281 GND.n701 GND.n56 9.3005
R1282 GND.n712 GND.n711 9.3005
R1283 GND.n118 GND.n117 9.3005
R1284 GND.n117 GND.n116 9.3005
R1285 GND.n134 GND.n133 9.3005
R1286 GND.n133 GND.n132 9.3005
R1287 GND.n139 GND.n138 9.3005
R1288 GND.n140 GND.n139 9.3005
R1289 GND.n120 GND.n119 9.3005
R1290 GND.n104 GND.n103 9.3005
R1291 GND.n131 GND.n130 9.3005
R1292 GND.n125 GND.n102 9.3005
R1293 GND.n135 GND.n101 9.3005
R1294 GND.n142 GND.n141 9.3005
R1295 GND.n137 GND.n136 9.3005
R1296 GND.n98 GND.n97 9.3005
R1297 GND.n150 GND.n149 9.3005
R1298 GND.n108 GND.n107 9.3005
R1299 GND.n115 GND.n114 9.3005
R1300 GND.n478 GND.n477 9.3005
R1301 GND.n467 GND.n460 9.3005
R1302 GND.n469 GND.n468 9.3005
R1303 GND.n471 GND.n470 9.3005
R1304 GND.n472 GND.n457 9.3005
R1305 GND.n474 GND.n473 9.3005
R1306 GND.n739 GND.n43 9.3005
R1307 GND.n840 GND.n839 9.3005
R1308 GND.n841 GND.n3 9.3005
R1309 GND.n843 GND.n842 9.3005
R1310 GND.n844 GND.n2 9.3005
R1311 GND.n846 GND.n845 9.3005
R1312 GND.n1 GND.n0 9.3005
R1313 GND.n8 GND.n7 9.3005
R1314 GND.n836 GND.n835 9.3005
R1315 GND.n834 GND.n6 9.3005
R1316 GND.n833 GND.n832 9.3005
R1317 GND.n831 GND.n9 9.3005
R1318 GND.n830 GND.n829 9.3005
R1319 GND.n828 GND.n10 9.3005
R1320 GND.n827 GND.n826 9.3005
R1321 GND.n825 GND.n824 9.3005
R1322 GND.n823 GND.n11 9.3005
R1323 GND.n822 GND.n821 9.3005
R1324 GND.n820 GND.n13 9.3005
R1325 GND.n819 GND.n818 9.3005
R1326 GND.n817 GND.n14 9.3005
R1327 GND.n816 GND.n815 9.3005
R1328 GND.n814 GND.n813 9.3005
R1329 GND.n812 GND.n15 9.3005
R1330 GND.n811 GND.n810 9.3005
R1331 GND.n809 GND.n17 9.3005
R1332 GND.n808 GND.n807 9.3005
R1333 GND.n806 GND.n18 9.3005
R1334 GND.n805 GND.n804 9.3005
R1335 GND.n803 GND.n802 9.3005
R1336 GND.n801 GND.n19 9.3005
R1337 GND.n800 GND.n799 9.3005
R1338 GND.n798 GND.n21 9.3005
R1339 GND.n797 GND.n796 9.3005
R1340 GND.n795 GND.n22 9.3005
R1341 GND.n794 GND.n793 9.3005
R1342 GND.n792 GND.n791 9.3005
R1343 GND.n790 GND.n23 9.3005
R1344 GND.n789 GND.n788 9.3005
R1345 GND.n787 GND.n25 9.3005
R1346 GND.n786 GND.n785 9.3005
R1347 GND.n784 GND.n26 9.3005
R1348 GND.n783 GND.n782 9.3005
R1349 GND.n781 GND.n780 9.3005
R1350 GND.n779 GND.n27 9.3005
R1351 GND.n778 GND.n777 9.3005
R1352 GND.n776 GND.n29 9.3005
R1353 GND.n775 GND.n774 9.3005
R1354 GND.n773 GND.n30 9.3005
R1355 GND.n772 GND.n771 9.3005
R1356 GND.n770 GND.n769 9.3005
R1357 GND.n768 GND.n31 9.3005
R1358 GND.n767 GND.n766 9.3005
R1359 GND.n765 GND.n33 9.3005
R1360 GND.n764 GND.n763 9.3005
R1361 GND.n762 GND.n34 9.3005
R1362 GND.n761 GND.n760 9.3005
R1363 GND.n759 GND.n758 9.3005
R1364 GND.n757 GND.n35 9.3005
R1365 GND.n756 GND.n755 9.3005
R1366 GND.n754 GND.n37 9.3005
R1367 GND.n753 GND.n752 9.3005
R1368 GND.n751 GND.n38 9.3005
R1369 GND.n750 GND.n749 9.3005
R1370 GND.n748 GND.n747 9.3005
R1371 GND.n746 GND.n39 9.3005
R1372 GND.n745 GND.n744 9.3005
R1373 GND.n743 GND.n41 9.3005
R1374 GND.n742 GND.n42 9.3005
R1375 GND.n741 GND.n740 9.3005
R1376 GND.n674 GND.n640 9.03579
R1377 GND.n423 GND.t282 8.7005
R1378 GND.n423 GND.t311 8.7005
R1379 GND.n435 GND.t232 8.7005
R1380 GND.n435 GND.t313 8.7005
R1381 GND.n427 GND.t82 8.7005
R1382 GND.n427 GND.t280 8.7005
R1383 GND.n453 GND.t115 8.7005
R1384 GND.n453 GND.t105 8.7005
R1385 GND.n450 GND.t211 8.7005
R1386 GND.n450 GND.t136 8.7005
R1387 GND.n458 GND.t263 8.7005
R1388 GND.n458 GND.t27 8.7005
R1389 GND.n719 GND.n48 6.77697
R1390 GND.n675 GND.n639 6.77697
R1391 GND.n681 GND.n680 6.77697
R1392 GND.n610 GND.n583 6.77697
R1393 GND.n619 GND.n581 6.77697
R1394 GND.n531 GND.t257 5.8005
R1395 GND.n531 GND.t69 5.8005
R1396 GND.n91 GND.t107 5.8005
R1397 GND.n91 GND.t295 5.8005
R1398 GND.n87 GND.t183 5.8005
R1399 GND.n87 GND.t265 5.8005
R1400 GND.n84 GND.t94 5.8005
R1401 GND.n84 GND.t67 5.8005
R1402 GND.n83 GND.t47 5.8005
R1403 GND.n83 GND.t338 5.8005
R1404 GND.n78 GND.t253 5.8005
R1405 GND.n78 GND.t278 5.8005
R1406 GND.n73 GND.t197 5.8005
R1407 GND.n73 GND.t144 5.8005
R1408 GND.n70 GND.t172 5.8005
R1409 GND.n70 GND.t75 5.8005
R1410 GND.n69 GND.t193 5.8005
R1411 GND.n69 GND.t234 5.8005
R1412 GND.n564 GND.t342 5.8005
R1413 GND.n564 GND.t289 5.8005
R1414 GND.n64 GND.t275 5.8005
R1415 GND.n64 GND.t228 5.8005
R1416 GND.n519 GND.n518 5.21334
R1417 GND.n498 GND.n447 5.21334
R1418 GND.n476 GND.n475 5.21334
R1419 GND.n698 GND 4.87704
R1420 GND.n738 GND.n737 4.33704
R1421 GND.n636 GND.n635 4.00641
R1422 GND.n93 GND.n4 3.71362
R1423 GND.n685 GND.n636 3.13461
R1424 GND GND.n592 2.85076
R1425 GND.n697 GND 2.85076
R1426 GND GND.n698 2.85076
R1427 GND GND.n738 2.30925
R1428 GND.n737 GND.n736 2.2505
R1429 GND.n519 GND.n425 2.04483
R1430 GND.n501 GND.n447 2.04483
R1431 GND.n476 GND.n456 2.04483
R1432 GND.n573 GND 1.79008
R1433 GND.n571 GND 1.79008
R1434 GND GND.n66 1.79008
R1435 GND GND.n72 1.79008
R1436 GND.n555 GND 1.79008
R1437 GND.n553 GND 1.79008
R1438 GND GND.n80 1.79008
R1439 GND GND.n86 1.79008
R1440 GND.n540 GND 1.79008
R1441 GND.n538 GND 1.79008
R1442 GND.n151 GND 1.72207
R1443 GND.n738 GND 1.52425
R1444 GND.n840 GND.n4 1.208
R1445 GND.n151 GND.n93 1.17175
R1446 GND.n415 GND.n151 1.15253
R1447 GND.n736 GND 1.13527
R1448 GND.n591 GND.n590 1.12991
R1449 GND.n698 GND.n697 0.872295
R1450 GND.n736 GND.n735 0.856945
R1451 GND.n592 GND 0.846654
R1452 GND.n595 GND.n591 0.753441
R1453 GND.n636 GND 0.683994
R1454 GND.n532 GND 0.645031
R1455 GND GND.n92 0.645031
R1456 GND.n92 GND 0.645031
R1457 GND.n545 GND 0.645031
R1458 GND GND.n545 0.645031
R1459 GND.n546 GND 0.645031
R1460 GND GND.n546 0.645031
R1461 GND.n547 GND 0.645031
R1462 GND.n547 GND 0.645031
R1463 GND GND.n79 0.645031
R1464 GND.n79 GND 0.645031
R1465 GND.n560 GND 0.645031
R1466 GND GND.n560 0.645031
R1467 GND.n561 GND 0.645031
R1468 GND GND.n561 0.645031
R1469 GND.n562 GND 0.645031
R1470 GND.n562 GND 0.645031
R1471 GND.n565 GND 0.645031
R1472 GND.n565 GND 0.645031
R1473 GND GND.n65 0.645031
R1474 GND.n294 GND 0.633946
R1475 GND GND.n289 0.633946
R1476 GND.n280 GND 0.633946
R1477 GND.n65 GND 0.608898
R1478 GND GND.n303 0.51148
R1479 GND.n592 GND 0.473256
R1480 GND GND.n399 0.390703
R1481 GND.n383 GND 0.390703
R1482 GND GND.n367 0.390703
R1483 GND.n351 GND 0.390703
R1484 GND GND.n335 0.390703
R1485 GND.n319 GND 0.390703
R1486 GND.n629 GND.n628 0.376971
R1487 GND.n465 GND.n4 0.196125
R1488 GND.n737 GND 0.188801
R1489 GND.n522 GND.n424 0.120292
R1490 GND.n525 GND.n421 0.120292
R1491 GND.n444 GND.n433 0.120292
R1492 GND.n441 GND.n436 0.120292
R1493 GND.n511 GND.n510 0.120292
R1494 GND.n516 GND.n515 0.120292
R1495 GND.n479 GND.n478 0.120292
R1496 GND.n484 GND.n483 0.120292
R1497 GND.n493 GND.n492 0.120292
R1498 GND.n500 GND.n448 0.120292
R1499 GND.n632 GND.n631 0.120292
R1500 GND.n631 GND.n630 0.120292
R1501 GND.n621 GND.n620 0.120292
R1502 GND.n612 GND.n611 0.120292
R1503 GND.n608 GND.n607 0.120292
R1504 GND.n607 GND.n606 0.120292
R1505 GND.n602 GND.n601 0.120292
R1506 GND.n598 GND.n597 0.120292
R1507 GND.n597 GND.n596 0.120292
R1508 GND.n684 GND.n683 0.120292
R1509 GND.n683 GND.n637 0.120292
R1510 GND.n678 GND.n677 0.120292
R1511 GND.n677 GND.n676 0.120292
R1512 GND.n671 GND.n642 0.120292
R1513 GND.n667 GND.n642 0.120292
R1514 GND.n658 GND.n648 0.120292
R1515 GND.n653 GND.n652 0.120292
R1516 GND.n733 GND.n732 0.120292
R1517 GND.n732 GND.n731 0.120292
R1518 GND.n731 GND.n45 0.120292
R1519 GND.n727 GND.n45 0.120292
R1520 GND.n727 GND.n726 0.120292
R1521 GND.n726 GND.n725 0.120292
R1522 GND.n722 GND.n721 0.120292
R1523 GND.n721 GND.n720 0.120292
R1524 GND.n717 GND.n716 0.120292
R1525 GND.n716 GND.n715 0.120292
R1526 GND.n715 GND.n50 0.120292
R1527 GND.n710 GND.n709 0.120292
R1528 GND.n709 GND.n53 0.120292
R1529 GND.n705 GND.n704 0.120292
R1530 GND.n704 GND.n703 0.120292
R1531 GND.n468 GND.n467 0.120292
R1532 GND.n473 GND.n472 0.120292
R1533 GND.n509 GND 0.112479
R1534 GND GND.n451 0.112479
R1535 GND.n516 GND.n425 0.109875
R1536 GND.n501 GND.n500 0.109875
R1537 GND.n473 GND.n456 0.109875
R1538 GND.n733 GND 0.105969
R1539 GND.n425 GND.n424 0.104667
R1540 GND.n501 GND.n433 0.104667
R1541 GND.n478 GND.n456 0.104667
R1542 GND.n116 GND 0.0866486
R1543 GND.n415 GND.n414 0.0815811
R1544 GND.n410 GND.n153 0.0815811
R1545 GND.n399 GND.n162 0.0815811
R1546 GND.n172 GND.n171 0.0815811
R1547 GND.n383 GND.n382 0.0815811
R1548 GND.n378 GND.n181 0.0815811
R1549 GND.n367 GND.n190 0.0815811
R1550 GND.n200 GND.n199 0.0815811
R1551 GND.n351 GND.n350 0.0815811
R1552 GND.n346 GND.n209 0.0815811
R1553 GND.n335 GND.n218 0.0815811
R1554 GND.n228 GND.n227 0.0815811
R1555 GND.n319 GND.n318 0.0815811
R1556 GND.n314 GND.n237 0.0815811
R1557 GND.n303 GND.n246 0.0815811
R1558 GND.n294 GND.n293 0.0815811
R1559 GND.n289 GND.n257 0.0815811
R1560 GND.n280 GND.n279 0.0815811
R1561 GND.n115 GND.n107 0.0815811
R1562 GND.n131 GND.n103 0.0815811
R1563 GND.n141 GND.n135 0.0815811
R1564 GND.n150 GND.n97 0.0815811
R1565 GND.n132 GND 0.0807365
R1566 GND GND.n140 0.0807365
R1567 GND.n525 GND.n524 0.0760208
R1568 GND.n442 GND.n441 0.0760208
R1569 GND.n511 GND.n428 0.0760208
R1570 GND.n483 GND.n454 0.0760208
R1571 GND.n494 GND.n493 0.0760208
R1572 GND.n468 GND.n459 0.0760208
R1573 GND.n523 GND 0.0603958
R1574 GND GND.n443 0.0603958
R1575 GND.n437 GND 0.0603958
R1576 GND.n510 GND 0.0603958
R1577 GND.n515 GND 0.0603958
R1578 GND.n480 GND 0.0603958
R1579 GND.n485 GND 0.0603958
R1580 GND.n492 GND 0.0603958
R1581 GND GND.n448 0.0603958
R1582 GND.n632 GND 0.0603958
R1583 GND.n626 GND 0.0603958
R1584 GND GND.n625 0.0603958
R1585 GND GND.n624 0.0603958
R1586 GND.n621 GND 0.0603958
R1587 GND.n617 GND 0.0603958
R1588 GND GND.n616 0.0603958
R1589 GND GND.n615 0.0603958
R1590 GND.n612 GND 0.0603958
R1591 GND.n608 GND 0.0603958
R1592 GND.n603 GND 0.0603958
R1593 GND GND.n602 0.0603958
R1594 GND.n598 GND 0.0603958
R1595 GND.n593 GND 0.0603958
R1596 GND GND.n684 0.0603958
R1597 GND.n678 GND 0.0603958
R1598 GND.n673 GND 0.0603958
R1599 GND GND.n672 0.0603958
R1600 GND GND.n671 0.0603958
R1601 GND GND.n666 0.0603958
R1602 GND GND.n665 0.0603958
R1603 GND.n647 GND 0.0603958
R1604 GND.n660 GND 0.0603958
R1605 GND GND.n659 0.0603958
R1606 GND GND.n658 0.0603958
R1607 GND.n654 GND 0.0603958
R1608 GND GND.n653 0.0603958
R1609 GND GND.n650 0.0603958
R1610 GND.n696 GND 0.0603958
R1611 GND.n722 GND 0.0603958
R1612 GND.n717 GND 0.0603958
R1613 GND.n711 GND 0.0603958
R1614 GND GND.n710 0.0603958
R1615 GND.n705 GND 0.0603958
R1616 GND.n56 GND 0.0603958
R1617 GND.n699 GND 0.0603958
R1618 GND.n467 GND 0.0603958
R1619 GND.n472 GND 0.0603958
R1620 GND.n842 GND.n841 0.058
R1621 GND.n842 GND.n2 0.058
R1622 GND.n846 GND.n0 0.058
R1623 GND.n8 GND.n0 0.058
R1624 GND.n834 GND.n833 0.058
R1625 GND.n833 GND.n9 0.058
R1626 GND.n829 GND.n828 0.058
R1627 GND.n828 GND.n827 0.058
R1628 GND.n823 GND.n822 0.058
R1629 GND.n822 GND.n13 0.058
R1630 GND.n818 GND.n817 0.058
R1631 GND.n817 GND.n816 0.058
R1632 GND.n812 GND.n811 0.058
R1633 GND.n811 GND.n17 0.058
R1634 GND.n807 GND.n806 0.058
R1635 GND.n806 GND.n805 0.058
R1636 GND.n801 GND.n800 0.058
R1637 GND.n800 GND.n21 0.058
R1638 GND.n796 GND.n795 0.058
R1639 GND.n795 GND.n794 0.058
R1640 GND.n790 GND.n789 0.058
R1641 GND.n789 GND.n25 0.058
R1642 GND.n785 GND.n784 0.058
R1643 GND.n784 GND.n783 0.058
R1644 GND.n779 GND.n778 0.058
R1645 GND.n778 GND.n29 0.058
R1646 GND.n774 GND.n773 0.058
R1647 GND.n773 GND.n772 0.058
R1648 GND.n768 GND.n767 0.058
R1649 GND.n767 GND.n33 0.058
R1650 GND.n763 GND.n762 0.058
R1651 GND.n762 GND.n761 0.058
R1652 GND.n757 GND.n756 0.058
R1653 GND.n756 GND.n37 0.058
R1654 GND.n752 GND.n751 0.058
R1655 GND.n751 GND.n750 0.058
R1656 GND.n746 GND.n745 0.058
R1657 GND.n745 GND.n41 0.058
R1658 GND.n740 GND.n42 0.058
R1659 GND.n740 GND.n739 0.058
R1660 GND.n464 GND 0.0577917
R1661 GND.n413 GND.n152 0.0553986
R1662 GND.n402 GND.n161 0.0553986
R1663 GND.n168 GND.n167 0.0553986
R1664 GND.n177 GND.n173 0.0553986
R1665 GND.n381 GND.n180 0.0553986
R1666 GND.n370 GND.n189 0.0553986
R1667 GND.n196 GND.n195 0.0553986
R1668 GND.n205 GND.n201 0.0553986
R1669 GND.n349 GND.n208 0.0553986
R1670 GND.n338 GND.n217 0.0553986
R1671 GND.n224 GND.n223 0.0553986
R1672 GND.n233 GND.n229 0.0553986
R1673 GND.n317 GND.n236 0.0553986
R1674 GND.n306 GND.n245 0.0553986
R1675 GND.n253 GND.n252 0.0553986
R1676 GND.n292 GND.n256 0.0553986
R1677 GND.n270 GND.n269 0.0553986
R1678 GND.n278 GND.n275 0.0553986
R1679 GND.n119 GND.n118 0.0553986
R1680 GND.n134 GND.n102 0.0553986
R1681 GND.n138 GND.n137 0.0553986
R1682 GND.n109 GND.n107 0.0545423
R1683 GND.n524 GND.n523 0.0447708
R1684 GND.n443 GND.n442 0.0447708
R1685 GND.n514 GND.n428 0.0447708
R1686 GND.n480 GND.n454 0.0447708
R1687 GND.n495 GND.n494 0.0447708
R1688 GND.n471 GND.n459 0.0447708
R1689 GND GND.n410 0.0410405
R1690 GND.n171 GND 0.0410405
R1691 GND GND.n378 0.0410405
R1692 GND.n199 GND 0.0410405
R1693 GND GND.n346 0.0410405
R1694 GND.n227 GND 0.0410405
R1695 GND GND.n314 0.0410405
R1696 GND GND.n115 0.0410405
R1697 GND GND.n131 0.0410405
R1698 GND.n141 GND 0.0410405
R1699 GND GND.n150 0.0410405
R1700 GND.n411 GND 0.0351284
R1701 GND GND.n170 0.0351284
R1702 GND.n379 GND 0.0351284
R1703 GND GND.n198 0.0351284
R1704 GND.n347 GND 0.0351284
R1705 GND GND.n226 0.0351284
R1706 GND.n315 GND 0.0351284
R1707 GND GND.n255 0.0351284
R1708 GND.n290 GND 0.0351284
R1709 GND GND.n272 0.0351284
R1710 GND.n276 GND 0.0351284
R1711 GND.n425 GND 0.0343542
R1712 GND.n501 GND 0.0343542
R1713 GND.n616 GND 0.0343542
R1714 GND.n456 GND 0.0343542
R1715 GND.n635 GND 0.0330521
R1716 GND.n626 GND 0.0330521
R1717 GND.n625 GND 0.0330521
R1718 GND.n603 GND 0.0330521
R1719 GND.n593 GND 0.0330521
R1720 GND.n685 GND 0.0330521
R1721 GND.n673 GND 0.0330521
R1722 GND.n665 GND 0.0330521
R1723 GND.n660 GND 0.0330521
R1724 GND GND.n696 0.0330521
R1725 GND.n711 GND 0.0330521
R1726 GND GND.n56 0.0330521
R1727 GND.n699 GND 0.0330521
R1728 GND.n841 GND 0.02925
R1729 GND GND.n846 0.02925
R1730 GND.n835 GND 0.02925
R1731 GND GND.n834 0.02925
R1732 GND.n829 GND 0.02925
R1733 GND.n824 GND 0.02925
R1734 GND GND.n823 0.02925
R1735 GND.n818 GND 0.02925
R1736 GND.n813 GND 0.02925
R1737 GND GND.n812 0.02925
R1738 GND.n807 GND 0.02925
R1739 GND.n802 GND 0.02925
R1740 GND GND.n801 0.02925
R1741 GND.n796 GND 0.02925
R1742 GND.n791 GND 0.02925
R1743 GND GND.n790 0.02925
R1744 GND.n785 GND 0.02925
R1745 GND.n780 GND 0.02925
R1746 GND GND.n779 0.02925
R1747 GND.n774 GND 0.02925
R1748 GND.n769 GND 0.02925
R1749 GND GND.n768 0.02925
R1750 GND.n763 GND 0.02925
R1751 GND.n758 GND 0.02925
R1752 GND GND.n757 0.02925
R1753 GND.n752 GND 0.02925
R1754 GND.n747 GND 0.02925
R1755 GND GND.n746 0.02925
R1756 GND.n42 GND 0.02925
R1757 GND.n414 GND.n413 0.0266824
R1758 GND.n161 GND.n153 0.0266824
R1759 GND.n168 GND.n162 0.0266824
R1760 GND.n177 GND.n172 0.0266824
R1761 GND.n382 GND.n381 0.0266824
R1762 GND.n189 GND.n181 0.0266824
R1763 GND.n196 GND.n190 0.0266824
R1764 GND.n205 GND.n200 0.0266824
R1765 GND.n350 GND.n349 0.0266824
R1766 GND.n217 GND.n209 0.0266824
R1767 GND.n224 GND.n218 0.0266824
R1768 GND.n233 GND.n228 0.0266824
R1769 GND.n318 GND.n317 0.0266824
R1770 GND.n245 GND.n237 0.0266824
R1771 GND.n253 GND.n246 0.0266824
R1772 GND.n293 GND.n292 0.0266824
R1773 GND.n270 GND.n257 0.0266824
R1774 GND.n279 GND.n278 0.0266824
R1775 GND.n118 GND.n103 0.0266824
R1776 GND.n135 GND.n134 0.0266824
R1777 GND.n138 GND.n97 0.0266824
R1778 GND.n697 GND 0.026141
R1779 GND.n401 GND 0.0249932
R1780 GND GND.n179 0.0249932
R1781 GND.n369 GND 0.0249932
R1782 GND GND.n207 0.0249932
R1783 GND.n337 GND 0.0249932
R1784 GND GND.n235 0.0249932
R1785 GND.n305 GND 0.0249932
R1786 GND GND.n522 0.0239375
R1787 GND GND.n421 0.0239375
R1788 GND.n420 GND 0.0239375
R1789 GND.n444 GND 0.0239375
R1790 GND GND.n436 0.0239375
R1791 GND.n437 GND 0.0239375
R1792 GND GND.n509 0.0239375
R1793 GND GND.n514 0.0239375
R1794 GND GND.n479 0.0239375
R1795 GND GND.n484 0.0239375
R1796 GND.n485 GND 0.0239375
R1797 GND.n451 GND 0.0239375
R1798 GND.n495 GND 0.0239375
R1799 GND.n624 GND 0.0239375
R1800 GND.n617 GND 0.0239375
R1801 GND.n615 GND 0.0239375
R1802 GND.n601 GND 0.0239375
R1803 GND GND.n647 0.0239375
R1804 GND.n659 GND 0.0239375
R1805 GND GND.n648 0.0239375
R1806 GND.n654 GND 0.0239375
R1807 GND.n652 GND 0.0239375
R1808 GND.n650 GND 0.0239375
R1809 GND GND.n53 0.0239375
R1810 GND.n703 GND 0.0239375
R1811 GND GND.n471 0.0239375
R1812 GND.n620 GND 0.0226354
R1813 GND.n611 GND 0.0226354
R1814 GND.n676 GND 0.0226354
R1815 GND.n720 GND 0.0226354
R1816 GND.n630 GND 0.0213333
R1817 GND.n606 GND 0.0213333
R1818 GND.n596 GND 0.0213333
R1819 GND.n672 GND 0.0213333
R1820 GND.n667 GND 0.0213333
R1821 GND.n666 GND 0.0213333
R1822 GND.n725 GND 0.0213333
R1823 GND GND.n50 0.0213333
R1824 GND GND.n466 0.0213333
R1825 GND.n425 GND 0.0194732
R1826 GND.n501 GND 0.0194732
R1827 GND.n456 GND 0.0194732
R1828 GND GND.n637 0.016125
R1829 GND GND.n840 0.016125
R1830 GND.n835 GND 0.016125
R1831 GND.n824 GND 0.016125
R1832 GND.n813 GND 0.016125
R1833 GND.n802 GND 0.016125
R1834 GND.n791 GND 0.016125
R1835 GND.n780 GND 0.016125
R1836 GND.n769 GND 0.016125
R1837 GND.n758 GND 0.016125
R1838 GND.n747 GND 0.016125
R1839 GND.n735 GND 0.0148229
R1840 GND.n2 GND 0.011125
R1841 GND GND.n8 0.011125
R1842 GND GND.n9 0.011125
R1843 GND.n827 GND 0.011125
R1844 GND GND.n13 0.011125
R1845 GND.n816 GND 0.011125
R1846 GND GND.n17 0.011125
R1847 GND.n805 GND 0.011125
R1848 GND GND.n21 0.011125
R1849 GND.n794 GND 0.011125
R1850 GND GND.n25 0.011125
R1851 GND.n783 GND 0.011125
R1852 GND GND.n29 0.011125
R1853 GND.n772 GND 0.011125
R1854 GND GND.n33 0.011125
R1855 GND.n761 GND 0.011125
R1856 GND GND.n37 0.011125
R1857 GND.n750 GND 0.011125
R1858 GND GND.n41 0.011125
R1859 GND.n739 GND 0.011125
R1860 GND.n411 GND.n152 0.00641216
R1861 GND.n402 GND.n401 0.00641216
R1862 GND.n170 GND.n167 0.00641216
R1863 GND.n179 GND.n173 0.00641216
R1864 GND.n379 GND.n180 0.00641216
R1865 GND.n370 GND.n369 0.00641216
R1866 GND.n198 GND.n195 0.00641216
R1867 GND.n207 GND.n201 0.00641216
R1868 GND.n347 GND.n208 0.00641216
R1869 GND.n338 GND.n337 0.00641216
R1870 GND.n226 GND.n223 0.00641216
R1871 GND.n235 GND.n229 0.00641216
R1872 GND.n315 GND.n236 0.00641216
R1873 GND.n306 GND.n305 0.00641216
R1874 GND.n255 GND.n252 0.00641216
R1875 GND.n290 GND.n256 0.00641216
R1876 GND.n272 GND.n269 0.00641216
R1877 GND.n276 GND.n275 0.00641216
R1878 GND.n119 GND.n116 0.00641216
R1879 GND.n132 GND.n102 0.00641216
R1880 GND.n140 GND.n137 0.00641216
R1881 GND.n464 GND.n420 0.00310417
R1882 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t5 732.702
R1883 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t4 230.155
R1884 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t8 230.155
R1885 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 208.965
R1886 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t7 157.856
R1887 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t6 157.856
R1888 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 153.72
R1889 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 153.529
R1890 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 96.8352
R1891 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t2 26.5955
R1892 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t3 26.5955
R1893 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 25.1816
R1894 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t0 24.9236
R1895 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t1 24.9236
R1896 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 14.0359
R1897 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 13.0565
R1898 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 11.2645
R1899 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 10.7179
R1900 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 9.3005
R1901 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 7.11508
R1902 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 6.1445
R1903 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 5.23106
R1904 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 4.65505
R1905 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 4.3525
R1906 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 2.86617
R1907 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 2.67513
R1908 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 2.0485
R1909 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 1.55202
R1910 decoder_3_0/decoder_2to4_2.bb[0].n0 decoder_3_0/decoder_2to4_2.bb[0].t1 235.56
R1911 decoder_3_0/decoder_2to4_2.bb[0].n1 decoder_3_0/decoder_2to4_2.bb[0].t4 229.369
R1912 decoder_3_0/decoder_2to4_2.bb[0].n3 decoder_3_0/decoder_2to4_2.bb[0].t5 229.369
R1913 decoder_3_0/decoder_2to4_2.bb[0].n1 decoder_3_0/decoder_2to4_2.bb[0].t2 157.07
R1914 decoder_3_0/decoder_2to4_2.bb[0].n3 decoder_3_0/decoder_2to4_2.bb[0].t3 157.07
R1915 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_2.bb[0].t0 152.889
R1916 decoder_3_0/decoder_2to4_2.bb[0].n2 decoder_3_0/decoder_2to4_2.bb[0].n1 152.712
R1917 decoder_3_0/decoder_2to4_2.bb[0].n4 decoder_3_0/decoder_2to4_2.bb[0].n3 152.475
R1918 decoder_3_0/decoder_2to4_2.bb[0].n7 decoder_3_0/decoder_2to4_2.bb[0] 24.2121
R1919 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_2.bb[0].n6 23.559
R1920 decoder_3_0/decoder_2to4_2.bb[0].n7 decoder_3_0/decoder_2to4_2.bb[0] 14.1918
R1921 decoder_3_0/decoder_2to4_2.bb[0].n5 decoder_3_0/decoder_2to4_2.bb[0].n2 10.2234
R1922 decoder_3_0/decoder_2to4_2.bb[0].n5 decoder_3_0/decoder_2to4_2.bb[0].n4 9.77342
R1923 decoder_3_0/decoder_2to4_2.bb[0].n4 decoder_3_0/decoder_2to4_2.bb[0] 5.45235
R1924 decoder_3_0/decoder_2to4_2.bb[0].n2 decoder_3_0/decoder_2to4_2.bb[0] 5.21532
R1925 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_2.bb[0].n7 4.73093
R1926 decoder_3_0/decoder_2to4_2.bb[0].n6 decoder_3_0/decoder_2to4_2.bb[0].n5 4.6005
R1927 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_2.bb[0].n0 2.22659
R1928 decoder_3_0/decoder_2to4_2.bb[0].n0 decoder_3_0/decoder_2to4_2.bb[0] 1.55202
R1929 decoder_3_0/decoder_2to4_2.bb[0].n6 decoder_3_0/decoder_2to4_2.bb[0] 0.44425
R1930 a_24840_n1428.t0 a_24840_n1428.t1 49.8467
R1931 VBPLV.n2 VBPLV.t6 139.206
R1932 VBPLV.n3 VBPLV.t16 139.206
R1933 VBPLV.n4 VBPLV.t11 139.206
R1934 VBPLV.n5 VBPLV.t20 139.206
R1935 VBPLV.n6 VBPLV.t15 139.206
R1936 VBPLV.n7 VBPLV.t3 139.206
R1937 VBPLV.n8 VBPLV.t19 139.206
R1938 VBPLV.n9 VBPLV.t8 139.206
R1939 VBPLV.n10 VBPLV.t2 139.206
R1940 VBPLV.n11 VBPLV.t14 139.206
R1941 VBPLV.n12 VBPLV.t7 139.206
R1942 VBPLV.n13 VBPLV.t17 139.206
R1943 VBPLV.n14 VBPLV.t13 139.206
R1944 VBPLV.n15 VBPLV.t0 139.206
R1945 VBPLV.n16 VBPLV.t1 139.206
R1946 VBPLV.n17 VBPLV.t4 139.206
R1947 VBPLV.n18 VBPLV.t5 139.206
R1948 VBPLV.n19 VBPLV.t9 139.206
R1949 VBPLV.n20 VBPLV.t10 139.206
R1950 VBPLV.n21 VBPLV.t18 139.206
R1951 VBPLV.n1 VBPLV.t12 139.206
R1952 VBPLV.n0 VBPLV.t21 139.206
R1953 VBPLV VBPLV.n1 0.804667
R1954 VBPLV VBPLV.n21 0.804667
R1955 VBPLV.n20 VBPLV 0.804667
R1956 VBPLV VBPLV.n19 0.804667
R1957 VBPLV.n18 VBPLV 0.804667
R1958 VBPLV VBPLV.n17 0.804667
R1959 VBPLV.n16 VBPLV 0.804667
R1960 VBPLV VBPLV.n15 0.804667
R1961 VBPLV.n14 VBPLV 0.804667
R1962 VBPLV VBPLV.n13 0.804667
R1963 VBPLV.n12 VBPLV 0.804667
R1964 VBPLV VBPLV.n11 0.804667
R1965 VBPLV.n10 VBPLV 0.804667
R1966 VBPLV VBPLV.n9 0.804667
R1967 VBPLV.n8 VBPLV 0.804667
R1968 VBPLV VBPLV.n7 0.804667
R1969 VBPLV.n6 VBPLV 0.804667
R1970 VBPLV VBPLV.n5 0.804667
R1971 VBPLV.n4 VBPLV 0.804667
R1972 VBPLV VBPLV.n3 0.804667
R1973 VBPLV.n2 VBPLV 0.804667
R1974 VBPLV.n0 VBPLV 0.679667
R1975 VBPLV.n1 VBPLV.n0 0.454667
R1976 VBPLV.n21 VBPLV.n20 0.454667
R1977 VBPLV.n19 VBPLV.n18 0.454667
R1978 VBPLV.n17 VBPLV.n16 0.454667
R1979 VBPLV.n15 VBPLV.n14 0.454667
R1980 VBPLV.n13 VBPLV.n12 0.454667
R1981 VBPLV.n11 VBPLV.n10 0.454667
R1982 VBPLV.n9 VBPLV.n8 0.454667
R1983 VBPLV.n7 VBPLV.n6 0.454667
R1984 VBPLV.n5 VBPLV.n4 0.454667
R1985 VBPLV.n3 VBPLV.n2 0.454667
R1986 VDDH.n24 VDDH.n9 2705.6
R1987 VDDH.n63 VDDH.n9 2705.6
R1988 VDDH.n378 VDDH.n123 1881
R1989 VDDH.n378 VDDH.n377 1881
R1990 VDDH.n377 VDDH.n124 1881
R1991 VDDH.n353 VDDH.n124 1881
R1992 VDDH.n353 VDDH.n352 1881
R1993 VDDH.n352 VDDH.n204 1881
R1994 VDDH.n293 VDDH.n204 1881
R1995 VDDH.n294 VDDH.n293 1881
R1996 VDDH.n309 VDDH.n294 1881
R1997 VDDH.n310 VDDH.n309 1881
R1998 VDDH.t52 VDDH.t34 583.548
R1999 VDDH.t73 VDDH.t40 583.548
R2000 VDDH.t26 VDDH.t5 583.548
R2001 VDDH.t29 VDDH.t21 552.236
R2002 VDDH.n25 VDDH.n10 536.095
R2003 VDDH.n62 VDDH.n10 536.095
R2004 VDDH.t0 VDDH.t62 523.162
R2005 VDDH.t38 VDDH.t4 523.162
R2006 VDDH.t57 VDDH.t25 523.162
R2007 VDDH.t69 VDDH.t10 523.162
R2008 VDDH.t76 VDDH.t70 523.162
R2009 VDDH.t49 VDDH.t83 523.162
R2010 VDDH.n307 VDDH.t74 499.882
R2011 VDDH.n337 VDDH.t128 499.882
R2012 VDDH.n328 VDDH.t53 499.882
R2013 VDDH.n318 VDDH.t79 499.882
R2014 VDDH.n23 VDDH.n8 463.938
R2015 VDDH.n64 VDDH.n8 463.938
R2016 VDDH.t110 VDDH.t29 378.611
R2017 VDDH.t34 VDDH.t88 378.611
R2018 VDDH.t120 VDDH.t52 378.611
R2019 VDDH.t40 VDDH.t96 378.611
R2020 VDDH.t86 VDDH.t73 378.611
R2021 VDDH.t104 VDDH.t26 378.611
R2022 VDDH.t5 VDDH.t94 378.611
R2023 VDDH.t114 VDDH.t14 378.611
R2024 VDDH.n17 VDDH.t61 330.449
R2025 VDDH.n0 VDDH.t82 330.183
R2026 VDDH.n4 VDDH.t30 330.183
R2027 VDDH.n11 VDDH.t45 330.183
R2028 VDDH.n38 VDDH.t31 330.183
R2029 VDDH.n33 VDDH.t12 330.12
R2030 VDDH.n32 VDDH.t46 330.12
R2031 VDDH.n30 VDDH.t36 330.12
R2032 VDDH.n29 VDDH.t13 330.12
R2033 VDDH.n28 VDDH.t81 330.12
R2034 VDDH.n27 VDDH.t60 330.12
R2035 VDDH.n17 VDDH.t37 330.12
R2036 VDDH.n298 VDDH.n297 321.882
R2037 VDDH.n264 VDDH.n254 321.882
R2038 VDDH.n264 VDDH.n248 321.882
R2039 VDDH.n269 VDDH.n248 321.882
R2040 VDDH.n269 VDDH.n245 321.882
R2041 VDDH.n278 VDDH.n245 321.882
R2042 VDDH.n227 VDDH.n211 321.882
R2043 VDDH.n211 VDDH.n208 321.882
R2044 VDDH.n349 VDDH.n208 321.882
R2045 VDDH.n349 VDDH.n209 321.882
R2046 VDDH.n251 VDDH.n209 321.882
R2047 VDDH.n363 VDDH.n162 321.882
R2048 VDDH.n359 VDDH.n162 321.882
R2049 VDDH.n359 VDDH.n200 321.882
R2050 VDDH.n214 VDDH.n200 321.882
R2051 VDDH.n223 VDDH.n214 321.882
R2052 VDDH.n183 VDDH.n173 321.882
R2053 VDDH.n183 VDDH.n167 321.882
R2054 VDDH.n188 VDDH.n167 321.882
R2055 VDDH.n188 VDDH.n164 321.882
R2056 VDDH.n197 VDDH.n164 321.882
R2057 VDDH.n147 VDDH.n131 321.882
R2058 VDDH.n131 VDDH.n128 321.882
R2059 VDDH.n374 VDDH.n128 321.882
R2060 VDDH.n374 VDDH.n129 321.882
R2061 VDDH.n170 VDDH.n129 321.882
R2062 VDDH.n388 VDDH.n86 321.882
R2063 VDDH.n384 VDDH.n86 321.882
R2064 VDDH.n384 VDDH.n88 321.882
R2065 VDDH.n134 VDDH.n88 321.882
R2066 VDDH.n143 VDDH.n134 321.882
R2067 VDDH.n101 VDDH.n98 321.882
R2068 VDDH.n98 VDDH.n95 321.882
R2069 VDDH.n120 VDDH.n95 321.882
R2070 VDDH.n120 VDDH.n96 321.882
R2071 VDDH.n111 VDDH.n96 321.882
R2072 VDDH.n336 VDDH.n243 321.882
R2073 VDDH.n327 VDDH.n285 321.882
R2074 VDDH.n317 VDDH.n292 321.882
R2075 VDDH.n77 VDDH.n2 321.882
R2076 VDDH.n80 VDDH.n2 321.882
R2077 VDDH.n67 VDDH.n6 321.882
R2078 VDDH.n68 VDDH.n67 321.882
R2079 VDDH.n51 VDDH.n13 321.882
R2080 VDDH.n52 VDDH.n51 321.882
R2081 VDDH.n20 VDDH.n14 321.882
R2082 VDDH.n47 VDDH.n14 321.882
R2083 VDDH.n306 VDDH.n305 271.068
R2084 VDDH.n339 VDDH.n338 271.068
R2085 VDDH.n330 VDDH.n329 271.068
R2086 VDDH.n320 VDDH.n319 271.068
R2087 VDDH.t3 VDDH.t2 260.76
R2088 VDDH.n73 VDDH.t7 252.983
R2089 VDDH.n313 VDDH.t80 252.982
R2090 VDDH.n300 VDDH.t75 252.982
R2091 VDDH.n323 VDDH.t54 252.982
R2092 VDDH.n332 VDDH.t129 252.982
R2093 VDDH.n274 VDDH.t51 252.982
R2094 VDDH.n260 VDDH.t66 252.982
R2095 VDDH.n344 VDDH.t78 252.982
R2096 VDDH.n232 VDDH.t56 252.982
R2097 VDDH.n219 VDDH.t68 252.982
R2098 VDDH.n355 VDDH.t59 252.982
R2099 VDDH.n193 VDDH.t72 252.982
R2100 VDDH.n179 VDDH.t131 252.982
R2101 VDDH.n369 VDDH.t42 252.982
R2102 VDDH.n152 VDDH.t16 252.982
R2103 VDDH.n139 VDDH.t64 252.982
R2104 VDDH.n380 VDDH.t33 252.982
R2105 VDDH.n115 VDDH.t20 252.982
R2106 VDDH.n104 VDDH.t133 252.982
R2107 VDDH.n59 VDDH.t24 252.982
R2108 VDDH.n43 VDDH.t44 252.982
R2109 VDDH.n35 VDDH.t48 252.982
R2110 VDDH.n80 VDDH.t22 224.667
R2111 VDDH.t27 VDDH.t28 224.07
R2112 VDDH.t39 VDDH.t3 224.07
R2113 VDDH.t2 VDDH.t35 224.07
R2114 VDDH.t1 VDDH.t11 224.07
R2115 VDDH.n290 VDDH.n289 200.111
R2116 VDDH.n296 VDDH.n295 200.111
R2117 VDDH.n283 VDDH.n282 200.111
R2118 VDDH.n241 VDDH.n240 200.111
R2119 VDDH.n93 VDDH.n92 200.111
R2120 VDDH.n379 VDDH.n91 200.111
R2121 VDDH.n126 VDDH.n125 200.111
R2122 VDDH.n177 VDDH.n176 200.111
R2123 VDDH.n354 VDDH.n203 200.111
R2124 VDDH.n206 VDDH.n205 200.111
R2125 VDDH.n258 VDDH.n257 200.111
R2126 VDDH.n102 VDDH.n101 191.167
R2127 VDDH.n280 VDDH.t110 189.305
R2128 VDDH.t88 VDDH.n280 189.305
R2129 VDDH.n286 VDDH.t120 189.305
R2130 VDDH.t96 VDDH.n286 189.305
R2131 VDDH.n308 VDDH.t86 189.305
R2132 VDDH.n308 VDDH.t104 189.305
R2133 VDDH.n311 VDDH.t94 189.305
R2134 VDDH.n311 VDDH.t114 189.305
R2135 VDDH.n304 VDDH.n298 185
R2136 VDDH.n303 VDDH.n297 185
R2137 VDDH.n307 VDDH.n297 185
R2138 VDDH.n101 VDDH.n100 185
R2139 VDDH.n98 VDDH.n97 185
R2140 VDDH.n99 VDDH.n98 185
R2141 VDDH.n107 VDDH.n95 185
R2142 VDDH.n95 VDDH.n94 185
R2143 VDDH.n120 VDDH.n119 185
R2144 VDDH.n121 VDDH.n120 185
R2145 VDDH.n108 VDDH.n96 185
R2146 VDDH.n109 VDDH.n96 185
R2147 VDDH.n112 VDDH.n111 185
R2148 VDDH.n111 VDDH.n110 185
R2149 VDDH.n389 VDDH.n388 185
R2150 VDDH.n388 VDDH.n387 185
R2151 VDDH.n86 VDDH.n85 185
R2152 VDDH.n386 VDDH.n86 185
R2153 VDDH.n384 VDDH.n383 185
R2154 VDDH.n385 VDDH.n384 185
R2155 VDDH.n89 VDDH.n88 185
R2156 VDDH.n132 VDDH.n88 185
R2157 VDDH.n135 VDDH.n134 185
R2158 VDDH.n134 VDDH.n133 185
R2159 VDDH.n143 VDDH.n142 185
R2160 VDDH.n144 VDDH.n143 185
R2161 VDDH.n148 VDDH.n147 185
R2162 VDDH.n147 VDDH.n146 185
R2163 VDDH.n131 VDDH.n130 185
R2164 VDDH.n145 VDDH.n131 185
R2165 VDDH.n155 VDDH.n128 185
R2166 VDDH.n128 VDDH.n127 185
R2167 VDDH.n374 VDDH.n373 185
R2168 VDDH.n375 VDDH.n374 185
R2169 VDDH.n156 VDDH.n129 185
R2170 VDDH.n168 VDDH.n129 185
R2171 VDDH.n170 VDDH.n169 185
R2172 VDDH.n171 VDDH.n170 185
R2173 VDDH.n174 VDDH.n173 185
R2174 VDDH.n173 VDDH.n172 185
R2175 VDDH.n183 VDDH.n182 185
R2176 VDDH.n184 VDDH.n183 185
R2177 VDDH.n167 VDDH.n166 185
R2178 VDDH.n185 VDDH.n167 185
R2179 VDDH.n189 VDDH.n188 185
R2180 VDDH.n188 VDDH.n187 185
R2181 VDDH.n165 VDDH.n164 185
R2182 VDDH.n164 VDDH.n163 185
R2183 VDDH.n197 VDDH.n196 185
R2184 VDDH.n198 VDDH.n197 185
R2185 VDDH.n364 VDDH.n363 185
R2186 VDDH.n363 VDDH.n362 185
R2187 VDDH.n162 VDDH.n161 185
R2188 VDDH.n361 VDDH.n162 185
R2189 VDDH.n359 VDDH.n358 185
R2190 VDDH.n360 VDDH.n359 185
R2191 VDDH.n201 VDDH.n200 185
R2192 VDDH.n212 VDDH.n200 185
R2193 VDDH.n215 VDDH.n214 185
R2194 VDDH.n214 VDDH.n213 185
R2195 VDDH.n223 VDDH.n222 185
R2196 VDDH.n224 VDDH.n223 185
R2197 VDDH.n228 VDDH.n227 185
R2198 VDDH.n227 VDDH.n226 185
R2199 VDDH.n211 VDDH.n210 185
R2200 VDDH.n225 VDDH.n211 185
R2201 VDDH.n235 VDDH.n208 185
R2202 VDDH.n208 VDDH.n207 185
R2203 VDDH.n349 VDDH.n348 185
R2204 VDDH.n350 VDDH.n349 185
R2205 VDDH.n236 VDDH.n209 185
R2206 VDDH.n249 VDDH.n209 185
R2207 VDDH.n251 VDDH.n250 185
R2208 VDDH.n252 VDDH.n251 185
R2209 VDDH.n255 VDDH.n254 185
R2210 VDDH.n254 VDDH.n253 185
R2211 VDDH.n264 VDDH.n263 185
R2212 VDDH.n265 VDDH.n264 185
R2213 VDDH.n248 VDDH.n247 185
R2214 VDDH.n266 VDDH.n248 185
R2215 VDDH.n270 VDDH.n269 185
R2216 VDDH.n269 VDDH.n268 185
R2217 VDDH.n246 VDDH.n245 185
R2218 VDDH.n245 VDDH.n244 185
R2219 VDDH.n278 VDDH.n277 185
R2220 VDDH.n279 VDDH.n278 185
R2221 VDDH.n243 VDDH.n242 185
R2222 VDDH.n336 VDDH.n335 185
R2223 VDDH.n337 VDDH.n336 185
R2224 VDDH.n285 VDDH.n284 185
R2225 VDDH.n327 VDDH.n326 185
R2226 VDDH.n328 VDDH.n327 185
R2227 VDDH.n292 VDDH.n291 185
R2228 VDDH.n317 VDDH.n316 185
R2229 VDDH.n318 VDDH.n317 185
R2230 VDDH.n20 VDDH.n19 185
R2231 VDDH.n21 VDDH.n20 185
R2232 VDDH.n15 VDDH.n14 185
R2233 VDDH.n18 VDDH.n14 185
R2234 VDDH.n47 VDDH.n46 185
R2235 VDDH.n48 VDDH.n47 185
R2236 VDDH.n39 VDDH.n13 185
R2237 VDDH.n49 VDDH.n13 185
R2238 VDDH.n51 VDDH.n12 185
R2239 VDDH.n51 VDDH.n50 185
R2240 VDDH.n53 VDDH.n52 185
R2241 VDDH.n52 VDDH.n7 185
R2242 VDDH.n55 VDDH.n6 185
R2243 VDDH.n65 VDDH.n6 185
R2244 VDDH.n67 VDDH.n5 185
R2245 VDDH.n67 VDDH.n66 185
R2246 VDDH.n69 VDDH.n68 185
R2247 VDDH.n68 VDDH.n3 185
R2248 VDDH.n77 VDDH.n76 185
R2249 VDDH.n78 VDDH.n77 185
R2250 VDDH.n2 VDDH.n1 185
R2251 VDDH.n79 VDDH.n2 185
R2252 VDDH.n81 VDDH.n80 185
R2253 VDDH.t11 VDDH.n21 164.69
R2254 VDDH.n23 VDDH.t27 132.345
R2255 VDDH.t35 VDDH.n22 132.345
R2256 VDDH.n110 VDDH.n109 92.2149
R2257 VDDH.n144 VDDH.n133 92.2149
R2258 VDDH.n171 VDDH.n168 92.2149
R2259 VDDH.n198 VDDH.n163 92.2149
R2260 VDDH.n224 VDDH.n213 92.2149
R2261 VDDH.n252 VDDH.n249 92.2149
R2262 VDDH.n279 VDDH.n244 92.2149
R2263 VDDH.n23 VDDH.t39 91.7246
R2264 VDDH.n22 VDDH.t1 91.7246
R2265 VDDH.n100 VDDH.t132 89.3332
R2266 VDDH.n387 VDDH.t32 89.3332
R2267 VDDH.n146 VDDH.t15 89.3332
R2268 VDDH.n172 VDDH.t130 89.3332
R2269 VDDH.n362 VDDH.t58 89.3332
R2270 VDDH.n226 VDDH.t55 89.3332
R2271 VDDH.n253 VDDH.t65 89.3332
R2272 VDDH.n306 VDDH.n298 86.068
R2273 VDDH.n338 VDDH.n243 86.068
R2274 VDDH.n329 VDDH.n285 86.068
R2275 VDDH.n319 VDDH.n292 86.068
R2276 VDDH.n100 VDDH.t18 84.5303
R2277 VDDH.n387 VDDH.t62 84.5303
R2278 VDDH.n146 VDDH.t38 84.5303
R2279 VDDH.n172 VDDH.t57 84.5303
R2280 VDDH.n362 VDDH.t69 84.5303
R2281 VDDH.n226 VDDH.t76 84.5303
R2282 VDDH.n253 VDDH.t49 84.5303
R2283 VDDH.n110 VDDH.t0 82.6092
R2284 VDDH.t4 VDDH.n144 82.6092
R2285 VDDH.t25 VDDH.n171 82.6092
R2286 VDDH.t10 VDDH.n198 82.6092
R2287 VDDH.t70 VDDH.n224 82.6092
R2288 VDDH.t83 VDDH.n252 82.6092
R2289 VDDH.t21 VDDH.n279 82.6092
R2290 VDDH.n49 VDDH.n48 78.8324
R2291 VDDH.n78 VDDH.n3 75.3176
R2292 VDDH.n64 VDDH.n7 61.7605
R2293 VDDH.t84 VDDH.n94 59.5556
R2294 VDDH.t90 VDDH.n385 59.5556
R2295 VDDH.t108 VDDH.n127 59.5556
R2296 VDDH.n185 VDDH.t118 59.5556
R2297 VDDH.t126 VDDH.n360 59.5556
R2298 VDDH.t92 VDDH.n207 59.5556
R2299 VDDH.n266 VDDH.t98 59.5556
R2300 VDDH.n121 VDDH.t102 57.6345
R2301 VDDH.t106 VDDH.n132 57.6345
R2302 VDDH.n375 VDDH.t116 57.6345
R2303 VDDH.n187 VDDH.t124 57.6345
R2304 VDDH.t100 VDDH.n212 57.6345
R2305 VDDH.n350 VDDH.t112 57.6345
R2306 VDDH.n268 VDDH.t122 57.6345
R2307 VDDH.n307 VDDH.n306 49.4675
R2308 VDDH.n338 VDDH.n337 49.4675
R2309 VDDH.n329 VDDH.n328 49.4675
R2310 VDDH.n319 VDDH.n318 49.4675
R2311 VDDH.n21 VDDH.n18 48.2035
R2312 VDDH.n50 VDDH.n49 48.2035
R2313 VDDH.n66 VDDH.n65 48.2035
R2314 VDDH.n79 VDDH.n78 48.2035
R2315 VDDH.n122 VDDH.n121 47.0682
R2316 VDDH.n132 VDDH.n87 47.0682
R2317 VDDH.n376 VDDH.n375 47.0682
R2318 VDDH.n187 VDDH.n186 47.0682
R2319 VDDH.n212 VDDH.n199 47.0682
R2320 VDDH.n351 VDDH.n350 47.0682
R2321 VDDH.n268 VDDH.n267 47.0682
R2322 VDDH.n122 VDDH.n94 45.1471
R2323 VDDH.n385 VDDH.n87 45.1471
R2324 VDDH.n376 VDDH.n127 45.1471
R2325 VDDH.n186 VDDH.n185 45.1471
R2326 VDDH.n360 VDDH.n199 45.1471
R2327 VDDH.n351 VDDH.n207 45.1471
R2328 VDDH.n267 VDDH.n266 45.1471
R2329 VDDH.t17 VDDH.n7 39.6675
R2330 VDDH.t9 VDDH.n3 39.6675
R2331 VDDH.n48 VDDH.t8 36.1527
R2332 VDDH.n305 VDDH.n304 36.1417
R2333 VDDH.n304 VDDH.n303 36.1417
R2334 VDDH.n263 VDDH.n255 36.1417
R2335 VDDH.n263 VDDH.n247 36.1417
R2336 VDDH.n270 VDDH.n247 36.1417
R2337 VDDH.n270 VDDH.n246 36.1417
R2338 VDDH.n277 VDDH.n246 36.1417
R2339 VDDH.n228 VDDH.n210 36.1417
R2340 VDDH.n235 VDDH.n210 36.1417
R2341 VDDH.n348 VDDH.n235 36.1417
R2342 VDDH.n348 VDDH.n236 36.1417
R2343 VDDH.n250 VDDH.n236 36.1417
R2344 VDDH.n364 VDDH.n161 36.1417
R2345 VDDH.n358 VDDH.n161 36.1417
R2346 VDDH.n358 VDDH.n201 36.1417
R2347 VDDH.n215 VDDH.n201 36.1417
R2348 VDDH.n222 VDDH.n215 36.1417
R2349 VDDH.n182 VDDH.n174 36.1417
R2350 VDDH.n182 VDDH.n166 36.1417
R2351 VDDH.n189 VDDH.n166 36.1417
R2352 VDDH.n189 VDDH.n165 36.1417
R2353 VDDH.n196 VDDH.n165 36.1417
R2354 VDDH.n148 VDDH.n130 36.1417
R2355 VDDH.n155 VDDH.n130 36.1417
R2356 VDDH.n373 VDDH.n155 36.1417
R2357 VDDH.n373 VDDH.n156 36.1417
R2358 VDDH.n169 VDDH.n156 36.1417
R2359 VDDH.n389 VDDH.n85 36.1417
R2360 VDDH.n383 VDDH.n85 36.1417
R2361 VDDH.n383 VDDH.n89 36.1417
R2362 VDDH.n135 VDDH.n89 36.1417
R2363 VDDH.n142 VDDH.n135 36.1417
R2364 VDDH.n107 VDDH.n97 36.1417
R2365 VDDH.n119 VDDH.n107 36.1417
R2366 VDDH.n119 VDDH.n108 36.1417
R2367 VDDH.n112 VDDH.n108 36.1417
R2368 VDDH.n339 VDDH.n242 36.1417
R2369 VDDH.n335 VDDH.n242 36.1417
R2370 VDDH.n330 VDDH.n284 36.1417
R2371 VDDH.n326 VDDH.n284 36.1417
R2372 VDDH.n320 VDDH.n291 36.1417
R2373 VDDH.n316 VDDH.n291 36.1417
R2374 VDDH.n76 VDDH.n1 36.1417
R2375 VDDH.n81 VDDH.n1 36.1417
R2376 VDDH.n55 VDDH.n5 36.1417
R2377 VDDH.n69 VDDH.n5 36.1417
R2378 VDDH.n39 VDDH.n12 36.1417
R2379 VDDH.n53 VDDH.n12 36.1417
R2380 VDDH.n19 VDDH.n15 36.1417
R2381 VDDH.n46 VDDH.n15 36.1417
R2382 VDDH.n99 VDDH.t84 32.6598
R2383 VDDH.n386 VDDH.t90 32.6598
R2384 VDDH.n145 VDDH.t108 32.6598
R2385 VDDH.t118 VDDH.n184 32.6598
R2386 VDDH.n361 VDDH.t126 32.6598
R2387 VDDH.n225 VDDH.t92 32.6598
R2388 VDDH.t98 VDDH.n265 32.6598
R2389 VDDH.t19 VDDH.t102 31.6992
R2390 VDDH.t63 VDDH.t106 31.6992
R2391 VDDH.t41 VDDH.t116 31.6992
R2392 VDDH.t124 VDDH.t71 31.6992
R2393 VDDH.t67 VDDH.t100 31.6992
R2394 VDDH.t77 VDDH.t112 31.6992
R2395 VDDH.t122 VDDH.t50 31.6992
R2396 VDDH.n289 VDDH.t95 27.6955
R2397 VDDH.n289 VDDH.t115 27.6955
R2398 VDDH.n295 VDDH.t87 27.6955
R2399 VDDH.n295 VDDH.t105 27.6955
R2400 VDDH.n282 VDDH.t121 27.6955
R2401 VDDH.n282 VDDH.t97 27.6955
R2402 VDDH.n240 VDDH.t111 27.6955
R2403 VDDH.n240 VDDH.t89 27.6955
R2404 VDDH.n92 VDDH.t85 27.6955
R2405 VDDH.n92 VDDH.t103 27.6955
R2406 VDDH.n91 VDDH.t91 27.6955
R2407 VDDH.n91 VDDH.t107 27.6955
R2408 VDDH.n125 VDDH.t109 27.6955
R2409 VDDH.n125 VDDH.t117 27.6955
R2410 VDDH.n176 VDDH.t119 27.6955
R2411 VDDH.n176 VDDH.t125 27.6955
R2412 VDDH.n203 VDDH.t127 27.6955
R2413 VDDH.n203 VDDH.t101 27.6955
R2414 VDDH.n205 VDDH.t93 27.6955
R2415 VDDH.n205 VDDH.t113 27.6955
R2416 VDDH.n257 VDDH.t99 27.6955
R2417 VDDH.n257 VDDH.t123 27.6955
R2418 VDDH.n22 VDDH.n8 16.4402
R2419 VDDH.n310 VDDH.n290 16.2626
R2420 VDDH.n309 VDDH.n296 16.2626
R2421 VDDH.n294 VDDH.n283 16.2626
R2422 VDDH.n293 VDDH.n241 16.2626
R2423 VDDH.n258 VDDH.n204 16.2626
R2424 VDDH.n352 VDDH.n206 16.2626
R2425 VDDH.n354 VDDH.n353 16.2626
R2426 VDDH.n177 VDDH.n124 16.2626
R2427 VDDH.n377 VDDH.n126 16.2626
R2428 VDDH.n379 VDDH.n378 16.2626
R2429 VDDH.n123 VDDH.n93 16.2626
R2430 VDDH.n309 VDDH.n308 15.4172
R2431 VDDH.n294 VDDH.n286 15.4172
R2432 VDDH.n293 VDDH.n280 15.4172
R2433 VDDH.n267 VDDH.n204 15.4172
R2434 VDDH.n352 VDDH.n351 15.4172
R2435 VDDH.n353 VDDH.n199 15.4172
R2436 VDDH.n186 VDDH.n124 15.4172
R2437 VDDH.n377 VDDH.n376 15.4172
R2438 VDDH.n378 VDDH.n87 15.4172
R2439 VDDH.n123 VDDH.n122 15.4172
R2440 VDDH.n311 VDDH.n310 15.4172
R2441 VDDH.n65 VDDH.n64 13.5576
R2442 VDDH.n308 VDDH.n307 11.31
R2443 VDDH.n337 VDDH.n280 11.31
R2444 VDDH.n328 VDDH.n286 11.31
R2445 VDDH.n318 VDDH.n311 11.31
R2446 VDDH.t47 VDDH.t8 10.5449
R2447 VDDH.n63 VDDH.n62 9.73734
R2448 VDDH.n64 VDDH.n63 9.73734
R2449 VDDH.n10 VDDH.n9 9.73734
R2450 VDDH.n22 VDDH.n9 9.73734
R2451 VDDH.n25 VDDH.n24 9.73734
R2452 VDDH.n24 VDDH.n23 9.73734
R2453 VDDH.n107 VDDH.n106 9.3005
R2454 VDDH.n119 VDDH.n118 9.3005
R2455 VDDH.n117 VDDH.n108 9.3005
R2456 VDDH.n113 VDDH.n112 9.3005
R2457 VDDH.n390 VDDH.n389 9.3005
R2458 VDDH.n85 VDDH.n84 9.3005
R2459 VDDH.n383 VDDH.n382 9.3005
R2460 VDDH.n136 VDDH.n89 9.3005
R2461 VDDH.n137 VDDH.n135 9.3005
R2462 VDDH.n142 VDDH.n141 9.3005
R2463 VDDH.n149 VDDH.n148 9.3005
R2464 VDDH.n150 VDDH.n130 9.3005
R2465 VDDH.n155 VDDH.n154 9.3005
R2466 VDDH.n373 VDDH.n372 9.3005
R2467 VDDH.n371 VDDH.n156 9.3005
R2468 VDDH.n169 VDDH.n157 9.3005
R2469 VDDH.n174 VDDH.n158 9.3005
R2470 VDDH.n182 VDDH.n181 9.3005
R2471 VDDH.n175 VDDH.n166 9.3005
R2472 VDDH.n190 VDDH.n189 9.3005
R2473 VDDH.n191 VDDH.n165 9.3005
R2474 VDDH.n196 VDDH.n195 9.3005
R2475 VDDH.n365 VDDH.n364 9.3005
R2476 VDDH.n161 VDDH.n160 9.3005
R2477 VDDH.n358 VDDH.n357 9.3005
R2478 VDDH.n216 VDDH.n201 9.3005
R2479 VDDH.n217 VDDH.n215 9.3005
R2480 VDDH.n222 VDDH.n221 9.3005
R2481 VDDH.n229 VDDH.n228 9.3005
R2482 VDDH.n230 VDDH.n210 9.3005
R2483 VDDH.n235 VDDH.n234 9.3005
R2484 VDDH.n348 VDDH.n347 9.3005
R2485 VDDH.n346 VDDH.n236 9.3005
R2486 VDDH.n250 VDDH.n237 9.3005
R2487 VDDH.n255 VDDH.n238 9.3005
R2488 VDDH.n263 VDDH.n262 9.3005
R2489 VDDH.n256 VDDH.n247 9.3005
R2490 VDDH.n271 VDDH.n270 9.3005
R2491 VDDH.n272 VDDH.n246 9.3005
R2492 VDDH.n277 VDDH.n276 9.3005
R2493 VDDH.n340 VDDH.n339 9.3005
R2494 VDDH.n242 VDDH.n241 9.3005
R2495 VDDH.n335 VDDH.n334 9.3005
R2496 VDDH.n331 VDDH.n330 9.3005
R2497 VDDH.n284 VDDH.n283 9.3005
R2498 VDDH.n326 VDDH.n325 9.3005
R2499 VDDH.n305 VDDH.n288 9.3005
R2500 VDDH.n304 VDDH.n296 9.3005
R2501 VDDH.n303 VDDH.n302 9.3005
R2502 VDDH.n321 VDDH.n320 9.3005
R2503 VDDH.n291 VDDH.n290 9.3005
R2504 VDDH.n316 VDDH.n315 9.3005
R2505 VDDH.n104 VDDH.n103 9.3005
R2506 VDDH.n105 VDDH.n104 9.3005
R2507 VDDH.n116 VDDH.n115 9.3005
R2508 VDDH.n115 VDDH.n114 9.3005
R2509 VDDH.n380 VDDH.n90 9.3005
R2510 VDDH.n381 VDDH.n380 9.3005
R2511 VDDH.n139 VDDH.n138 9.3005
R2512 VDDH.n140 VDDH.n139 9.3005
R2513 VDDH.n152 VDDH.n151 9.3005
R2514 VDDH.n153 VDDH.n152 9.3005
R2515 VDDH.n370 VDDH.n369 9.3005
R2516 VDDH.n369 VDDH.n368 9.3005
R2517 VDDH.n180 VDDH.n179 9.3005
R2518 VDDH.n179 VDDH.n178 9.3005
R2519 VDDH.n193 VDDH.n192 9.3005
R2520 VDDH.n194 VDDH.n193 9.3005
R2521 VDDH.n355 VDDH.n202 9.3005
R2522 VDDH.n356 VDDH.n355 9.3005
R2523 VDDH.n219 VDDH.n218 9.3005
R2524 VDDH.n220 VDDH.n219 9.3005
R2525 VDDH.n232 VDDH.n231 9.3005
R2526 VDDH.n233 VDDH.n232 9.3005
R2527 VDDH.n345 VDDH.n344 9.3005
R2528 VDDH.n344 VDDH.n343 9.3005
R2529 VDDH.n261 VDDH.n260 9.3005
R2530 VDDH.n260 VDDH.n259 9.3005
R2531 VDDH.n274 VDDH.n273 9.3005
R2532 VDDH.n275 VDDH.n274 9.3005
R2533 VDDH.n332 VDDH.n281 9.3005
R2534 VDDH.n333 VDDH.n332 9.3005
R2535 VDDH.n323 VDDH.n287 9.3005
R2536 VDDH.n324 VDDH.n323 9.3005
R2537 VDDH.n300 VDDH.n299 9.3005
R2538 VDDH.n301 VDDH.n300 9.3005
R2539 VDDH.n313 VDDH.n312 9.3005
R2540 VDDH.n314 VDDH.n313 9.3005
R2541 VDDH.n36 VDDH.n35 9.3005
R2542 VDDH.n35 VDDH.n34 9.3005
R2543 VDDH.n43 VDDH.n42 9.3005
R2544 VDDH.n44 VDDH.n43 9.3005
R2545 VDDH.n59 VDDH.n58 9.3005
R2546 VDDH.n60 VDDH.n59 9.3005
R2547 VDDH.n74 VDDH.n73 9.3005
R2548 VDDH.n73 VDDH.n71 9.3005
R2549 VDDH.n19 VDDH.n16 9.3005
R2550 VDDH.n37 VDDH.n15 9.3005
R2551 VDDH.n46 VDDH.n45 9.3005
R2552 VDDH.n40 VDDH.n39 9.3005
R2553 VDDH.n41 VDDH.n12 9.3005
R2554 VDDH.n54 VDDH.n53 9.3005
R2555 VDDH.n56 VDDH.n55 9.3005
R2556 VDDH.n57 VDDH.n5 9.3005
R2557 VDDH.n70 VDDH.n69 9.3005
R2558 VDDH.n76 VDDH.n75 9.3005
R2559 VDDH.n72 VDDH.n1 9.3005
R2560 VDDH.n82 VDDH.n81 9.3005
R2561 VDDH.t43 VDDH.t17 7.0301
R2562 VDDH.t23 VDDH.t9 7.0301
R2563 VDDH.t22 VDDH.t6 7.0301
R2564 VDDH.n102 VDDH.n97 6.13579
R2565 VDDH VDDH.n322 3.7711
R2566 VDDH VDDH.n239 3.7711
R2567 VDDH.n341 VDDH 3.7711
R2568 VDDH VDDH.n342 3.7711
R2569 VDDH VDDH.n159 3.7711
R2570 VDDH.n366 VDDH 3.7711
R2571 VDDH VDDH.n367 3.7711
R2572 VDDH VDDH.n83 3.7711
R2573 VDDH.n391 VDDH 3.7711
R2574 VDDH.t132 VDDH.n99 2.8822
R2575 VDDH.n109 VDDH.t19 2.8822
R2576 VDDH.t32 VDDH.n386 2.8822
R2577 VDDH.n133 VDDH.t63 2.8822
R2578 VDDH.t15 VDDH.n145 2.8822
R2579 VDDH.n168 VDDH.t41 2.8822
R2580 VDDH.n184 VDDH.t130 2.8822
R2581 VDDH.t71 VDDH.n163 2.8822
R2582 VDDH.t58 VDDH.n361 2.8822
R2583 VDDH.n213 VDDH.t67 2.8822
R2584 VDDH.t55 VDDH.n225 2.8822
R2585 VDDH.n249 VDDH.t77 2.8822
R2586 VDDH.n265 VDDH.t65 2.8822
R2587 VDDH.t50 VDDH.n244 2.8822
R2588 VDDH.n103 VDDH.n102 1.60272
R2589 VDDH.n18 VDDH.t47 1.50684
R2590 VDDH.n50 VDDH.t43 1.50684
R2591 VDDH.n66 VDDH.t23 1.50684
R2592 VDDH.t6 VDDH.n79 1.50684
R2593 VDDH VDDH.n391 0.861477
R2594 VDDH.n391 VDDH.n83 0.61925
R2595 VDDH.n367 VDDH.n83 0.61925
R2596 VDDH.n367 VDDH.n366 0.61925
R2597 VDDH.n366 VDDH.n159 0.61925
R2598 VDDH.n342 VDDH.n159 0.61925
R2599 VDDH.n342 VDDH.n341 0.61925
R2600 VDDH.n341 VDDH.n239 0.61925
R2601 VDDH.n322 VDDH.n239 0.61925
R2602 VDDH.n322 VDDH 0.56425
R2603 VDDH.n26 VDDH.n25 0.517167
R2604 VDDH.n31 VDDH.n10 0.517167
R2605 VDDH.n62 VDDH.n61 0.517167
R2606 VDDH.n28 VDDH.n27 0.328024
R2607 VDDH.n30 VDDH.n29 0.328024
R2608 VDDH.n33 VDDH.n32 0.328024
R2609 VDDH VDDH.n28 0.238481
R2610 VDDH VDDH.n33 0.238481
R2611 VDDH.n26 VDDH.n17 0.204627
R2612 VDDH.n31 VDDH.n30 0.204627
R2613 VDDH VDDH.n340 0.195324
R2614 VDDH VDDH.n331 0.195324
R2615 VDDH VDDH.n288 0.195324
R2616 VDDH VDDH.n321 0.195324
R2617 VDDH.n29 VDDH 0.16296
R2618 VDDH VDDH.n390 0.1255
R2619 VDDH.n149 VDDH 0.1255
R2620 VDDH VDDH.n158 0.1255
R2621 VDDH VDDH.n365 0.1255
R2622 VDDH.n229 VDDH 0.1255
R2623 VDDH VDDH.n238 0.1255
R2624 VDDH.n27 VDDH.n26 0.123897
R2625 VDDH.n32 VDDH.n31 0.123897
R2626 VDDH VDDH.n44 0.0503047
R2627 VDDH.n118 VDDH.n117 0.047375
R2628 VDDH.n390 VDDH.n84 0.047375
R2629 VDDH.n137 VDDH.n136 0.047375
R2630 VDDH.n150 VDDH.n149 0.047375
R2631 VDDH.n372 VDDH.n371 0.047375
R2632 VDDH.n181 VDDH.n158 0.047375
R2633 VDDH.n191 VDDH.n190 0.047375
R2634 VDDH.n365 VDDH.n160 0.047375
R2635 VDDH.n217 VDDH.n216 0.047375
R2636 VDDH.n230 VDDH.n229 0.047375
R2637 VDDH.n347 VDDH.n346 0.047375
R2638 VDDH.n262 VDDH.n238 0.047375
R2639 VDDH.n272 VDDH.n271 0.047375
R2640 VDDH.n340 VDDH.n241 0.047375
R2641 VDDH.n331 VDDH.n283 0.047375
R2642 VDDH.n296 VDDH.n288 0.047375
R2643 VDDH.n321 VDDH.n290 0.047375
R2644 VDDH.n71 VDDH 0.0468867
R2645 VDDH.n54 VDDH.n11 0.0390742
R2646 VDDH.n70 VDDH.n4 0.0390742
R2647 VDDH.n82 VDDH.n0 0.0390742
R2648 VDDH.n61 VDDH 0.0371211
R2649 VDDH.n45 VDDH.n38 0.0356562
R2650 VDDH.n106 VDDH.n103 0.0322383
R2651 VDDH.n116 VDDH.n113 0.0322383
R2652 VDDH.n382 VDDH.n90 0.0322383
R2653 VDDH.n141 VDDH.n138 0.0322383
R2654 VDDH.n154 VDDH.n151 0.0322383
R2655 VDDH.n370 VDDH.n157 0.0322383
R2656 VDDH.n180 VDDH.n175 0.0322383
R2657 VDDH.n195 VDDH.n192 0.0322383
R2658 VDDH.n357 VDDH.n202 0.0322383
R2659 VDDH.n221 VDDH.n218 0.0322383
R2660 VDDH.n234 VDDH.n231 0.0322383
R2661 VDDH.n345 VDDH.n237 0.0322383
R2662 VDDH.n261 VDDH.n256 0.0322383
R2663 VDDH.n276 VDDH.n273 0.0322383
R2664 VDDH.n334 VDDH.n281 0.0322383
R2665 VDDH.n325 VDDH.n287 0.0322383
R2666 VDDH.n302 VDDH.n299 0.0322383
R2667 VDDH.n315 VDDH.n312 0.0322383
R2668 VDDH.n36 VDDH.n16 0.0322383
R2669 VDDH.n42 VDDH.n40 0.0322383
R2670 VDDH.n58 VDDH.n56 0.0322383
R2671 VDDH.n75 VDDH.n74 0.0322383
R2672 VDDH.n118 VDDH 0.0239375
R2673 VDDH.n136 VDDH 0.0239375
R2674 VDDH.n372 VDDH 0.0239375
R2675 VDDH.n190 VDDH 0.0239375
R2676 VDDH.n216 VDDH 0.0239375
R2677 VDDH.n347 VDDH 0.0239375
R2678 VDDH.n271 VDDH 0.0239375
R2679 VDDH.n45 VDDH 0.0239375
R2680 VDDH VDDH.n54 0.0239375
R2681 VDDH VDDH.n70 0.0239375
R2682 VDDH VDDH.n82 0.0239375
R2683 VDDH.n34 VDDH 0.0231237
R2684 VDDH.n333 VDDH 0.0205195
R2685 VDDH.n324 VDDH 0.0205195
R2686 VDDH.n301 VDDH 0.0205195
R2687 VDDH.n314 VDDH 0.0205195
R2688 VDDH.n105 VDDH.n93 0.0200312
R2689 VDDH.n381 VDDH.n379 0.0200312
R2690 VDDH.n153 VDDH.n126 0.0200312
R2691 VDDH.n178 VDDH.n177 0.0200312
R2692 VDDH.n356 VDDH.n354 0.0200312
R2693 VDDH.n233 VDDH.n206 0.0200312
R2694 VDDH.n259 VDDH.n258 0.0200312
R2695 VDDH.n117 VDDH.n116 0.0156367
R2696 VDDH.n114 VDDH 0.0156367
R2697 VDDH.n90 VDDH.n84 0.0156367
R2698 VDDH.n138 VDDH.n137 0.0156367
R2699 VDDH.n140 VDDH 0.0156367
R2700 VDDH.n151 VDDH.n150 0.0156367
R2701 VDDH.n371 VDDH.n370 0.0156367
R2702 VDDH.n368 VDDH 0.0156367
R2703 VDDH.n181 VDDH.n180 0.0156367
R2704 VDDH.n192 VDDH.n191 0.0156367
R2705 VDDH.n194 VDDH 0.0156367
R2706 VDDH.n202 VDDH.n160 0.0156367
R2707 VDDH.n218 VDDH.n217 0.0156367
R2708 VDDH.n220 VDDH 0.0156367
R2709 VDDH.n231 VDDH.n230 0.0156367
R2710 VDDH.n346 VDDH.n345 0.0156367
R2711 VDDH.n343 VDDH 0.0156367
R2712 VDDH.n262 VDDH.n261 0.0156367
R2713 VDDH.n273 VDDH.n272 0.0156367
R2714 VDDH.n275 VDDH 0.0156367
R2715 VDDH.n281 VDDH.n241 0.0156367
R2716 VDDH.n287 VDDH.n283 0.0156367
R2717 VDDH.n299 VDDH.n296 0.0156367
R2718 VDDH.n312 VDDH.n290 0.0156367
R2719 VDDH.n37 VDDH.n36 0.0156367
R2720 VDDH.n42 VDDH.n41 0.0156367
R2721 VDDH.n58 VDDH.n57 0.0156367
R2722 VDDH.n74 VDDH.n72 0.0156367
R2723 VDDH.n38 VDDH.n37 0.0122188
R2724 VDDH.n61 VDDH.n60 0.0102656
R2725 VDDH.n41 VDDH.n11 0.00880078
R2726 VDDH.n57 VDDH.n4 0.00880078
R2727 VDDH.n72 VDDH.n0 0.00880078
R2728 VDDH.n106 VDDH.n105 0.00391797
R2729 VDDH.n114 VDDH.n113 0.00391797
R2730 VDDH.n382 VDDH.n381 0.00391797
R2731 VDDH.n141 VDDH.n140 0.00391797
R2732 VDDH.n154 VDDH.n153 0.00391797
R2733 VDDH.n368 VDDH.n157 0.00391797
R2734 VDDH.n178 VDDH.n175 0.00391797
R2735 VDDH.n195 VDDH.n194 0.00391797
R2736 VDDH.n357 VDDH.n356 0.00391797
R2737 VDDH.n221 VDDH.n220 0.00391797
R2738 VDDH.n234 VDDH.n233 0.00391797
R2739 VDDH.n343 VDDH.n237 0.00391797
R2740 VDDH.n259 VDDH.n256 0.00391797
R2741 VDDH.n276 VDDH.n275 0.00391797
R2742 VDDH.n334 VDDH.n333 0.00391797
R2743 VDDH.n325 VDDH.n324 0.00391797
R2744 VDDH.n302 VDDH.n301 0.00391797
R2745 VDDH.n315 VDDH.n314 0.00391797
R2746 VDDH.n34 VDDH.n16 0.00391797
R2747 VDDH.n44 VDDH.n40 0.00391797
R2748 VDDH.n60 VDDH.n56 0.00391797
R2749 VDDH.n75 VDDH.n71 0.00391797
R2750 VDDH VDDH.n93 0.000988281
R2751 VDDH.n379 VDDH 0.000988281
R2752 VDDH VDDH.n126 0.000988281
R2753 VDDH.n177 VDDH 0.000988281
R2754 VDDH.n354 VDDH 0.000988281
R2755 VDDH VDDH.n206 0.000988281
R2756 VDDH.n258 VDDH 0.000988281
R2757 a_16484_n199.t0 a_16484_n199.t1 55.3905
R2758 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t6 732.773
R2759 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t8 212.081
R2760 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t5 212.081
R2761 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 208.965
R2762 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 186.001
R2763 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t7 139.78
R2764 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t4 139.78
R2765 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 96.8352
R2766 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 61.346
R2767 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 28.4963
R2768 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t2 26.5955
R2769 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t3 26.5955
R2770 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t1 24.9236
R2771 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t0 24.9236
R2772 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 12.5445
R2773 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 11.2645
R2774 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 9.65467
R2775 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 9.30258
R2776 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 6.1445
R2777 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 4.8645
R2778 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 4.65505
R2779 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 3.0725
R2780 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 2.0485
R2781 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 1.55202
R2782 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t4 732.702
R2783 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 208.965
R2784 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 96.8352
R2785 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 37.042
R2786 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t2 26.5955
R2787 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t3 26.5955
R2788 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t0 24.9236
R2789 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t1 24.9236
R2790 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 13.0565
R2791 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 11.2645
R2792 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 6.1445
R2793 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 4.65505
R2794 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 4.3525
R2795 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 2.0485
R2796 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 1.55202
R2797 VBPDEC.n4 VBPDEC.t11 120.969
R2798 VBPDEC.n5 VBPDEC.t2 120.969
R2799 VBPDEC.n6 VBPDEC.t8 120.969
R2800 VBPDEC.n7 VBPDEC.t3 120.969
R2801 VBPDEC.n8 VBPDEC.t0 120.969
R2802 VBPDEC.n9 VBPDEC.t9 120.969
R2803 VBPDEC.n10 VBPDEC.t6 120.969
R2804 VBPDEC.n11 VBPDEC.t1 120.969
R2805 VBPDEC.n3 VBPDEC.t10 120.969
R2806 VBPDEC.n2 VBPDEC.t4 120.969
R2807 VBPDEC.n1 VBPDEC.t7 120.969
R2808 VBPDEC.n0 VBPDEC.t5 120.969
R2809 VBPDEC.n1 VBPDEC.n0 0.713
R2810 VBPDEC.n2 VBPDEC.n1 0.713
R2811 VBPDEC.n3 VBPDEC.n2 0.713
R2812 VBPDEC.n11 VBPDEC.n10 0.713
R2813 VBPDEC.n10 VBPDEC.n9 0.713
R2814 VBPDEC.n9 VBPDEC.n8 0.713
R2815 VBPDEC.n7 VBPDEC.n6 0.713
R2816 VBPDEC.n6 VBPDEC.n5 0.713
R2817 VBPDEC.n5 VBPDEC.n4 0.713
R2818 VBPDEC VBPDEC.n11 0.690083
R2819 VBPDEC VBPDEC.n7 0.690083
R2820 VBPDEC.n0 VBPDEC 0.533833
R2821 VBPDEC VBPDEC.n3 0.140083
R2822 VBPDEC.n8 VBPDEC 0.140083
R2823 VBPDEC.n4 VBPDEC 0.140083
R2824 a_22706_943.t0 a_22706_943.t1 65.941
R2825 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t0 227.856
R2826 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n0 152.333
R2827 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t2 140.382
R2828 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t3 114.031
R2829 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t1 83.3993
R2830 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t4 81.5883
R2831 lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n1 14.4422
R2832 lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n3 7.56882
R2833 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n2 5.08175
R2834 lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R2835 a_14504_n199.t0 a_14504_n199.t1 55.3905
R2836 a_13908_n296.n0 a_13908_n296.t1 228.04
R2837 a_13908_n296.n0 a_13908_n296.t2 145.648
R2838 a_13908_n296.t0 a_13908_n296.n0 83.2159
R2839 VDD.n247 VDD.t148 674.802
R2840 VDD.n41 VDD.n40 674.766
R2841 VDD.n97 VDD.n69 674.766
R2842 VDD.n418 VDD.t0 633.369
R2843 VDD.n16 VDD.t182 599.119
R2844 VDD.t144 VDD.n285 553.428
R2845 VDD.n286 VDD 432.123
R2846 VDD.t134 VDD.n313 420.43
R2847 VDD.n417 VDD.t91 420.25
R2848 VDD.n416 VDD.t129 420.25
R2849 VDD.n415 VDD.t66 420.25
R2850 VDD.n414 VDD.t158 420.25
R2851 VDD.n413 VDD.t174 420.25
R2852 VDD.n412 VDD.t64 420.25
R2853 VDD.n411 VDD.t136 420.25
R2854 VDD.n410 VDD.t221 420.25
R2855 VDD.n409 VDD.t202 420.25
R2856 VDD.n41 VDD.t81 414.33
R2857 VDD.n97 VDD.t166 414.33
R2858 VDD.t4 VDD 411.372
R2859 VDD VDD.t72 369.938
R2860 VDD VDD.t138 369.938
R2861 VDD VDD.t146 369.938
R2862 VDD VDD.t238 369.938
R2863 VDD VDD.t32 369.938
R2864 VDD VDD.t236 369.938
R2865 VDD VDD.t212 369.938
R2866 VDD VDD.t14 369.938
R2867 VDD VDD.t20 369.938
R2868 VDD VDD.t95 369.938
R2869 VDD VDD.t204 366.978
R2870 VDD.t102 VDD 366.978
R2871 VDD VDD.t34 361.06
R2872 VDD VDD.t200 361.06
R2873 VDD VDD.t194 361.06
R2874 VDD VDD.t44 361.06
R2875 VDD VDD.t76 361.06
R2876 VDD VDD.t176 361.06
R2877 VDD VDD.t87 361.06
R2878 VDD VDD.t168 361.06
R2879 VDD VDD.t234 361.06
R2880 VDD VDD.t127 361.06
R2881 VDD.t121 VDD 361.06
R2882 VDD.n291 VDD.t141 340.301
R2883 VDD.n294 VDD.t49 340.301
R2884 VDD.n316 VDD.t119 336.416
R2885 VDD.n319 VDD.n301 320.976
R2886 VDD.n334 VDD.n293 320.976
R2887 VDD.n339 VDD.n338 320.976
R2888 VDD.n224 VDD.n223 318.305
R2889 VDD.n326 VDD.n297 318.305
R2890 VDD.n380 VDD.n379 318.303
R2891 VDD VDD.t144 313.707
R2892 VDD.n372 VDD.n231 313.575
R2893 VDD.n96 VDD 276.123
R2894 VDD.n98 VDD 276.123
R2895 VDD.n68 VDD 276.123
R2896 VDD.n42 VDD 276.123
R2897 VDD VDD.n96 270.356
R2898 VDD.n96 VDD.n95 267.296
R2899 VDD.n99 VDD.n98 267.296
R2900 VDD.n68 VDD.n67 267.296
R2901 VDD.n43 VDD.n42 267.296
R2902 VDD.n402 VDD.t96 255.905
R2903 VDD.n112 VDD.t203 255.905
R2904 VDD.n215 VDD.t21 255.905
R2905 VDD.n116 VDD.t222 255.905
R2906 VDD.n206 VDD.t15 255.905
R2907 VDD.n120 VDD.t137 255.905
R2908 VDD.n197 VDD.t213 255.905
R2909 VDD.n124 VDD.t65 255.905
R2910 VDD.n188 VDD.t237 255.905
R2911 VDD.n128 VDD.t175 255.905
R2912 VDD.n179 VDD.t33 255.905
R2913 VDD.n132 VDD.t159 255.905
R2914 VDD.n170 VDD.t239 255.905
R2915 VDD.n136 VDD.t67 255.905
R2916 VDD.n161 VDD.t147 255.905
R2917 VDD.n140 VDD.t130 255.905
R2918 VDD.n152 VDD.t139 255.905
R2919 VDD.n144 VDD.t92 255.905
R2920 VDD.n424 VDD.t73 255.905
R2921 VDD.n3 VDD.t1 255.905
R2922 VDD.n378 VDD.t199 255.905
R2923 VDD.n279 VDD.t145 255.905
R2924 VDD.n308 VDD.t170 255.905
R2925 VDD.n225 VDD.t53 255.904
R2926 VDD.n308 VDD.t135 255.904
R2927 VDD.n398 VDD.t105 252.95
R2928 VDD.n403 VDD.t94 252.95
R2929 VDD.n113 VDD.t113 252.95
R2930 VDD.n214 VDD.t47 252.95
R2931 VDD.n208 VDD.t151 252.95
R2932 VDD.n205 VDD.t37 252.95
R2933 VDD.n199 VDD.t11 252.95
R2934 VDD.n196 VDD.t69 252.95
R2935 VDD.n190 VDD.t71 252.95
R2936 VDD.n187 VDD.t209 252.95
R2937 VDD.n181 VDD.t187 252.95
R2938 VDD.n178 VDD.t161 252.95
R2939 VDD.n172 VDD.t79 252.95
R2940 VDD.n169 VDD.t25 252.95
R2941 VDD.n163 VDD.t117 252.95
R2942 VDD.n160 VDD.t55 252.95
R2943 VDD.n154 VDD.t27 252.95
R2944 VDD.n151 VDD.t29 252.95
R2945 VDD.n145 VDD.t75 252.95
R2946 VDD.n423 VDD.t3 252.95
R2947 VDD.n299 VDD.t98 250.722
R2948 VDD.n376 VDD.t7 249.901
R2949 VDD.n370 VDD.t126 249.52
R2950 VDD.n294 VDD.t84 249.52
R2951 VDD.n384 VDD.t224 249.387
R2952 VDD.n234 VDD.t39 249.363
R2953 VDD.n366 VDD.t99 249.363
R2954 VDD.n267 VDD.t122 249.363
R2955 VDD.n272 VDD.t103 249.363
R2956 VDD.n256 VDD.t128 249.363
R2957 VDD.n243 VDD.t205 249.363
R2958 VDD.n5 VDD.t167 249.362
R2959 VDD.n79 VDD.t88 249.362
R2960 VDD.n84 VDD.t169 249.362
R2961 VDD.n89 VDD.t235 249.362
R2962 VDD.n46 VDD.t82 249.362
R2963 VDD.n51 VDD.t45 249.362
R2964 VDD.n56 VDD.t77 249.362
R2965 VDD.n61 VDD.t177 249.362
R2966 VDD.n18 VDD.t183 249.362
R2967 VDD.n23 VDD.t35 249.362
R2968 VDD.n28 VDD.t201 249.362
R2969 VDD.n33 VDD.t195 249.362
R2970 VDD.n234 VDD.t133 249.362
R2971 VDD.n366 VDD.t41 249.362
R2972 VDD.n325 VDD.t231 249.362
R2973 VDD.n290 VDD.t185 249.062
R2974 VDD.n289 VDD.t107 249.062
R2975 VDD.n350 VDD.t230 248.929
R2976 VDD.t0 VDD.t2 248.599
R2977 VDD.t72 VDD.t74 248.599
R2978 VDD.t91 VDD.t28 248.599
R2979 VDD.t138 VDD.t26 248.599
R2980 VDD.t129 VDD.t54 248.599
R2981 VDD.t146 VDD.t116 248.599
R2982 VDD.t66 VDD.t24 248.599
R2983 VDD.t238 VDD.t78 248.599
R2984 VDD.t158 VDD.t160 248.599
R2985 VDD.t32 VDD.t186 248.599
R2986 VDD.t174 VDD.t208 248.599
R2987 VDD.t236 VDD.t70 248.599
R2988 VDD.t64 VDD.t68 248.599
R2989 VDD.t212 VDD.t10 248.599
R2990 VDD.t136 VDD.t36 248.599
R2991 VDD.t14 VDD.t150 248.599
R2992 VDD.t221 VDD.t46 248.599
R2993 VDD.t20 VDD.t112 248.599
R2994 VDD.t202 VDD.t93 248.599
R2995 VDD.t95 VDD.t104 248.599
R2996 VDD.t182 VDD.t50 248.599
R2997 VDD.t34 VDD.t110 248.599
R2998 VDD.t200 VDD.t196 248.599
R2999 VDD.t194 VDD.t108 248.599
R3000 VDD.t81 VDD.t219 248.599
R3001 VDD.t44 VDD.t164 248.599
R3002 VDD.t76 VDD.t178 248.599
R3003 VDD.t176 VDD.t58 248.599
R3004 VDD.t166 VDD.t56 248.599
R3005 VDD.t87 VDD.t156 248.599
R3006 VDD.t168 VDD.t180 248.599
R3007 VDD.t234 VDD.t154 248.599
R3008 VDD.t204 VDD.t225 248.599
R3009 VDD.t127 VDD.t16 248.599
R3010 VDD.t214 VDD.t102 248.599
R3011 VDD.t142 VDD.t121 248.599
R3012 VDD.n359 VDD.t218 247.394
R3013 VDD.n364 VDD.t120 247.394
R3014 VDD.n268 VDD.t215 247.394
R3015 VDD.n240 VDD.t17 247.394
R3016 VDD.n255 VDD.t226 247.394
R3017 VDD.n290 VDD.t9 247.394
R3018 VDD.n346 VDD.t173 247.394
R3019 VDD.n289 VDD.t132 247.394
R3020 VDD.n78 VDD.t57 247.394
R3021 VDD.n83 VDD.t157 247.394
R3022 VDD.n88 VDD.t181 247.394
R3023 VDD.n70 VDD.t155 247.394
R3024 VDD.n50 VDD.t220 247.394
R3025 VDD.n55 VDD.t165 247.394
R3026 VDD.n60 VDD.t179 247.394
R3027 VDD.n6 VDD.t59 247.394
R3028 VDD.n22 VDD.t51 247.394
R3029 VDD.n27 VDD.t111 247.394
R3030 VDD.n32 VDD.t197 247.394
R3031 VDD.n11 VDD.t109 247.394
R3032 VDD.n359 VDD.t191 247.394
R3033 VDD.n364 VDD.t63 247.394
R3034 VDD.n370 VDD.t189 247.394
R3035 VDD.n327 VDD.t13 247.394
R3036 VDD.n238 VDD.t143 247.393
R3037 VDD.n332 VDD.t153 245.178
R3038 VDD.n345 VDD.t101 245.178
R3039 VDD.n324 VDD.t217 245.178
R3040 VDD.n229 VDD.t43 245.178
R3041 VDD.n277 VDD.t5 243.512
R3042 VDD.n248 VDD.t149 243.512
R3043 VDD.t40 VDD.n236 234.982
R3044 VDD.n352 VDD 230.766
R3045 VDD VDD.n417 221.964
R3046 VDD VDD.n416 221.964
R3047 VDD VDD.n415 221.964
R3048 VDD VDD.n414 221.964
R3049 VDD VDD.n413 221.964
R3050 VDD VDD.n412 221.964
R3051 VDD VDD.n411 221.964
R3052 VDD VDD.n410 221.964
R3053 VDD VDD.n409 221.964
R3054 VDD.n40 VDD 219.004
R3055 VDD.n69 VDD 219.004
R3056 VDD.n285 VDD 219.004
R3057 VDD.t60 VDD 216.519
R3058 VDD.n384 VDD.n227 213.119
R3059 VDD.n317 VDD.n302 213.119
R3060 VDD.n351 VDD.n350 213.119
R3061 VDD.n409 VDD.n408 213.119
R3062 VDD.n410 VDD.n111 213.119
R3063 VDD.n411 VDD.n110 213.119
R3064 VDD.n412 VDD.n109 213.119
R3065 VDD.n413 VDD.n108 213.119
R3066 VDD.n414 VDD.n107 213.119
R3067 VDD.n415 VDD.n106 213.119
R3068 VDD.n416 VDD.n105 213.119
R3069 VDD.n417 VDD.n104 213.119
R3070 VDD.n285 VDD.n284 213.119
R3071 VDD.n331 VDD.n295 213.119
R3072 VDD.t148 VDD.t80 213.084
R3073 VDD.t171 VDD.t4 213.084
R3074 VDD.n315 VDD.n314 209.368
R3075 VDD.t232 VDD 208.127
R3076 VDD.t50 VDD 207.166
R3077 VDD.t110 VDD 207.166
R3078 VDD.t196 VDD 207.166
R3079 VDD.t108 VDD 207.166
R3080 VDD.t219 VDD 207.166
R3081 VDD.t164 VDD 207.166
R3082 VDD.t178 VDD 207.166
R3083 VDD.t58 VDD 207.166
R3084 VDD.t56 VDD 207.166
R3085 VDD.t156 VDD 207.166
R3086 VDD.t180 VDD 207.166
R3087 VDD.t154 VDD 207.166
R3088 VDD.t225 VDD 207.166
R3089 VDD.t16 VDD 207.166
R3090 VDD VDD.t214 207.166
R3091 VDD VDD.t142 207.166
R3092 VDD VDD.t162 206.45
R3093 VDD.t38 VDD 204.77
R3094 VDD.t2 VDD 198.287
R3095 VDD.t74 VDD 198.287
R3096 VDD.t28 VDD 198.287
R3097 VDD.t26 VDD 198.287
R3098 VDD.t54 VDD 198.287
R3099 VDD.t116 VDD 198.287
R3100 VDD.t24 VDD 198.287
R3101 VDD.t78 VDD 198.287
R3102 VDD.t160 VDD 198.287
R3103 VDD.t186 VDD 198.287
R3104 VDD.t208 VDD 198.287
R3105 VDD.t70 VDD 198.287
R3106 VDD.t68 VDD 198.287
R3107 VDD.t10 VDD 198.287
R3108 VDD.t36 VDD 198.287
R3109 VDD.t150 VDD 198.287
R3110 VDD.t46 VDD 198.287
R3111 VDD.t112 VDD 198.287
R3112 VDD.t93 VDD 198.287
R3113 VDD.t104 VDD 198.287
R3114 VDD.n237 VDD 197.325
R3115 VDD.t80 VDD 189.409
R3116 VDD VDD.t171 189.409
R3117 VDD.n40 VDD.n39 184.788
R3118 VDD VDD.t134 177.916
R3119 VDD.t42 VDD.t123 154.417
R3120 VDD.t62 VDD.t40 140.989
R3121 VDD.t190 VDD.t38 140.989
R3122 VDD.t114 VDD.t206 140.989
R3123 VDD.t162 VDD.t12 140.989
R3124 VDD.t172 VDD.t229 140.989
R3125 VDD.t188 VDD.t227 134.276
R3126 VDD.t22 VDD.t152 134.276
R3127 VDD.t192 VDD.t8 134.276
R3128 VDD.t100 VDD.t30 134.276
R3129 VDD.t131 VDD.t85 134.276
R3130 VDD.n314 VDD 125.883
R3131 VDD.n236 VDD 124.206
R3132 VDD.n351 VDD 124.206
R3133 VDD VDD.t62 117.492
R3134 VDD VDD.t190 117.492
R3135 VDD VDD.t6 107.421
R3136 VDD VDD.t125 107.421
R3137 VDD.t216 VDD 107.421
R3138 VDD.t83 VDD 107.421
R3139 VDD.t184 VDD 107.421
R3140 VDD VDD.t106 107.421
R3141 VDD.n236 VDD.n232 106.559
R3142 VDD.n302 VDD.t114 100.707
R3143 VDD.n295 VDD.t22 100.707
R3144 VDD.t18 VDD 97.3503
R3145 VDD VDD.t89 95.6719
R3146 VDD VDD.t210 95.6719
R3147 VDD.n314 VDD.t118 93.9934
R3148 VDD VDD.t140 90.6365
R3149 VDD.t89 VDD.t52 82.2443
R3150 VDD.t210 VDD.t198 82.2443
R3151 VDD.n227 VDD.t223 80.5659
R3152 VDD.t229 VDD.n351 80.5659
R3153 VDD.t52 VDD.t60 78.8874
R3154 VDD.t198 VDD.t232 78.8874
R3155 VDD.t206 VDD.t97 72.1736
R3156 VDD.t30 VDD 70.4952
R3157 VDD.t97 VDD.t216 68.8168
R3158 VDD VDD.t48 67.1383
R3159 VDD.t118 VDD.n302 60.4245
R3160 VDD.t48 VDD.n295 60.4245
R3161 VDD.t123 VDD 53.7107
R3162 VDD.n42 VDD.n41 51.3536
R3163 VDD.n69 VDD.n68 51.3536
R3164 VDD.n98 VDD.n97 51.3536
R3165 VDD.t223 VDD 45.3185
R3166 VDD.t6 VDD 45.3185
R3167 VDD.n395 VDD.n394 43.9358
R3168 VDD VDD.t83 43.6401
R3169 VDD.n231 VDD.t124 38.4155
R3170 VDD.n379 VDD.t233 38.4155
R3171 VDD.n223 VDD.t61 38.4155
R3172 VDD.n297 VDD.t163 38.4155
R3173 VDD.n394 VDD.n222 34.6358
R3174 VDD.n390 VDD.n222 34.6358
R3175 VDD.n390 VDD.n389 34.6358
R3176 VDD.n273 VDD.n261 34.6358
R3177 VDD.n280 VDD.n239 34.6358
R3178 VDD.n250 VDD.n249 34.6358
R3179 VDD.n309 VDD.n306 34.6358
R3180 VDD.n315 VDD.n304 34.6358
R3181 VDD.n372 VDD.n371 33.1299
R3182 VDD.n335 VDD.n334 30.8711
R3183 VDD.n341 VDD.n339 30.8711
R3184 VDD.n320 VDD.n319 30.8711
R3185 VDD.n17 VDD.n16 29.8521
R3186 VDD.n39 VDD.n38 29.8521
R3187 VDD.n380 VDD.n226 27.4829
R3188 VDD.n389 VDD.n224 27.4829
R3189 VDD VDD.n227 26.8556
R3190 VDD.t140 VDD.t172 26.8556
R3191 VDD.n231 VDD.t228 26.5955
R3192 VDD.n379 VDD.t211 26.5955
R3193 VDD.n223 VDD.t90 26.5955
R3194 VDD.n293 VDD.t23 26.5955
R3195 VDD.n293 VDD.t193 26.5955
R3196 VDD.n338 VDD.t31 26.5955
R3197 VDD.n338 VDD.t86 26.5955
R3198 VDD.n297 VDD.t19 26.5955
R3199 VDD.n301 VDD.t115 26.5955
R3200 VDD.n301 VDD.t207 26.5955
R3201 VDD.n74 VDD.n5 25.977
R3202 VDD.n79 VDD.n73 25.977
R3203 VDD.n84 VDD.n72 25.977
R3204 VDD.n90 VDD.n89 25.977
R3205 VDD.n46 VDD.n10 25.977
R3206 VDD.n51 VDD.n9 25.977
R3207 VDD.n56 VDD.n8 25.977
R3208 VDD.n62 VDD.n61 25.977
R3209 VDD.n18 VDD.n15 25.977
R3210 VDD.n23 VDD.n14 25.977
R3211 VDD.n28 VDD.n13 25.977
R3212 VDD.n34 VDD.n33 25.977
R3213 VDD.n360 VDD.n234 25.977
R3214 VDD.n366 VDD.n365 25.977
R3215 VDD.n377 VDD.n376 25.977
R3216 VDD.n267 VDD.n263 25.977
R3217 VDD.n272 VDD.n262 25.977
R3218 VDD.n257 VDD.n256 25.977
R3219 VDD.n254 VDD.n243 25.977
R3220 VDD.n402 VDD.n220 25.224
R3221 VDD.n398 VDD.n220 25.224
R3222 VDD.n404 VDD.n112 25.224
R3223 VDD.n404 VDD.n403 25.224
R3224 VDD.n216 VDD.n215 25.224
R3225 VDD.n216 VDD.n113 25.224
R3226 VDD.n213 VDD.n116 25.224
R3227 VDD.n214 VDD.n213 25.224
R3228 VDD.n207 VDD.n206 25.224
R3229 VDD.n208 VDD.n207 25.224
R3230 VDD.n204 VDD.n120 25.224
R3231 VDD.n205 VDD.n204 25.224
R3232 VDD.n198 VDD.n197 25.224
R3233 VDD.n199 VDD.n198 25.224
R3234 VDD.n195 VDD.n124 25.224
R3235 VDD.n196 VDD.n195 25.224
R3236 VDD.n189 VDD.n188 25.224
R3237 VDD.n190 VDD.n189 25.224
R3238 VDD.n186 VDD.n128 25.224
R3239 VDD.n187 VDD.n186 25.224
R3240 VDD.n180 VDD.n179 25.224
R3241 VDD.n181 VDD.n180 25.224
R3242 VDD.n177 VDD.n132 25.224
R3243 VDD.n178 VDD.n177 25.224
R3244 VDD.n171 VDD.n170 25.224
R3245 VDD.n172 VDD.n171 25.224
R3246 VDD.n168 VDD.n136 25.224
R3247 VDD.n169 VDD.n168 25.224
R3248 VDD.n162 VDD.n161 25.224
R3249 VDD.n163 VDD.n162 25.224
R3250 VDD.n159 VDD.n140 25.224
R3251 VDD.n160 VDD.n159 25.224
R3252 VDD.n153 VDD.n152 25.224
R3253 VDD.n154 VDD.n153 25.224
R3254 VDD.n150 VDD.n144 25.224
R3255 VDD.n151 VDD.n150 25.224
R3256 VDD.n424 VDD.n2 25.224
R3257 VDD.n145 VDD.n2 25.224
R3258 VDD.n422 VDD.n3 25.224
R3259 VDD.n423 VDD.n422 25.224
R3260 VDD.n95 VDD.n94 25.1591
R3261 VDD.n100 VDD.n99 25.1591
R3262 VDD.n67 VDD.n66 25.1591
R3263 VDD.n45 VDD.n43 25.1591
R3264 VDD.n78 VDD.n74 24.4711
R3265 VDD.n83 VDD.n73 24.4711
R3266 VDD.n88 VDD.n72 24.4711
R3267 VDD.n90 VDD.n70 24.4711
R3268 VDD.n50 VDD.n10 24.4711
R3269 VDD.n55 VDD.n9 24.4711
R3270 VDD.n60 VDD.n8 24.4711
R3271 VDD.n62 VDD.n6 24.4711
R3272 VDD.n22 VDD.n15 24.4711
R3273 VDD.n27 VDD.n14 24.4711
R3274 VDD.n32 VDD.n13 24.4711
R3275 VDD.n34 VDD.n11 24.4711
R3276 VDD.n360 VDD.n359 24.4711
R3277 VDD.n365 VDD.n364 24.4711
R3278 VDD.n371 VDD.n370 24.4711
R3279 VDD.n263 VDD.n238 24.4711
R3280 VDD.n268 VDD.n262 24.4711
R3281 VDD.n278 VDD.n277 24.4711
R3282 VDD.n257 VDD.n240 24.4711
R3283 VDD.n255 VDD.n254 24.4711
R3284 VDD.n335 VDD.n290 24.4711
R3285 VDD.n341 VDD.n289 24.4711
R3286 VDD.n384 VDD.n226 23.7181
R3287 VDD.n385 VDD.n384 23.7181
R3288 VDD.n273 VDD.n272 23.7181
R3289 VDD.n284 VDD.n239 23.7181
R3290 VDD.n250 VDD.n243 23.7181
R3291 VDD.n318 VDD.n317 23.7181
R3292 VDD.n313 VDD.n306 23.7181
R3293 VDD.n376 VDD.n229 22.9652
R3294 VDD.n332 VDD.n331 22.5887
R3295 VDD.n346 VDD.n345 22.5887
R3296 VDD.n325 VDD.n324 22.5887
R3297 VDD.n317 VDD.n316 22.5887
R3298 VDD.n403 VDD.n402 20.3299
R3299 VDD.n215 VDD.n214 20.3299
R3300 VDD.n206 VDD.n205 20.3299
R3301 VDD.n197 VDD.n196 20.3299
R3302 VDD.n188 VDD.n187 20.3299
R3303 VDD.n179 VDD.n178 20.3299
R3304 VDD.n170 VDD.n169 20.3299
R3305 VDD.n161 VDD.n160 20.3299
R3306 VDD.n152 VDD.n151 20.3299
R3307 VDD.n424 VDD.n423 20.3299
R3308 VDD.t12 VDD.t18 20.1418
R3309 VDD.n277 VDD.n261 19.9534
R3310 VDD.n249 VDD.n248 19.9534
R3311 VDD.n326 VDD.n325 18.824
R3312 VDD.n320 VDD.n299 18.4476
R3313 VDD.n356 VDD.n237 18.084
R3314 VDD.n408 VDD.n112 17.3181
R3315 VDD.n116 VDD.n111 17.3181
R3316 VDD.n120 VDD.n110 17.3181
R3317 VDD.n124 VDD.n109 17.3181
R3318 VDD.n128 VDD.n108 17.3181
R3319 VDD.n132 VDD.n107 17.3181
R3320 VDD.n136 VDD.n106 17.3181
R3321 VDD.n140 VDD.n105 17.3181
R3322 VDD.n144 VDD.n104 17.3181
R3323 VDD.n418 VDD.n3 17.3181
R3324 VDD.n323 VDD.n299 16.1887
R3325 VDD.n408 VDD.n113 15.8123
R3326 VDD.n208 VDD.n111 15.8123
R3327 VDD.n199 VDD.n110 15.8123
R3328 VDD.n190 VDD.n109 15.8123
R3329 VDD.n181 VDD.n108 15.8123
R3330 VDD.n172 VDD.n107 15.8123
R3331 VDD.n163 VDD.n106 15.8123
R3332 VDD.n154 VDD.n105 15.8123
R3333 VDD.n145 VDD.n104 15.8123
R3334 VDD.n350 VDD.n291 14.3064
R3335 VDD.n327 VDD.n294 14.3064
R3336 VDD.n327 VDD.n326 14.3064
R3337 VDD.n248 VDD.n247 13.5534
R3338 VDD.n103 VDD.n4 12.8047
R3339 VDD.n100 VDD.n5 12.8005
R3340 VDD.n79 VDD.n78 12.8005
R3341 VDD.n84 VDD.n83 12.8005
R3342 VDD.n89 VDD.n88 12.8005
R3343 VDD.n94 VDD.n70 12.8005
R3344 VDD.n46 VDD.n45 12.8005
R3345 VDD.n51 VDD.n50 12.8005
R3346 VDD.n56 VDD.n55 12.8005
R3347 VDD.n61 VDD.n60 12.8005
R3348 VDD.n66 VDD.n6 12.8005
R3349 VDD.n18 VDD.n17 12.8005
R3350 VDD.n23 VDD.n22 12.8005
R3351 VDD.n28 VDD.n27 12.8005
R3352 VDD.n33 VDD.n32 12.8005
R3353 VDD.n38 VDD.n11 12.8005
R3354 VDD.n359 VDD.n358 12.8005
R3355 VDD.n364 VDD.n234 12.8005
R3356 VDD.n366 VDD.n232 12.8005
R3357 VDD.n370 VDD.n232 12.8005
R3358 VDD.n286 VDD.n238 12.8005
R3359 VDD.n268 VDD.n267 12.8005
R3360 VDD.n284 VDD.n240 12.8005
R3361 VDD.n256 VDD.n255 12.8005
R3362 VDD.n350 VDD.n290 12.8005
R3363 VDD.n346 VDD.n291 12.8005
R3364 VDD.n352 VDD.n289 12.8005
R3365 VDD.n331 VDD.n294 12.0476
R3366 VDD.n103 VDD.n102 11.6828
R3367 VDD.n280 VDD.n279 10.5417
R3368 VDD.n309 VDD.n308 10.5417
R3369 VDD.n95 VDD 9.71084
R3370 VDD.n99 VDD 9.71084
R3371 VDD.n67 VDD 9.71084
R3372 VDD.n43 VDD 9.71084
R3373 VDD.n17 VDD 9.32654
R3374 VDD.n38 VDD.n37 9.3005
R3375 VDD.n19 VDD.n18 9.3005
R3376 VDD.n20 VDD.n15 9.3005
R3377 VDD.n22 VDD.n21 9.3005
R3378 VDD.n24 VDD.n23 9.3005
R3379 VDD.n25 VDD.n14 9.3005
R3380 VDD.n27 VDD.n26 9.3005
R3381 VDD.n29 VDD.n28 9.3005
R3382 VDD.n30 VDD.n13 9.3005
R3383 VDD.n32 VDD.n31 9.3005
R3384 VDD.n33 VDD.n12 9.3005
R3385 VDD.n35 VDD.n34 9.3005
R3386 VDD.n36 VDD.n11 9.3005
R3387 VDD.n66 VDD.n65 9.3005
R3388 VDD.n45 VDD.n44 9.3005
R3389 VDD.n47 VDD.n46 9.3005
R3390 VDD.n48 VDD.n10 9.3005
R3391 VDD.n50 VDD.n49 9.3005
R3392 VDD.n52 VDD.n51 9.3005
R3393 VDD.n53 VDD.n9 9.3005
R3394 VDD.n55 VDD.n54 9.3005
R3395 VDD.n57 VDD.n56 9.3005
R3396 VDD.n58 VDD.n8 9.3005
R3397 VDD.n60 VDD.n59 9.3005
R3398 VDD.n61 VDD.n7 9.3005
R3399 VDD.n63 VDD.n62 9.3005
R3400 VDD.n64 VDD.n6 9.3005
R3401 VDD.n94 VDD.n93 9.3005
R3402 VDD.n101 VDD.n100 9.3005
R3403 VDD.n75 VDD.n5 9.3005
R3404 VDD.n76 VDD.n74 9.3005
R3405 VDD.n78 VDD.n77 9.3005
R3406 VDD.n80 VDD.n79 9.3005
R3407 VDD.n81 VDD.n73 9.3005
R3408 VDD.n83 VDD.n82 9.3005
R3409 VDD.n85 VDD.n84 9.3005
R3410 VDD.n86 VDD.n72 9.3005
R3411 VDD.n88 VDD.n87 9.3005
R3412 VDD.n89 VDD.n71 9.3005
R3413 VDD.n91 VDD.n90 9.3005
R3414 VDD.n92 VDD.n70 9.3005
R3415 VDD.n247 VDD.n246 9.3005
R3416 VDD.n248 VDD.n245 9.3005
R3417 VDD.n249 VDD.n244 9.3005
R3418 VDD.n251 VDD.n250 9.3005
R3419 VDD.n252 VDD.n243 9.3005
R3420 VDD.n254 VDD.n253 9.3005
R3421 VDD.n255 VDD.n242 9.3005
R3422 VDD.n256 VDD.n241 9.3005
R3423 VDD.n258 VDD.n257 9.3005
R3424 VDD.n259 VDD.n240 9.3005
R3425 VDD.n284 VDD.n283 9.3005
R3426 VDD.n282 VDD.n239 9.3005
R3427 VDD.n281 VDD.n280 9.3005
R3428 VDD.n278 VDD.n260 9.3005
R3429 VDD.n277 VDD.n276 9.3005
R3430 VDD.n275 VDD.n261 9.3005
R3431 VDD.n274 VDD.n273 9.3005
R3432 VDD.n272 VDD.n271 9.3005
R3433 VDD.n270 VDD.n262 9.3005
R3434 VDD.n269 VDD.n268 9.3005
R3435 VDD.n267 VDD.n266 9.3005
R3436 VDD.n265 VDD.n263 9.3005
R3437 VDD.n264 VDD.n238 9.3005
R3438 VDD.n287 VDD.n286 9.3005
R3439 VDD.n353 VDD.n352 9.3005
R3440 VDD.n313 VDD.n312 9.3005
R3441 VDD.n311 VDD.n306 9.3005
R3442 VDD.n310 VDD.n309 9.3005
R3443 VDD.n307 VDD.n304 9.3005
R3444 VDD.n315 VDD.n305 9.3005
R3445 VDD.n317 VDD.n303 9.3005
R3446 VDD.n318 VDD.n300 9.3005
R3447 VDD.n321 VDD.n320 9.3005
R3448 VDD.n323 VDD.n322 9.3005
R3449 VDD.n325 VDD.n298 9.3005
R3450 VDD.n326 VDD.n296 9.3005
R3451 VDD.n328 VDD.n327 9.3005
R3452 VDD.n329 VDD.n294 9.3005
R3453 VDD.n331 VDD.n330 9.3005
R3454 VDD.n333 VDD.n292 9.3005
R3455 VDD.n336 VDD.n335 9.3005
R3456 VDD.n337 VDD.n290 9.3005
R3457 VDD.n350 VDD.n349 9.3005
R3458 VDD.n348 VDD.n291 9.3005
R3459 VDD.n347 VDD.n346 9.3005
R3460 VDD.n344 VDD.n343 9.3005
R3461 VDD.n342 VDD.n341 9.3005
R3462 VDD.n340 VDD.n289 9.3005
R3463 VDD.n394 VDD.n393 9.3005
R3464 VDD.n392 VDD.n222 9.3005
R3465 VDD.n391 VDD.n390 9.3005
R3466 VDD.n389 VDD.n388 9.3005
R3467 VDD.n387 VDD.n224 9.3005
R3468 VDD.n386 VDD.n385 9.3005
R3469 VDD.n384 VDD.n383 9.3005
R3470 VDD.n382 VDD.n226 9.3005
R3471 VDD.n381 VDD.n380 9.3005
R3472 VDD.n377 VDD.n228 9.3005
R3473 VDD.n376 VDD.n375 9.3005
R3474 VDD.n374 VDD.n373 9.3005
R3475 VDD.n371 VDD.n230 9.3005
R3476 VDD.n370 VDD.n369 9.3005
R3477 VDD.n368 VDD.n232 9.3005
R3478 VDD.n367 VDD.n366 9.3005
R3479 VDD.n365 VDD.n233 9.3005
R3480 VDD.n364 VDD.n363 9.3005
R3481 VDD.n362 VDD.n234 9.3005
R3482 VDD.n361 VDD.n360 9.3005
R3483 VDD.n359 VDD.n235 9.3005
R3484 VDD.n358 VDD.n357 9.3005
R3485 VDD.n419 VDD.n418 9.3005
R3486 VDD.n420 VDD.n3 9.3005
R3487 VDD.n422 VDD.n421 9.3005
R3488 VDD.n423 VDD.n0 9.3005
R3489 VDD.n425 VDD.n424 9.3005
R3490 VDD.n2 VDD.n1 9.3005
R3491 VDD.n146 VDD.n145 9.3005
R3492 VDD.n147 VDD.n104 9.3005
R3493 VDD.n148 VDD.n144 9.3005
R3494 VDD.n150 VDD.n149 9.3005
R3495 VDD.n151 VDD.n143 9.3005
R3496 VDD.n152 VDD.n142 9.3005
R3497 VDD.n153 VDD.n141 9.3005
R3498 VDD.n155 VDD.n154 9.3005
R3499 VDD.n156 VDD.n105 9.3005
R3500 VDD.n157 VDD.n140 9.3005
R3501 VDD.n159 VDD.n158 9.3005
R3502 VDD.n160 VDD.n139 9.3005
R3503 VDD.n161 VDD.n138 9.3005
R3504 VDD.n162 VDD.n137 9.3005
R3505 VDD.n164 VDD.n163 9.3005
R3506 VDD.n165 VDD.n106 9.3005
R3507 VDD.n166 VDD.n136 9.3005
R3508 VDD.n168 VDD.n167 9.3005
R3509 VDD.n169 VDD.n135 9.3005
R3510 VDD.n170 VDD.n134 9.3005
R3511 VDD.n171 VDD.n133 9.3005
R3512 VDD.n173 VDD.n172 9.3005
R3513 VDD.n174 VDD.n107 9.3005
R3514 VDD.n175 VDD.n132 9.3005
R3515 VDD.n177 VDD.n176 9.3005
R3516 VDD.n178 VDD.n131 9.3005
R3517 VDD.n179 VDD.n130 9.3005
R3518 VDD.n180 VDD.n129 9.3005
R3519 VDD.n182 VDD.n181 9.3005
R3520 VDD.n183 VDD.n108 9.3005
R3521 VDD.n184 VDD.n128 9.3005
R3522 VDD.n186 VDD.n185 9.3005
R3523 VDD.n187 VDD.n127 9.3005
R3524 VDD.n188 VDD.n126 9.3005
R3525 VDD.n189 VDD.n125 9.3005
R3526 VDD.n191 VDD.n190 9.3005
R3527 VDD.n192 VDD.n109 9.3005
R3528 VDD.n193 VDD.n124 9.3005
R3529 VDD.n195 VDD.n194 9.3005
R3530 VDD.n196 VDD.n123 9.3005
R3531 VDD.n197 VDD.n122 9.3005
R3532 VDD.n198 VDD.n121 9.3005
R3533 VDD.n200 VDD.n199 9.3005
R3534 VDD.n201 VDD.n110 9.3005
R3535 VDD.n202 VDD.n120 9.3005
R3536 VDD.n204 VDD.n203 9.3005
R3537 VDD.n205 VDD.n119 9.3005
R3538 VDD.n206 VDD.n118 9.3005
R3539 VDD.n207 VDD.n117 9.3005
R3540 VDD.n209 VDD.n208 9.3005
R3541 VDD.n210 VDD.n111 9.3005
R3542 VDD.n211 VDD.n116 9.3005
R3543 VDD.n213 VDD.n212 9.3005
R3544 VDD.n214 VDD.n115 9.3005
R3545 VDD.n215 VDD.n114 9.3005
R3546 VDD.n217 VDD.n216 9.3005
R3547 VDD.n218 VDD.n113 9.3005
R3548 VDD.n408 VDD.n407 9.3005
R3549 VDD.n406 VDD.n112 9.3005
R3550 VDD.n405 VDD.n404 9.3005
R3551 VDD.n403 VDD.n219 9.3005
R3552 VDD.n402 VDD.n401 9.3005
R3553 VDD.n400 VDD.n220 9.3005
R3554 VDD.n399 VDD.n398 9.3005
R3555 VDD.n378 VDD.n377 8.28285
R3556 VDD.n385 VDD.n225 8.28285
R3557 VDD.n279 VDD.n278 8.28285
R3558 VDD.n308 VDD.n304 8.28285
R3559 VDD.t227 VDD.t42 6.71428
R3560 VDD.t125 VDD.t188 6.71428
R3561 VDD.t152 VDD.t192 6.71428
R3562 VDD.t8 VDD.t184 6.71428
R3563 VDD.t85 VDD.t100 6.71428
R3564 VDD.t106 VDD.t131 6.71428
R3565 VDD.n16 VDD 4.84842
R3566 VDD.n39 VDD 4.84842
R3567 VDD.n355 VDD 4.63938
R3568 VDD.n397 VDD 4.08544
R3569 VDD.n246 VDD.n221 3.76683
R3570 VDD.n334 VDD.n333 3.76521
R3571 VDD.n344 VDD.n339 3.76521
R3572 VDD.n319 VDD.n318 3.76521
R3573 VDD.n358 VDD.n237 3.58719
R3574 VDD.n288 VDD 3.09034
R3575 VDD.n354 VDD 3.09034
R3576 VDD VDD.n355 3.09034
R3577 VDD VDD.n397 3.03019
R3578 VDD.n312 VDD.n221 2.89503
R3579 VDD.n396 VDD.n395 2.89503
R3580 VDD.n419 VDD.n103 2.77316
R3581 VDD.n397 VDD 2.27784
R3582 VDD.n373 VDD.n372 1.50638
R3583 VDD.n373 VDD.n229 1.12991
R3584 VDD.n333 VDD.n332 1.12991
R3585 VDD.n345 VDD.n344 1.12991
R3586 VDD.n324 VDD.n323 1.12991
R3587 VDD.n316 VDD.n315 1.12991
R3588 VDD.n396 VDD.n221 0.872295
R3589 VDD.n354 VDD.n288 0.872295
R3590 VDD.n355 VDD 0.462038
R3591 VDD VDD.n354 0.410756
R3592 VDD.n380 VDD.n378 0.376971
R3593 VDD.n225 VDD.n224 0.376971
R3594 VDD VDD.n396 0.252103
R3595 VDD.n20 VDD.n19 0.120292
R3596 VDD.n21 VDD.n20 0.120292
R3597 VDD.n25 VDD.n24 0.120292
R3598 VDD.n26 VDD.n25 0.120292
R3599 VDD.n30 VDD.n29 0.120292
R3600 VDD.n31 VDD.n30 0.120292
R3601 VDD.n35 VDD.n12 0.120292
R3602 VDD.n36 VDD.n35 0.120292
R3603 VDD.n48 VDD.n47 0.120292
R3604 VDD.n49 VDD.n48 0.120292
R3605 VDD.n53 VDD.n52 0.120292
R3606 VDD.n54 VDD.n53 0.120292
R3607 VDD.n58 VDD.n57 0.120292
R3608 VDD.n59 VDD.n58 0.120292
R3609 VDD.n63 VDD.n7 0.120292
R3610 VDD.n64 VDD.n63 0.120292
R3611 VDD.n76 VDD.n75 0.120292
R3612 VDD.n77 VDD.n76 0.120292
R3613 VDD.n81 VDD.n80 0.120292
R3614 VDD.n82 VDD.n81 0.120292
R3615 VDD.n86 VDD.n85 0.120292
R3616 VDD.n87 VDD.n86 0.120292
R3617 VDD.n91 VDD.n71 0.120292
R3618 VDD.n92 VDD.n91 0.120292
R3619 VDD.n245 VDD.n244 0.120292
R3620 VDD.n251 VDD.n244 0.120292
R3621 VDD.n253 VDD.n252 0.120292
R3622 VDD.n253 VDD.n242 0.120292
R3623 VDD.n258 VDD.n241 0.120292
R3624 VDD.n259 VDD.n258 0.120292
R3625 VDD.n282 VDD.n281 0.120292
R3626 VDD.n281 VDD.n260 0.120292
R3627 VDD.n276 VDD.n275 0.120292
R3628 VDD.n275 VDD.n274 0.120292
R3629 VDD.n271 VDD.n270 0.120292
R3630 VDD.n270 VDD.n269 0.120292
R3631 VDD.n266 VDD.n265 0.120292
R3632 VDD.n265 VDD.n264 0.120292
R3633 VDD.n311 VDD.n310 0.120292
R3634 VDD.n310 VDD.n307 0.120292
R3635 VDD.n321 VDD.n300 0.120292
R3636 VDD.n322 VDD.n321 0.120292
R3637 VDD.n298 VDD.n296 0.120292
R3638 VDD.n328 VDD.n296 0.120292
R3639 VDD.n336 VDD.n292 0.120292
R3640 VDD.n337 VDD.n336 0.120292
R3641 VDD.n348 VDD.n347 0.120292
R3642 VDD.n343 VDD.n342 0.120292
R3643 VDD.n342 VDD.n340 0.120292
R3644 VDD.n393 VDD.n392 0.120292
R3645 VDD.n392 VDD.n391 0.120292
R3646 VDD.n388 VDD.n387 0.120292
R3647 VDD.n387 VDD.n386 0.120292
R3648 VDD.n382 VDD.n381 0.120292
R3649 VDD.n381 VDD.n228 0.120292
R3650 VDD.n374 VDD.n230 0.120292
R3651 VDD.n369 VDD.n230 0.120292
R3652 VDD.n367 VDD.n233 0.120292
R3653 VDD.n363 VDD.n233 0.120292
R3654 VDD.n362 VDD.n361 0.120292
R3655 VDD.n361 VDD.n235 0.120292
R3656 VDD.n44 VDD 0.11899
R3657 VDD VDD.n101 0.11899
R3658 VDD.n393 VDD 0.109875
R3659 VDD.n388 VDD 0.104667
R3660 VDD.n102 VDD 0.09425
R3661 VDD VDD.n4 0.078625
R3662 VDD.n421 VDD.n420 0.072375
R3663 VDD.n421 VDD.n0 0.072375
R3664 VDD.n425 VDD.n1 0.072375
R3665 VDD.n146 VDD.n1 0.072375
R3666 VDD.n149 VDD.n148 0.072375
R3667 VDD.n149 VDD.n143 0.072375
R3668 VDD.n142 VDD.n141 0.072375
R3669 VDD.n155 VDD.n141 0.072375
R3670 VDD.n158 VDD.n157 0.072375
R3671 VDD.n158 VDD.n139 0.072375
R3672 VDD.n138 VDD.n137 0.072375
R3673 VDD.n164 VDD.n137 0.072375
R3674 VDD.n167 VDD.n166 0.072375
R3675 VDD.n167 VDD.n135 0.072375
R3676 VDD.n134 VDD.n133 0.072375
R3677 VDD.n173 VDD.n133 0.072375
R3678 VDD.n176 VDD.n175 0.072375
R3679 VDD.n176 VDD.n131 0.072375
R3680 VDD.n130 VDD.n129 0.072375
R3681 VDD.n182 VDD.n129 0.072375
R3682 VDD.n185 VDD.n184 0.072375
R3683 VDD.n185 VDD.n127 0.072375
R3684 VDD.n126 VDD.n125 0.072375
R3685 VDD.n191 VDD.n125 0.072375
R3686 VDD.n194 VDD.n193 0.072375
R3687 VDD.n194 VDD.n123 0.072375
R3688 VDD.n122 VDD.n121 0.072375
R3689 VDD.n200 VDD.n121 0.072375
R3690 VDD.n203 VDD.n202 0.072375
R3691 VDD.n203 VDD.n119 0.072375
R3692 VDD.n118 VDD.n117 0.072375
R3693 VDD.n209 VDD.n117 0.072375
R3694 VDD.n212 VDD.n211 0.072375
R3695 VDD.n212 VDD.n115 0.072375
R3696 VDD.n217 VDD.n114 0.072375
R3697 VDD.n218 VDD.n217 0.072375
R3698 VDD.n406 VDD.n405 0.072375
R3699 VDD.n405 VDD.n219 0.072375
R3700 VDD.n401 VDD.n400 0.072375
R3701 VDD.n400 VDD.n399 0.072375
R3702 VDD.n19 VDD 0.0603958
R3703 VDD.n24 VDD 0.0603958
R3704 VDD.n29 VDD 0.0603958
R3705 VDD VDD.n12 0.0603958
R3706 VDD.n37 VDD 0.0603958
R3707 VDD.n47 VDD 0.0603958
R3708 VDD.n52 VDD 0.0603958
R3709 VDD.n57 VDD 0.0603958
R3710 VDD VDD.n7 0.0603958
R3711 VDD.n65 VDD 0.0603958
R3712 VDD.n75 VDD 0.0603958
R3713 VDD.n80 VDD 0.0603958
R3714 VDD.n85 VDD 0.0603958
R3715 VDD VDD.n71 0.0603958
R3716 VDD.n93 VDD 0.0603958
R3717 VDD VDD.n245 0.0603958
R3718 VDD.n252 VDD 0.0603958
R3719 VDD VDD.n241 0.0603958
R3720 VDD.n283 VDD 0.0603958
R3721 VDD VDD.n282 0.0603958
R3722 VDD.n276 VDD 0.0603958
R3723 VDD.n271 VDD 0.0603958
R3724 VDD.n266 VDD 0.0603958
R3725 VDD.n287 VDD 0.0603958
R3726 VDD VDD.n311 0.0603958
R3727 VDD VDD.n305 0.0603958
R3728 VDD VDD.n303 0.0603958
R3729 VDD VDD.n300 0.0603958
R3730 VDD VDD.n298 0.0603958
R3731 VDD.n329 VDD 0.0603958
R3732 VDD.n330 VDD 0.0603958
R3733 VDD VDD.n292 0.0603958
R3734 VDD.n349 VDD 0.0603958
R3735 VDD VDD.n348 0.0603958
R3736 VDD.n343 VDD 0.0603958
R3737 VDD.n353 VDD 0.0603958
R3738 VDD.n383 VDD 0.0603958
R3739 VDD VDD.n382 0.0603958
R3740 VDD.n375 VDD 0.0603958
R3741 VDD VDD.n374 0.0603958
R3742 VDD VDD.n368 0.0603958
R3743 VDD VDD.n367 0.0603958
R3744 VDD VDD.n362 0.0603958
R3745 VDD.n357 VDD 0.0603958
R3746 VDD VDD.n356 0.0603958
R3747 VDD VDD.n4 0.0408646
R3748 VDD.n283 VDD 0.0382604
R3749 VDD.n288 VDD 0.0365577
R3750 VDD.n420 VDD 0.0364375
R3751 VDD VDD.n425 0.0364375
R3752 VDD.n147 VDD 0.0364375
R3753 VDD.n148 VDD 0.0364375
R3754 VDD VDD.n142 0.0364375
R3755 VDD.n156 VDD 0.0364375
R3756 VDD.n157 VDD 0.0364375
R3757 VDD VDD.n138 0.0364375
R3758 VDD.n165 VDD 0.0364375
R3759 VDD.n166 VDD 0.0364375
R3760 VDD VDD.n134 0.0364375
R3761 VDD.n174 VDD 0.0364375
R3762 VDD.n175 VDD 0.0364375
R3763 VDD VDD.n130 0.0364375
R3764 VDD.n183 VDD 0.0364375
R3765 VDD.n184 VDD 0.0364375
R3766 VDD VDD.n126 0.0364375
R3767 VDD.n192 VDD 0.0364375
R3768 VDD.n193 VDD 0.0364375
R3769 VDD VDD.n122 0.0364375
R3770 VDD.n201 VDD 0.0364375
R3771 VDD.n202 VDD 0.0364375
R3772 VDD VDD.n118 0.0364375
R3773 VDD.n210 VDD 0.0364375
R3774 VDD.n211 VDD 0.0364375
R3775 VDD VDD.n114 0.0364375
R3776 VDD.n407 VDD 0.0364375
R3777 VDD VDD.n406 0.0364375
R3778 VDD.n401 VDD 0.0364375
R3779 VDD.n246 VDD 0.03175
R3780 VDD VDD.n287 0.03175
R3781 VDD.n312 VDD 0.03175
R3782 VDD.n305 VDD 0.03175
R3783 VDD.n303 VDD 0.03175
R3784 VDD.n330 VDD 0.03175
R3785 VDD.n349 VDD 0.03175
R3786 VDD VDD.n353 0.03175
R3787 VDD.n368 VDD 0.03175
R3788 VDD.n357 VDD 0.03175
R3789 VDD.n356 VDD 0.03175
R3790 VDD.n37 VDD 0.0265417
R3791 VDD.n44 VDD 0.0265417
R3792 VDD.n65 VDD 0.0265417
R3793 VDD.n101 VDD 0.0265417
R3794 VDD.n93 VDD 0.0265417
R3795 VDD.n102 VDD 0.0252396
R3796 VDD.n21 VDD 0.0239375
R3797 VDD.n26 VDD 0.0239375
R3798 VDD.n31 VDD 0.0239375
R3799 VDD VDD.n36 0.0239375
R3800 VDD.n49 VDD 0.0239375
R3801 VDD.n54 VDD 0.0239375
R3802 VDD.n59 VDD 0.0239375
R3803 VDD VDD.n64 0.0239375
R3804 VDD.n77 VDD 0.0239375
R3805 VDD.n82 VDD 0.0239375
R3806 VDD.n87 VDD 0.0239375
R3807 VDD VDD.n92 0.0239375
R3808 VDD.n242 VDD 0.0239375
R3809 VDD VDD.n259 0.0239375
R3810 VDD.n269 VDD 0.0239375
R3811 VDD.n264 VDD 0.0239375
R3812 VDD VDD.n328 0.0239375
R3813 VDD.n347 VDD 0.0239375
R3814 VDD.n363 VDD 0.0239375
R3815 VDD VDD.n235 0.0239375
R3816 VDD VDD.n260 0.0226354
R3817 VDD.n307 VDD 0.0226354
R3818 VDD.n386 VDD 0.0226354
R3819 VDD VDD.n228 0.0226354
R3820 VDD VDD.n251 0.0213333
R3821 VDD.n274 VDD 0.0213333
R3822 VDD.n322 VDD 0.0213333
R3823 VDD VDD.n329 0.0213333
R3824 VDD VDD.n337 0.0213333
R3825 VDD.n340 VDD 0.0213333
R3826 VDD.n383 VDD 0.0213333
R3827 VDD.n375 VDD 0.0213333
R3828 VDD.n369 VDD 0.0213333
R3829 VDD VDD.n419 0.01925
R3830 VDD VDD.n147 0.01925
R3831 VDD VDD.n156 0.01925
R3832 VDD VDD.n165 0.01925
R3833 VDD VDD.n174 0.01925
R3834 VDD VDD.n183 0.01925
R3835 VDD VDD.n192 0.01925
R3836 VDD VDD.n201 0.01925
R3837 VDD VDD.n210 0.01925
R3838 VDD.n407 VDD 0.01925
R3839 VDD.n391 VDD 0.016125
R3840 VDD VDD.n0 0.0137813
R3841 VDD VDD.n146 0.0137813
R3842 VDD.n143 VDD 0.0137813
R3843 VDD VDD.n155 0.0137813
R3844 VDD.n139 VDD 0.0137813
R3845 VDD VDD.n164 0.0137813
R3846 VDD.n135 VDD 0.0137813
R3847 VDD VDD.n173 0.0137813
R3848 VDD.n131 VDD 0.0137813
R3849 VDD VDD.n182 0.0137813
R3850 VDD.n127 VDD 0.0137813
R3851 VDD VDD.n191 0.0137813
R3852 VDD.n123 VDD 0.0137813
R3853 VDD VDD.n200 0.0137813
R3854 VDD.n119 VDD 0.0137813
R3855 VDD VDD.n209 0.0137813
R3856 VDD.n115 VDD 0.0137813
R3857 VDD VDD.n218 0.0137813
R3858 VDD VDD.n219 0.0137813
R3859 VDD.n399 VDD 0.0137813
R3860 VDD.n395 VDD 0.0109167
R3861 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t4 732.773
R3862 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t6 241.536
R3863 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t8 232.214
R3864 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t17 232.214
R3865 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t19 229.369
R3866 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t9 229.369
R3867 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t16 229.369
R3868 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t15 212.081
R3869 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t13 212.081
R3870 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 208.964
R3871 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 186.001
R3872 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t18 169.237
R3873 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t7 159.915
R3874 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t11 159.915
R3875 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t5 157.07
R3876 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t20 157.07
R3877 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t10 157.07
R3878 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 155.88
R3879 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 152.712
R3880 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 152.475
R3881 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 152
R3882 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 152
R3883 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 152
R3884 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t14 139.78
R3885 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t12 139.78
R3886 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 96.8352
R3887 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 61.346
R3888 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t3 26.5955
R3889 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t0 26.5955
R3890 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t2 24.9236
R3891 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t1 24.9236
R3892 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 23.417
R3893 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 21.3854
R3894 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 20.0025
R3895 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 18.2158
R3896 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 17.7529
R3897 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 12.5445
R3898 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 12.4213
R3899 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 11.7484
R3900 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 11.2645
R3901 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 10.9817
R3902 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 10.2234
R3903 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 9.77342
R3904 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 9.65467
R3905 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 9.30258
R3906 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 6.98232
R3907 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 6.1445
R3908 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 6.12758
R3909 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 5.92643
R3910 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 5.45235
R3911 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 5.21532
R3912 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 5.04425
R3913 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 4.8645
R3914 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 4.65505
R3915 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 3.0725
R3916 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 2.27147
R3917 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 2.27147
R3918 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 2.0485
R3919 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 1.55202
R3920 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 1.53956
R3921 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 1.42823
R3922 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 0.770031
R3923 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 0.623547
R3924 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.334484
R3925 a_20048_n709.t0 a_20048_n709.t1 114.052
R3926 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t4 732.702
R3927 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 208.964
R3928 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 96.8352
R3929 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 28.767
R3930 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t2 26.5955
R3931 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t0 26.5955
R3932 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t1 24.9236
R3933 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t3 24.9236
R3934 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 13.0565
R3935 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 11.2645
R3936 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 6.1445
R3937 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 4.65505
R3938 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 4.3525
R3939 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 2.0485
R3940 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 1.55202
R3941 a_17344_n1619.t0 a_17344_n1619.t1 114.052
R3942 dcell_lv_0.bb[8].n11 dcell_lv_0.bb[8].t10 230.363
R3943 dcell_lv_0.bb[8].n8 dcell_lv_0.bb[8].t13 230.155
R3944 dcell_lv_0.bb[8].n5 dcell_lv_0.bb[8].t11 229.369
R3945 dcell_lv_0.bb[8].n2 dcell_lv_0.bb[8].t9 212.081
R3946 dcell_lv_0.bb[8].n3 dcell_lv_0.bb[8].t5 212.081
R3947 dcell_lv_0.bb[8].n1 dcell_lv_0.bb[8].n0 208.965
R3948 dcell_lv_0.bb[8].n4 dcell_lv_0.bb[8].n3 186.001
R3949 dcell_lv_0.bb[8].n11 dcell_lv_0.bb[8].t7 158.064
R3950 dcell_lv_0.bb[8].n8 dcell_lv_0.bb[8].t12 157.856
R3951 dcell_lv_0.bb[8].n5 dcell_lv_0.bb[8].t6 157.07
R3952 dcell_lv_0.bb[8].n6 dcell_lv_0.bb[8].n5 152
R3953 dcell_lv_0.bb[8].n9 dcell_lv_0.bb[8].n8 152
R3954 dcell_lv_0.bb[8].n12 dcell_lv_0.bb[8].n11 152
R3955 dcell_lv_0.bb[8].n2 dcell_lv_0.bb[8].t8 139.78
R3956 dcell_lv_0.bb[8].n3 dcell_lv_0.bb[8].t4 139.78
R3957 dcell_lv_0.bb[8] dcell_lv_0.bb[8].n17 96.8352
R3958 dcell_lv_0.bb[8].n3 dcell_lv_0.bb[8].n2 61.346
R3959 dcell_lv_0.bb[8].n10 dcell_lv_0.bb[8].n9 36.3091
R3960 dcell_lv_0.bb[8].n14 dcell_lv_0.bb[8].n13 29.6212
R3961 dcell_lv_0.bb[8].n0 dcell_lv_0.bb[8].t1 26.5955
R3962 dcell_lv_0.bb[8].n0 dcell_lv_0.bb[8].t3 26.5955
R3963 dcell_lv_0.bb[8].n17 dcell_lv_0.bb[8].t0 24.9236
R3964 dcell_lv_0.bb[8].n17 dcell_lv_0.bb[8].t2 24.9236
R3965 dcell_lv_0.bb[8].n13 dcell_lv_0.bb[8].n12 21.0816
R3966 dcell_lv_0.bb[8].n7 dcell_lv_0.bb[8].n6 20.0252
R3967 dcell_lv_0.bb[8].n15 dcell_lv_0.bb[8] 12.5445
R3968 dcell_lv_0.bb[8].n16 dcell_lv_0.bb[8] 11.2645
R3969 dcell_lv_0.bb[8].n15 dcell_lv_0.bb[8].n14 9.65467
R3970 dcell_lv_0.bb[8].n14 dcell_lv_0.bb[8].n4 9.30258
R3971 dcell_lv_0.bb[8].n16 dcell_lv_0.bb[8] 6.1445
R3972 dcell_lv_0.bb[8].n6 dcell_lv_0.bb[8] 5.92643
R3973 dcell_lv_0.bb[8] dcell_lv_0.bb[8].n15 4.8645
R3974 dcell_lv_0.bb[8] dcell_lv_0.bb[8].n16 4.65505
R3975 dcell_lv_0.bb[8].n12 dcell_lv_0.bb[8] 3.2005
R3976 dcell_lv_0.bb[8].n4 dcell_lv_0.bb[8] 3.0725
R3977 dcell_lv_0.bb[8].n10 dcell_lv_0.bb[8].n7 2.17042
R3978 dcell_lv_0.bb[8].n9 dcell_lv_0.bb[8] 2.10199
R3979 dcell_lv_0.bb[8] dcell_lv_0.bb[8].n1 2.0485
R3980 dcell_lv_0.bb[8].n1 dcell_lv_0.bb[8] 1.55202
R3981 dcell_lv_0.bb[8].n13 dcell_lv_0.bb[8] 1.32081
R3982 dcell_lv_0.bb[8] dcell_lv_0.bb[8].n10 0.611828
R3983 dcell_lv_0.bb[8].n7 dcell_lv_0.bb[8] 0.373547
R3984 dcell_lv_0.b[8].n7 dcell_lv_0.b[8].t7 241.536
R3985 dcell_lv_0.b[8].n5 dcell_lv_0.b[8].t14 241.536
R3986 dcell_lv_0.b[8].n10 dcell_lv_0.b[8].t17 230.363
R3987 dcell_lv_0.b[8].n2 dcell_lv_0.b[8].t5 230.155
R3988 dcell_lv_0.b[8].n17 dcell_lv_0.b[8].t11 230.155
R3989 dcell_lv_0.b[8].n13 dcell_lv_0.b[8].t12 229.369
R3990 dcell_lv_0.b[8].n16 dcell_lv_0.b[8].t4 229.369
R3991 dcell_lv_0.b[8].n23 dcell_lv_0.b[8].n22 208.964
R3992 dcell_lv_0.b[8] dcell_lv_0.b[8].n7 177.839
R3993 dcell_lv_0.b[8].n7 dcell_lv_0.b[8].t13 169.237
R3994 dcell_lv_0.b[8].n5 dcell_lv_0.b[8].t10 169.237
R3995 dcell_lv_0.b[8].n6 dcell_lv_0.b[8].n5 159.37
R3996 dcell_lv_0.b[8].n10 dcell_lv_0.b[8].t16 158.064
R3997 dcell_lv_0.b[8] dcell_lv_0.b[8].n16 157.927
R3998 dcell_lv_0.b[8].n2 dcell_lv_0.b[8].t9 157.856
R3999 dcell_lv_0.b[8].n17 dcell_lv_0.b[8].t6 157.856
R4000 dcell_lv_0.b[8].n13 dcell_lv_0.b[8].t8 157.07
R4001 dcell_lv_0.b[8].n16 dcell_lv_0.b[8].t15 157.07
R4002 dcell_lv_0.b[8].n14 dcell_lv_0.b[8].n13 153.423
R4003 dcell_lv_0.b[8].n3 dcell_lv_0.b[8].n2 152
R4004 dcell_lv_0.b[8].n11 dcell_lv_0.b[8].n10 152
R4005 dcell_lv_0.b[8].n18 dcell_lv_0.b[8].n17 152
R4006 dcell_lv_0.b[8] dcell_lv_0.b[8].n0 96.8352
R4007 dcell_lv_0.b[8].n21 dcell_lv_0.b[8].n20 44.3335
R4008 dcell_lv_0.b[8].n8 dcell_lv_0.b[8].n6 40.9264
R4009 dcell_lv_0.b[8].n12 dcell_lv_0.b[8].n11 33.9843
R4010 dcell_lv_0.b[8].n22 dcell_lv_0.b[8].t0 26.5955
R4011 dcell_lv_0.b[8].n22 dcell_lv_0.b[8].t1 26.5955
R4012 dcell_lv_0.b[8].n0 dcell_lv_0.b[8].t2 24.9236
R4013 dcell_lv_0.b[8].n0 dcell_lv_0.b[8].t3 24.9236
R4014 dcell_lv_0.b[8].n4 dcell_lv_0.b[8].n3 17.557
R4015 dcell_lv_0.b[8].n20 dcell_lv_0.b[8].n19 16.335
R4016 dcell_lv_0.b[8].n15 dcell_lv_0.b[8].n14 15.3266
R4017 dcell_lv_0.b[8].n19 dcell_lv_0.b[8] 13.1418
R4018 dcell_lv_0.b[8] dcell_lv_0.b[8].n21 13.0565
R4019 dcell_lv_0.b[8].n8 dcell_lv_0.b[8] 12.9576
R4020 dcell_lv_0.b[8] dcell_lv_0.b[8].n1 11.2645
R4021 dcell_lv_0.b[8].n19 dcell_lv_0.b[8].n18 7.9365
R4022 dcell_lv_0.b[8].n9 dcell_lv_0.b[8].n8 6.5302
R4023 dcell_lv_0.b[8].n1 dcell_lv_0.b[8] 6.1445
R4024 dcell_lv_0.b[8].n1 dcell_lv_0.b[8] 4.65505
R4025 dcell_lv_0.b[8].n14 dcell_lv_0.b[8] 4.5042
R4026 dcell_lv_0.b[8].n21 dcell_lv_0.b[8] 4.3525
R4027 dcell_lv_0.b[8].n6 dcell_lv_0.b[8] 3.49141
R4028 dcell_lv_0.b[8].n11 dcell_lv_0.b[8] 3.2005
R4029 dcell_lv_0.b[8].n18 dcell_lv_0.b[8] 2.3045
R4030 dcell_lv_0.b[8].n3 dcell_lv_0.b[8] 2.10199
R4031 dcell_lv_0.b[8].n23 dcell_lv_0.b[8] 2.0485
R4032 dcell_lv_0.b[8] dcell_lv_0.b[8].n23 1.55202
R4033 dcell_lv_0.b[8].n12 dcell_lv_0.b[8].n9 1.39698
R4034 dcell_lv_0.b[8].n20 dcell_lv_0.b[8].n15 1.06105
R4035 dcell_lv_0.b[8].n9 dcell_lv_0.b[8].n4 0.852062
R4036 dcell_lv_0.b[8] dcell_lv_0.b[8].n12 0.613781
R4037 dcell_lv_0.b[8].n15 dcell_lv_0.b[8] 0.3755
R4038 dcell_lv_0.b[8].n4 dcell_lv_0.b[8] 0.221203
R4039 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 593.163
R4040 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n3 224.776
R4041 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 132.067
R4042 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n3 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 26.5955
R4043 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n3 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 26.5955
R4044 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 3.76521
R4045 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 2.13158
R4046 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 2.0264
R4047 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 1.17559
R4048 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.921363
R4049 a_17038_n199.t0 a_17038_n199.t1 55.3905
R4050 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t5 732.702
R4051 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t7 230.155
R4052 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t4 229.369
R4053 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 208.964
R4054 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 157.927
R4055 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t6 157.856
R4056 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t8 157.07
R4057 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 152
R4058 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 96.8352
R4059 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 28.9524
R4060 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t0 26.5955
R4061 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t2 26.5955
R4062 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t3 24.9236
R4063 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t1 24.9236
R4064 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 14.5363
R4065 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 13.0565
R4066 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 12.5635
R4067 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 12.2776
R4068 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 11.2645
R4069 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 7.11161
R4070 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 6.74842
R4071 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 6.1445
R4072 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 4.65505
R4073 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 4.3525
R4074 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 2.13383
R4075 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 2.0485
R4076 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 1.55202
R4077 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 593.154
R4078 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 224.776
R4079 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 132.067
R4080 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 26.5955
R4081 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 26.5955
R4082 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 18.824
R4083 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 6.77697
R4084 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 4.15748
R4085 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 3.76521
R4086 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 1.17559
R4087 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.921363
R4088 decoder_3_0/decoder_2to4_1.bb[1].n14 decoder_3_0/decoder_2to4_1.bb[1].t13 241.536
R4089 decoder_3_0/decoder_2to4_1.bb[1].n16 decoder_3_0/decoder_2to4_1.bb[1].t15 241.536
R4090 decoder_3_0/decoder_2to4_1.bb[1].n8 decoder_3_0/decoder_2to4_1.bb[1].t17 230.155
R4091 decoder_3_0/decoder_2to4_1.bb[1].n6 decoder_3_0/decoder_2to4_1.bb[1].t18 230.155
R4092 decoder_3_0/decoder_2to4_1.bb[1].n5 decoder_3_0/decoder_2to4_1.bb[1].t19 229.369
R4093 decoder_3_0/decoder_2to4_1.bb[1].n11 decoder_3_0/decoder_2to4_1.bb[1].t11 228.649
R4094 decoder_3_0/decoder_2to4_1.bb[1].n2 decoder_3_0/decoder_2to4_1.bb[1].t7 212.081
R4095 decoder_3_0/decoder_2to4_1.bb[1].n3 decoder_3_0/decoder_2to4_1.bb[1].t9 212.081
R4096 decoder_3_0/decoder_2to4_1.bb[1].n1 decoder_3_0/decoder_2to4_1.bb[1].n0 208.965
R4097 decoder_3_0/decoder_2to4_1.bb[1].n4 decoder_3_0/decoder_2to4_1.bb[1].n3 186.001
R4098 decoder_3_0/decoder_2to4_1.bb[1].n14 decoder_3_0/decoder_2to4_1.bb[1].t12 169.237
R4099 decoder_3_0/decoder_2to4_1.bb[1].n16 decoder_3_0/decoder_2to4_1.bb[1].t10 169.237
R4100 decoder_3_0/decoder_2to4_1.bb[1] decoder_3_0/decoder_2to4_1.bb[1].n5 157.927
R4101 decoder_3_0/decoder_2to4_1.bb[1].n8 decoder_3_0/decoder_2to4_1.bb[1].t5 157.856
R4102 decoder_3_0/decoder_2to4_1.bb[1].n6 decoder_3_0/decoder_2to4_1.bb[1].t14 157.856
R4103 decoder_3_0/decoder_2to4_1.bb[1].n5 decoder_3_0/decoder_2to4_1.bb[1].t16 157.07
R4104 decoder_3_0/decoder_2to4_1.bb[1].n11 decoder_3_0/decoder_2to4_1.bb[1].t4 156.35
R4105 decoder_3_0/decoder_2to4_1.bb[1] decoder_3_0/decoder_2to4_1.bb[1].n14 154.744
R4106 decoder_3_0/decoder_2to4_1.bb[1] decoder_3_0/decoder_2to4_1.bb[1].n16 154.744
R4107 decoder_3_0/decoder_2to4_1.bb[1].n9 decoder_3_0/decoder_2to4_1.bb[1].n8 152
R4108 decoder_3_0/decoder_2to4_1.bb[1].n12 decoder_3_0/decoder_2to4_1.bb[1].n11 152
R4109 decoder_3_0/decoder_2to4_1.bb[1].n7 decoder_3_0/decoder_2to4_1.bb[1].n6 152
R4110 decoder_3_0/decoder_2to4_1.bb[1].n2 decoder_3_0/decoder_2to4_1.bb[1].t6 139.78
R4111 decoder_3_0/decoder_2to4_1.bb[1].n3 decoder_3_0/decoder_2to4_1.bb[1].t8 139.78
R4112 decoder_3_0/decoder_2to4_1.bb[1] decoder_3_0/decoder_2to4_1.bb[1].n22 96.8352
R4113 decoder_3_0/decoder_2to4_1.bb[1].n3 decoder_3_0/decoder_2to4_1.bb[1].n2 61.346
R4114 decoder_3_0/decoder_2to4_1.bb[1].n0 decoder_3_0/decoder_2to4_1.bb[1].t1 26.5955
R4115 decoder_3_0/decoder_2to4_1.bb[1].n0 decoder_3_0/decoder_2to4_1.bb[1].t3 26.5955
R4116 decoder_3_0/decoder_2to4_1.bb[1].n22 decoder_3_0/decoder_2to4_1.bb[1].t0 24.9236
R4117 decoder_3_0/decoder_2to4_1.bb[1].n22 decoder_3_0/decoder_2to4_1.bb[1].t2 24.9236
R4118 decoder_3_0/decoder_2to4_1.bb[1].n13 decoder_3_0/decoder_2to4_1.bb[1].n12 24.0766
R4119 decoder_3_0/decoder_2to4_1.bb[1].n18 decoder_3_0/decoder_2to4_1.bb[1] 23.888
R4120 decoder_3_0/decoder_2to4_1.bb[1].n15 decoder_3_0/decoder_2to4_1.bb[1] 19.8144
R4121 decoder_3_0/decoder_2to4_1.bb[1] decoder_3_0/decoder_2to4_1.bb[1].n7 19.6746
R4122 decoder_3_0/decoder_2to4_1.bb[1].n10 decoder_3_0/decoder_2to4_1.bb[1].n9 19.5604
R4123 decoder_3_0/decoder_2to4_1.bb[1].n18 decoder_3_0/decoder_2to4_1.bb[1].n17 18.2347
R4124 decoder_3_0/decoder_2to4_1.bb[1].n17 decoder_3_0/decoder_2to4_1.bb[1] 17.3957
R4125 decoder_3_0/decoder_2to4_1.bb[1].n19 decoder_3_0/decoder_2to4_1.bb[1].n18 12.788
R4126 decoder_3_0/decoder_2to4_1.bb[1].n20 decoder_3_0/decoder_2to4_1.bb[1] 12.5445
R4127 decoder_3_0/decoder_2to4_1.bb[1].n21 decoder_3_0/decoder_2to4_1.bb[1] 11.2645
R4128 decoder_3_0/decoder_2to4_1.bb[1].n20 decoder_3_0/decoder_2to4_1.bb[1].n19 9.65467
R4129 decoder_3_0/decoder_2to4_1.bb[1].n19 decoder_3_0/decoder_2to4_1.bb[1].n4 9.30258
R4130 decoder_3_0/decoder_2to4_1.bb[1].n21 decoder_3_0/decoder_2to4_1.bb[1] 6.1445
R4131 decoder_3_0/decoder_2to4_1.bb[1].n12 decoder_3_0/decoder_2to4_1.bb[1] 6.13383
R4132 decoder_3_0/decoder_2to4_1.bb[1] decoder_3_0/decoder_2to4_1.bb[1].n20 4.8645
R4133 decoder_3_0/decoder_2to4_1.bb[1] decoder_3_0/decoder_2to4_1.bb[1].n21 4.65505
R4134 decoder_3_0/decoder_2to4_1.bb[1].n4 decoder_3_0/decoder_2to4_1.bb[1] 3.0725
R4135 decoder_3_0/decoder_2to4_1.bb[1].n7 decoder_3_0/decoder_2to4_1.bb[1] 2.13383
R4136 decoder_3_0/decoder_2to4_1.bb[1].n9 decoder_3_0/decoder_2to4_1.bb[1] 2.10199
R4137 decoder_3_0/decoder_2to4_1.bb[1] decoder_3_0/decoder_2to4_1.bb[1].n1 2.0485
R4138 decoder_3_0/decoder_2to4_1.bb[1].n1 decoder_3_0/decoder_2to4_1.bb[1] 1.55202
R4139 decoder_3_0/decoder_2to4_1.bb[1].n17 decoder_3_0/decoder_2to4_1.bb[1] 1.43019
R4140 decoder_3_0/decoder_2to4_1.bb[1].n15 decoder_3_0/decoder_2to4_1.bb[1].n13 1.08448
R4141 decoder_3_0/decoder_2to4_1.bb[1].n13 decoder_3_0/decoder_2to4_1.bb[1].n10 1.05323
R4142 decoder_3_0/decoder_2to4_1.bb[1] decoder_3_0/decoder_2to4_1.bb[1].n15 0.949719
R4143 decoder_3_0/decoder_2to4_1.bb[1].n10 decoder_3_0/decoder_2to4_1.bb[1] 0.0688594
R4144 a_7030_204.t0 a_7030_204.t1 60.9236
R4145 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n2 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n1 258.363
R4146 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n3 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t6 229.369
R4147 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n2 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n0 202.094
R4148 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n3 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t5 157.07
R4149 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n4 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n3 152
R4150 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n6 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t3 132.982
R4151 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n6 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n5 61.3652
R4152 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n0 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t2 32.5055
R4153 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n0 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t1 32.5055
R4154 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n1 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t0 26.5955
R4155 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n1 dcell_lv_0.seg_selector_logic_0.x3/x3.B.t4 26.5955
R4156 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n5 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n4 19.8407
R4157 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n4 dcell_lv_0.seg_selector_logic_0.x3/x3.B 5.92643
R4158 dcell_lv_0.seg_selector_logic_0.x3/x3.B dcell_lv_0.seg_selector_logic_0.x3/x3.B.n6 4.04261
R4159 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n5 dcell_lv_0.seg_selector_logic_0.x3/x3.B.n2 1.12991
R4160 a_23732_943.t0 a_23732_943.t1 65.941
R4161 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t4 732.773
R4162 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t6 212.081
R4163 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t8 212.081
R4164 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 208.965
R4165 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 186.001
R4166 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t5 139.78
R4167 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t7 139.78
R4168 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 96.8352
R4169 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 61.346
R4170 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t3 26.5955
R4171 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t1 26.5955
R4172 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t2 24.9236
R4173 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t0 24.9236
R4174 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 21.888
R4175 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 12.5445
R4176 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 11.2645
R4177 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 9.65467
R4178 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 9.30258
R4179 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 6.1445
R4180 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 4.8645
R4181 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 4.65505
R4182 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 3.0725
R4183 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 2.0485
R4184 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 1.55202
R4185 a_16088_n709.t0 a_16088_n709.t1 114.052
R4186 dec1[0].n0 dec1[0].t1 334.771
R4187 dec1[0].n1 dec1[0].t2 126.278
R4188 dec1[0].n2 dec1[0].t4 125.566
R4189 dec1[0].n1 dec1[0].t3 125.566
R4190 dec1[0].n0 dec1[0].t0 87.8568
R4191 dec1[0] dec1[0].n3 5.013
R4192 dec1[0].n3 dec1[0].n2 4.68383
R4193 dec1[0].n3 dec1[0].n0 0.876942
R4194 dec1[0].n2 dec1[0].n1 0.713
R4195 a_23732_685.t0 a_23732_685.t1 65.941
R4196 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t15 732.702
R4197 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t12 241.536
R4198 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t5 230.155
R4199 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t14 230.155
R4200 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t8 230.155
R4201 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t7 230.155
R4202 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t17 230.155
R4203 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t18 230.155
R4204 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 208.964
R4205 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 177.839
R4206 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t6 169.237
R4207 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t10 157.856
R4208 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t13 157.856
R4209 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t16 157.856
R4210 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t4 157.856
R4211 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t9 157.856
R4212 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t11 157.856
R4213 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 154.867
R4214 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 153.72
R4215 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 153.529
R4216 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 152
R4217 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 152
R4218 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 152
R4219 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 96.8352
R4220 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t0 26.5955
R4221 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t1 26.5955
R4222 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 25.9222
R4223 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t2 24.9236
R4224 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t3 24.9236
R4225 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 22.9626
R4226 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 22.4345
R4227 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 21.542
R4228 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 20.5115
R4229 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 19.8793
R4230 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 18.3823
R4231 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 13.0565
R4232 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 12.1443
R4233 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 11.2645
R4234 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 11.1817
R4235 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 10.7179
R4236 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 9.3005
R4237 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 6.38175
R4238 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 6.1445
R4239 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 5.23106
R4240 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 4.65505
R4241 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 4.3525
R4242 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 2.86617
R4243 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 2.67513
R4244 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 2.10199
R4245 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 2.10199
R4246 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 2.10199
R4247 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 2.0485
R4248 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 1.55202
R4249 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 1.52886
R4250 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 1.23683
R4251 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 0.926281
R4252 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 0.918469
R4253 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 0.842297
R4254 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.484875
R4255 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.00245312
R4256 a_6682_n1748.t0 a_6682_n1748.t1 49.8467
R4257 dcell_lv_0.logic_shift_seg2_0.x7.Y dcell_lv_0.logic_shift_seg2_0.x7.Y.n0 237.577
R4258 dcell_lv_0.logic_shift_seg2_0.x7.Y.n2 dcell_lv_0.logic_shift_seg2_0.x7.Y.t4 230.363
R4259 dcell_lv_0.logic_shift_seg2_0.x7.Y.n2 dcell_lv_0.logic_shift_seg2_0.x7.Y.t3 158.064
R4260 dcell_lv_0.logic_shift_seg2_0.x7.Y.n3 dcell_lv_0.logic_shift_seg2_0.x7.Y.n2 152.553
R4261 dcell_lv_0.logic_shift_seg2_0.x7.Y.n1 dcell_lv_0.logic_shift_seg2_0.x7.Y.t2 140.53
R4262 dcell_lv_0.logic_shift_seg2_0.x7.Y.n0 dcell_lv_0.logic_shift_seg2_0.x7.Y.t1 26.5955
R4263 dcell_lv_0.logic_shift_seg2_0.x7.Y.n0 dcell_lv_0.logic_shift_seg2_0.x7.Y.t0 26.5955
R4264 dcell_lv_0.logic_shift_seg2_0.x7.Y.n4 dcell_lv_0.logic_shift_seg2_0.x7.Y.n3 20.0033
R4265 dcell_lv_0.logic_shift_seg2_0.x7.Y dcell_lv_0.logic_shift_seg2_0.x7.Y.n4 11.2946
R4266 dcell_lv_0.logic_shift_seg2_0.x7.Y.n1 dcell_lv_0.logic_shift_seg2_0.x7.Y 9.03579
R4267 dcell_lv_0.logic_shift_seg2_0.x7.Y.n4 dcell_lv_0.logic_shift_seg2_0.x7.Y.n1 5.27109
R4268 dcell_lv_0.logic_shift_seg2_0.x7.Y.n1 dcell_lv_0.logic_shift_seg2_0.x7.Y 1.72748
R4269 dcell_lv_0.logic_shift_seg2_0.x7.Y.n3 dcell_lv_0.logic_shift_seg2_0.x7.Y 1.54533
R4270 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t0 227.856
R4271 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n0 152.333
R4272 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t2 140.382
R4273 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t3 114.031
R4274 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t1 83.3993
R4275 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t4 81.5883
R4276 lvsf_7bit_0/lvsf_buff_4/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n1 14.4422
R4277 lvsf_7bit_0/lvsf_buff_4/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n3 7.56882
R4278 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n2 5.08175
R4279 lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_4/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R4280 a_19454_n199.t0 a_19454_n199.t1 55.3905
R4281 a_18858_n296.t0 a_18858_n296.n0 228.04
R4282 a_18858_n296.n0 a_18858_n296.t2 145.648
R4283 a_18858_n296.n0 a_18858_n296.t1 83.2159
R4284 dcell_lv_0.seg_selector_logic_0.x2/x4.A dcell_lv_0.seg_selector_logic_0.x2/x4.A.n3 237.577
R4285 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n0 dcell_lv_0.seg_selector_logic_0.x2/x4.A.t4 228.649
R4286 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n0 dcell_lv_0.seg_selector_logic_0.x2/x4.A.t3 156.35
R4287 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n1 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n0 152
R4288 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n2 dcell_lv_0.seg_selector_logic_0.x2/x4.A.t2 131.691
R4289 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n2 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n1 35.0201
R4290 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n3 dcell_lv_0.seg_selector_logic_0.x2/x4.A.t1 26.5955
R4291 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n3 dcell_lv_0.seg_selector_logic_0.x2/x4.A.t0 26.5955
R4292 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n4 dcell_lv_0.seg_selector_logic_0.x2/x4.A 16.5652
R4293 dcell_lv_0.seg_selector_logic_0.x2/x4.A dcell_lv_0.seg_selector_logic_0.x2/x4.A.n4 9.03579
R4294 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n4 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n2 8.8386
R4295 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n4 dcell_lv_0.seg_selector_logic_0.x2/x4.A 1.72748
R4296 dcell_lv_0.seg_selector_logic_0.x2/x4.A.n1 dcell_lv_0.seg_selector_logic_0.x2/x4.A 1.43334
R4297 a_7766_n660.t0 a_7766_n660.t1 60.9236
R4298 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n2 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t7 732.662
R4299 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n7 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n6 258.363
R4300 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n0 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t6 230.576
R4301 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n7 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n5 202.094
R4302 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n0 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t5 158.275
R4303 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n1 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n0 152
R4304 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n4 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t2 126.469
R4305 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n8 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n7 62.4946
R4306 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n5 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t1 32.5055
R4307 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n5 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t0 32.5055
R4308 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n6 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t3 26.5955
R4309 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n6 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t4 26.5955
R4310 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n2 19.9547
R4311 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n3 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 13.6567
R4312 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n3 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n1 12.0102
R4313 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n4 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n3 9.82192
R4314 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n1 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 6.66717
R4315 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n8 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n4 6.51278
R4316 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n8 4.04261
R4317 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n2 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.110917
R4318 a_15888_n296.n0 a_15888_n296.t1 228.04
R4319 a_15888_n296.n0 a_15888_n296.t2 145.648
R4320 a_15888_n296.t0 a_15888_n296.n0 83.2159
R4321 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t0 227.856
R4322 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n0 152.333
R4323 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t3 140.382
R4324 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t2 114.031
R4325 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t1 83.3993
R4326 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t4 81.5883
R4327 lvsf_7bit_0/lvsf_buff_3/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n1 14.4422
R4328 lvsf_7bit_0/lvsf_buff_3/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n3 7.56882
R4329 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n2 5.08175
R4330 lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_3/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R4331 a_16048_n199.t0 a_16048_n199.t1 55.3905
R4332 dec0[2].n0 dec0[2].t1 334.788
R4333 dec0[2].n2 dec0[2].t4 126.27
R4334 dec0[2].n2 dec0[2].t2 125.558
R4335 dec0[2].n1 dec0[2].t3 121.127
R4336 dec0[2].n0 dec0[2].t0 87.8063
R4337 dec0[2].n3 dec0[2].n2 5.73592
R4338 dec0[2] dec0[2].n3 5.37342
R4339 dec0[2].n1 dec0[2].n0 0.322615
R4340 dec0[2].n3 dec0[2].n1 0.177583
R4341 a_24472_427.t0 a_24472_427.t1 65.941
R4342 a_24472_685.t0 a_24472_685.t1 65.941
R4343 VBNLV.n2 VBNLV.t13 124.9
R4344 VBNLV.n3 VBNLV.t4 124.9
R4345 VBNLV.n4 VBNLV.t14 124.9
R4346 VBNLV.n5 VBNLV.t9 124.9
R4347 VBNLV.n6 VBNLV.t18 124.9
R4348 VBNLV.n7 VBNLV.t15 124.9
R4349 VBNLV.n8 VBNLV.t0 124.9
R4350 VBNLV.n9 VBNLV.t19 124.9
R4351 VBNLV.n10 VBNLV.t5 124.9
R4352 VBNLV.n11 VBNLV.t1 124.9
R4353 VBNLV.n12 VBNLV.t16 124.9
R4354 VBNLV.n13 VBNLV.t6 124.9
R4355 VBNLV.n14 VBNLV.t20 124.9
R4356 VBNLV.n15 VBNLV.t11 124.9
R4357 VBNLV.n16 VBNLV.t2 124.9
R4358 VBNLV.n17 VBNLV.t21 124.9
R4359 VBNLV.n18 VBNLV.t7 124.9
R4360 VBNLV.n19 VBNLV.t3 124.9
R4361 VBNLV.n20 VBNLV.t12 124.9
R4362 VBNLV.n21 VBNLV.t8 124.9
R4363 VBNLV.n1 VBNLV.t17 124.9
R4364 VBNLV.n0 VBNLV.t10 124.9
R4365 VBNLV.n1 VBNLV.n0 1.27824
R4366 VBNLV.n21 VBNLV.n20 1.27824
R4367 VBNLV.n19 VBNLV.n18 1.27824
R4368 VBNLV.n17 VBNLV.n16 1.27824
R4369 VBNLV.n15 VBNLV.n14 1.27824
R4370 VBNLV.n13 VBNLV.n12 1.27824
R4371 VBNLV.n11 VBNLV.n10 1.27824
R4372 VBNLV.n9 VBNLV.n8 1.27824
R4373 VBNLV.n7 VBNLV.n6 1.27824
R4374 VBNLV.n5 VBNLV.n4 1.27824
R4375 VBNLV.n3 VBNLV.n2 1.27824
R4376 VBNLV VBNLV.n1 0.391454
R4377 VBNLV VBNLV.n21 0.391454
R4378 VBNLV.n20 VBNLV 0.391454
R4379 VBNLV VBNLV.n19 0.391454
R4380 VBNLV.n18 VBNLV 0.391454
R4381 VBNLV VBNLV.n17 0.391454
R4382 VBNLV.n16 VBNLV 0.391454
R4383 VBNLV VBNLV.n15 0.391454
R4384 VBNLV.n14 VBNLV 0.391454
R4385 VBNLV VBNLV.n13 0.391454
R4386 VBNLV.n12 VBNLV 0.391454
R4387 VBNLV VBNLV.n11 0.391454
R4388 VBNLV.n10 VBNLV 0.391454
R4389 VBNLV VBNLV.n9 0.391454
R4390 VBNLV.n8 VBNLV 0.391454
R4391 VBNLV VBNLV.n7 0.391454
R4392 VBNLV.n6 VBNLV 0.391454
R4393 VBNLV VBNLV.n5 0.391454
R4394 VBNLV.n4 VBNLV 0.391454
R4395 VBNLV VBNLV.n3 0.391454
R4396 VBNLV.n2 VBNLV 0.391454
R4397 VBNLV.n0 VBNLV 0.266454
R4398 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n1 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t0 227.856
R4399 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R4400 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n2 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t2 140.163
R4401 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n0 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t3 114.031
R4402 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n1 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t1 83.3993
R4403 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n0 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t4 81.5883
R4404 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n3 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R4405 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n3 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R4406 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R4407 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n2 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R4408 a_13118_n709.t0 a_13118_n709.t1 114.052
R4409 dcell_lv_0.seg_selector_logic_0.x1/x3.B dcell_lv_0.seg_selector_logic_0.x1/x3.B.n3 237.577
R4410 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n0 dcell_lv_0.seg_selector_logic_0.x1/x3.B.t4 230.363
R4411 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n0 dcell_lv_0.seg_selector_logic_0.x1/x3.B.t3 158.064
R4412 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n1 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n0 153.28
R4413 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n2 dcell_lv_0.seg_selector_logic_0.x1/x3.B.t2 132.81
R4414 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n3 dcell_lv_0.seg_selector_logic_0.x1/x3.B.t1 26.5955
R4415 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n3 dcell_lv_0.seg_selector_logic_0.x1/x3.B.t0 26.5955
R4416 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n2 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n1 19.4367
R4417 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n4 dcell_lv_0.seg_selector_logic_0.x1/x3.B 16.5652
R4418 dcell_lv_0.seg_selector_logic_0.x1/x3.B dcell_lv_0.seg_selector_logic_0.x1/x3.B.n4 9.03579
R4419 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n4 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n2 7.72113
R4420 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n1 dcell_lv_0.seg_selector_logic_0.x1/x3.B 5.1205
R4421 dcell_lv_0.seg_selector_logic_0.x1/x3.B.n4 dcell_lv_0.seg_selector_logic_0.x1/x3.B 1.72748
R4422 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n1 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t5 732.662
R4423 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n2 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t4 230.576
R4424 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n6 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t1 218.572
R4425 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n2 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t3 158.275
R4426 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n3 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n2 152
R4427 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n5 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n0 94.1864
R4428 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n6 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n5 86.3316
R4429 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n0 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t2 24.9236
R4430 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n0 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t0 24.9236
R4431 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n5 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n4 21.3341
R4432 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n1 10.6809
R4433 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n4 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n3 9.3005
R4434 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n6 7.54721
R4435 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n3 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 6.66717
R4436 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n4 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 3.48572
R4437 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n1 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.110917
R4438 dec0[3].n0 dec0[3].t1 334.822
R4439 dec0[3].n1 dec0[3].t3 126.27
R4440 dec0[3].n1 dec0[3].t2 125.558
R4441 dec0[3].n2 dec0[3].t4 125.558
R4442 dec0[3].n0 dec0[3].t0 87.8063
R4443 dec0[3].n3 dec0[3].n2 5.73592
R4444 dec0[3] dec0[3].n3 5.64217
R4445 dec0[3].n2 dec0[3].n1 0.713
R4446 dec0[3].n3 dec0[3].n0 0.197295
R4447 a_25156_427.t0 a_25156_427.t1 65.941
R4448 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t9 732.773
R4449 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t6 230.155
R4450 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t4 229.369
R4451 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t8 212.081
R4452 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t11 212.081
R4453 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 208.965
R4454 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 186.001
R4455 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 157.927
R4456 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t5 157.856
R4457 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t12 157.07
R4458 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 152
R4459 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t7 139.78
R4460 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t10 139.78
R4461 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 96.8352
R4462 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 61.346
R4463 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t3 26.5955
R4464 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t1 26.5955
R4465 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t2 24.9236
R4466 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t0 24.9236
R4467 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 19.6746
R4468 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 19.6318
R4469 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 12.5445
R4470 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 11.3943
R4471 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 11.2645
R4472 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 9.65467
R4473 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 9.30258
R4474 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 6.49425
R4475 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 6.1445
R4476 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 4.8645
R4477 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 4.65505
R4478 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 3.0725
R4479 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 2.13383
R4480 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 2.0485
R4481 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 1.55202
R4482 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t4 732.662
R4483 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t5 230.576
R4484 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n8 224.776
R4485 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n7 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 217.601
R4486 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t3 158.275
R4487 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 152.8
R4488 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t1 132.067
R4489 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n7 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 64.0005
R4490 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n8 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t2 26.5955
R4491 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n8 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t0 26.5955
R4492 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 15.377
R4493 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 10.1396
R4494 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 9.57008
R4495 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 5.86717
R4496 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 5.80407
R4497 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n7 3.38874
R4498 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 2.6841
R4499 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 1.47388
R4500 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 1.17559
R4501 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 0.921363
R4502 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 0.0400833
R4503 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t2 732.662
R4504 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t0 230.518
R4505 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t1 162.351
R4506 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 23.694
R4507 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n1 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB 14.6392
R4508 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n1 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB 11.6875
R4509 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n1 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB 7.23528
R4510 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n1 5.04292
R4511 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB 0.110917
R4512 a_7510_428.t0 a_7510_428.t1 49.8467
R4513 dcell_lv_0.seg_selector_logic_0.x1/x3.A dcell_lv_0.seg_selector_logic_0.x1/x3.A.n0 237.577
R4514 dcell_lv_0.seg_selector_logic_0.x1/x3.A.n2 dcell_lv_0.seg_selector_logic_0.x1/x3.A.t3 231.835
R4515 dcell_lv_0.seg_selector_logic_0.x1/x3.A.n2 dcell_lv_0.seg_selector_logic_0.x1/x3.A.t4 157.07
R4516 dcell_lv_0.seg_selector_logic_0.x1/x3.A dcell_lv_0.seg_selector_logic_0.x1/x3.A.n2 154.304
R4517 dcell_lv_0.seg_selector_logic_0.x1/x3.A.n1 dcell_lv_0.seg_selector_logic_0.x1/x3.A.t2 140.53
R4518 dcell_lv_0.seg_selector_logic_0.x1/x3.A.n3 dcell_lv_0.seg_selector_logic_0.x1/x3.A 32.1479
R4519 dcell_lv_0.seg_selector_logic_0.x1/x3.A.n0 dcell_lv_0.seg_selector_logic_0.x1/x3.A.t1 26.5955
R4520 dcell_lv_0.seg_selector_logic_0.x1/x3.A.n0 dcell_lv_0.seg_selector_logic_0.x1/x3.A.t0 26.5955
R4521 dcell_lv_0.seg_selector_logic_0.x1/x3.A dcell_lv_0.seg_selector_logic_0.x1/x3.A.n3 14.3064
R4522 dcell_lv_0.seg_selector_logic_0.x1/x3.A.n1 dcell_lv_0.seg_selector_logic_0.x1/x3.A 9.03579
R4523 dcell_lv_0.seg_selector_logic_0.x1/x3.A.n3 dcell_lv_0.seg_selector_logic_0.x1/x3.A.n1 2.25932
R4524 dcell_lv_0.seg_selector_logic_0.x1/x3.A.n1 dcell_lv_0.seg_selector_logic_0.x1/x3.A 1.72748
R4525 bb[2].n4 bb[2].n3 863.124
R4526 bb[2].n3 bb[2].n2 585
R4527 bb[2].n1 bb[2].t1 490.913
R4528 bb[2].n7 bb[2].n6 152
R4529 bb[2].n0 bb[2].t0 144.376
R4530 bb[2].n3 bb[2].t1 140.738
R4531 bb[2].n6 bb[2].t2 114.031
R4532 bb[2].n6 bb[2].t3 81.5883
R4533 bb[2] bb[2].n7 16.7132
R4534 bb[2] bb[2].n5 13.7979
R4535 bb[2] bb[2].n0 11.3477
R4536 bb[2] bb[2].n1 11.2054
R4537 bb[2].n2 bb[2] 8.81089
R4538 bb[2] bb[2].n4 7.61955
R4539 bb[2].n5 bb[2] 7.17626
R4540 bb[2].n5 bb[2] 6.59444
R4541 bb[2].n4 bb[2] 4.98751
R4542 bb[2].n2 bb[2] 3.49141
R4543 bb[2].n0 bb[2] 2.94838
R4544 bb[2].n5 bb[2] 2.16154
R4545 bb[2].n7 bb[2] 1.16414
R4546 bb[2].n1 bb[2] 1.09557
R4547 b[2].n4 b[2].n3 863.124
R4548 b[2].n3 b[2].n2 585
R4549 b[2].n1 b[2].t1 490.913
R4550 b[2].n0 b[2].t0 144.376
R4551 b[2].n3 b[2].t1 140.738
R4552 b[2] b[2].n5 14.3755
R4553 b[2].n5 b[2] 13.5763
R4554 b[2] b[2].n0 11.3477
R4555 b[2] b[2].n1 11.2054
R4556 b[2].n2 b[2] 8.81089
R4557 b[2] b[2].n4 7.61955
R4558 b[2].n4 b[2] 4.98751
R4559 b[2].n2 b[2] 3.49141
R4560 b[2].n0 b[2] 2.94838
R4561 b[2].n1 b[2] 1.09557
R4562 b[2].n5 b[2] 0.776258
R4563 a_14374_n1619.t0 a_14374_n1619.t1 114.052
R4564 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n1 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t0 227.856
R4565 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R4566 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n2 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t4 140.163
R4567 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n0 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t2 114.031
R4568 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n1 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t1 83.3993
R4569 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n0 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t3 81.5883
R4570 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n3 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R4571 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n3 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R4572 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R4573 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n2 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R4574 SH[1].n5 SH[1].n4 863.124
R4575 SH[1].n4 SH[1].n3 585
R4576 SH[1].n2 SH[1].t1 490.913
R4577 SH[1].n0 SH[1].t0 144.376
R4578 SH[1].n4 SH[1].t1 140.738
R4579 SH[1].n1 SH[1] 14.4526
R4580 SH[1].n1 SH[1] 13.9641
R4581 SH[1] SH[1].n0 11.3477
R4582 SH[1] SH[1].n2 11.2054
R4583 SH[1].n3 SH[1] 8.81089
R4584 SH[1] SH[1].n5 7.61955
R4585 SH[1].n5 SH[1] 4.98751
R4586 SH[1].n3 SH[1] 3.49141
R4587 SH[1].n0 SH[1] 2.94838
R4588 SH[1].n2 SH[1] 1.09557
R4589 SH[1] SH[1].n1 0.388379
R4590 a_7786_428.t0 a_7786_428.t1 49.8467
R4591 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t0 227.856
R4592 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n0 152.333
R4593 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t4 140.382
R4594 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t2 114.031
R4595 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t1 83.3993
R4596 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t3 81.5883
R4597 lvsf_7bit_0/lvsf_buff_2/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n1 14.4422
R4598 lvsf_7bit_0/lvsf_buff_2/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n3 7.56882
R4599 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n2 5.08175
R4600 lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_2/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R4601 bb[3].n4 bb[3].n3 863.124
R4602 bb[3].n3 bb[3].n2 585
R4603 bb[3].n1 bb[3].t1 490.913
R4604 bb[3].n7 bb[3].n6 152
R4605 bb[3].n0 bb[3].t0 144.376
R4606 bb[3].n3 bb[3].t1 140.738
R4607 bb[3].n6 bb[3].t2 114.031
R4608 bb[3].n6 bb[3].t3 81.5883
R4609 bb[3] bb[3].n7 16.7132
R4610 bb[3] bb[3].n5 13.7979
R4611 bb[3] bb[3].n0 11.3477
R4612 bb[3] bb[3].n1 11.2054
R4613 bb[3].n2 bb[3] 8.81089
R4614 bb[3] bb[3].n4 7.61955
R4615 bb[3].n5 bb[3] 7.17626
R4616 bb[3].n5 bb[3] 6.59444
R4617 bb[3].n4 bb[3] 4.98751
R4618 bb[3].n2 bb[3] 3.49141
R4619 bb[3].n0 bb[3] 2.94838
R4620 bb[3].n5 bb[3] 2.16154
R4621 bb[3].n7 bb[3] 1.16414
R4622 bb[3].n1 bb[3] 1.09557
R4623 decoder_3_0/decoder_2to4_2.b[0].n9 decoder_3_0/decoder_2to4_2.b[0].t2 230.712
R4624 decoder_3_0/decoder_2to4_2.b[0].n7 decoder_3_0/decoder_2to4_2.b[0].t4 230.576
R4625 decoder_3_0/decoder_2to4_2.b[0].n2 decoder_3_0/decoder_2to4_2.b[0].t5 230.155
R4626 decoder_3_0/decoder_2to4_2.b[0].n0 decoder_3_0/decoder_2to4_2.b[0].t7 230.155
R4627 decoder_3_0/decoder_2to4_2.b[0].n11 decoder_3_0/decoder_2to4_2.b[0].n10 205.28
R4628 decoder_3_0/decoder_2to4_2.b[0].n7 decoder_3_0/decoder_2to4_2.b[0].t9 158.275
R4629 decoder_3_0/decoder_2to4_2.b[0].n2 decoder_3_0/decoder_2to4_2.b[0].t8 157.856
R4630 decoder_3_0/decoder_2to4_2.b[0].n0 decoder_3_0/decoder_2to4_2.b[0].t6 157.856
R4631 decoder_3_0/decoder_2to4_2.b[0].n3 decoder_3_0/decoder_2to4_2.b[0].n2 153.72
R4632 decoder_3_0/decoder_2to4_2.b[0].n1 decoder_3_0/decoder_2to4_2.b[0].n0 153.529
R4633 decoder_3_0/decoder_2to4_2.b[0].n8 decoder_3_0/decoder_2to4_2.b[0].n7 153.067
R4634 decoder_3_0/decoder_2to4_2.b[0].n6 decoder_3_0/decoder_2to4_2.b[0].t1 135.947
R4635 decoder_3_0/decoder_2to4_2.b[0] decoder_3_0/decoder_2to4_2.b[0].n11 67.4857
R4636 decoder_3_0/decoder_2to4_2.b[0].n11 decoder_3_0/decoder_2to4_2.b[0].n9 44.0818
R4637 decoder_3_0/decoder_2to4_2.b[0] decoder_3_0/decoder_2to4_2.b[0].n6 33.5064
R4638 decoder_3_0/decoder_2to4_2.b[0].n10 decoder_3_0/decoder_2to4_2.b[0].t3 26.5955
R4639 decoder_3_0/decoder_2to4_2.b[0].n10 decoder_3_0/decoder_2to4_2.b[0].t0 26.5955
R4640 decoder_3_0/decoder_2to4_2.b[0] decoder_3_0/decoder_2to4_2.b[0].n5 23.9017
R4641 decoder_3_0/decoder_2to4_2.b[0].n9 decoder_3_0/decoder_2to4_2.b[0].n8 19.3316
R4642 decoder_3_0/decoder_2to4_2.b[0].n6 decoder_3_0/decoder_2to4_2.b[0] 16.4149
R4643 decoder_3_0/decoder_2to4_2.b[0].n4 decoder_3_0/decoder_2to4_2.b[0].n1 10.7179
R4644 decoder_3_0/decoder_2to4_2.b[0].n4 decoder_3_0/decoder_2to4_2.b[0].n3 9.3005
R4645 decoder_3_0/decoder_2to4_2.b[0].n8 decoder_3_0/decoder_2to4_2.b[0] 5.6005
R4646 decoder_3_0/decoder_2to4_2.b[0].n5 decoder_3_0/decoder_2to4_2.b[0].n4 5.04981
R4647 decoder_3_0/decoder_2to4_2.b[0].n1 decoder_3_0/decoder_2to4_2.b[0] 2.86617
R4648 decoder_3_0/decoder_2to4_2.b[0].n3 decoder_3_0/decoder_2to4_2.b[0] 2.67513
R4649 decoder_3_0/decoder_2to4_2.b[0].n5 decoder_3_0/decoder_2to4_2.b[0] 0.18175
R4650 b[3].n4 b[3].n3 863.124
R4651 b[3].n3 b[3].n2 585
R4652 b[3].n1 b[3].t1 490.913
R4653 b[3].n0 b[3].t0 144.376
R4654 b[3].n3 b[3].t1 140.738
R4655 b[3] b[3].n5 14.3755
R4656 b[3].n5 b[3] 13.5763
R4657 b[3] b[3].n0 11.3477
R4658 b[3] b[3].n1 11.2054
R4659 b[3].n2 b[3] 8.81089
R4660 b[3] b[3].n4 7.61955
R4661 b[3].n4 b[3] 4.98751
R4662 b[3].n2 b[3] 3.49141
R4663 b[3].n0 b[3] 2.94838
R4664 b[3].n1 b[3] 1.09557
R4665 b[3].n5 b[3] 0.776258
R4666 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n1 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t2 732.662
R4667 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n2 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t0 223.315
R4668 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t1 162.351
R4669 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n2 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 15.4066
R4670 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n0 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 11.6875
R4671 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n1 10.7065
R4672 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n0 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 7.23528
R4673 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n2 7.20375
R4674 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n0 5.04292
R4675 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n1 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.0400833
R4676 dcell_lv_0.logic_shift_seg2_0.x6.Y.n2 dcell_lv_0.logic_shift_seg2_0.x6.Y.t0 268.077
R4677 dcell_lv_0.logic_shift_seg2_0.x6.Y.n2 dcell_lv_0.logic_shift_seg2_0.x6.Y.t0 258.846
R4678 dcell_lv_0.logic_shift_seg2_0.x6.Y.n1 dcell_lv_0.logic_shift_seg2_0.x6.Y.t4 241.536
R4679 dcell_lv_0.logic_shift_seg2_0.x6.Y dcell_lv_0.logic_shift_seg2_0.x6.Y.n0 237.577
R4680 dcell_lv_0.logic_shift_seg2_0.x6.Y.n1 dcell_lv_0.logic_shift_seg2_0.x6.Y.t3 169.237
R4681 dcell_lv_0.logic_shift_seg2_0.x6.Y dcell_lv_0.logic_shift_seg2_0.x6.Y.n1 153.877
R4682 dcell_lv_0.logic_shift_seg2_0.x6.Y.n2 dcell_lv_0.logic_shift_seg2_0.x6.Y 29.7595
R4683 dcell_lv_0.logic_shift_seg2_0.x6.Y.n0 dcell_lv_0.logic_shift_seg2_0.x6.Y.t1 26.5955
R4684 dcell_lv_0.logic_shift_seg2_0.x6.Y.n0 dcell_lv_0.logic_shift_seg2_0.x6.Y.t2 26.5955
R4685 dcell_lv_0.logic_shift_seg2_0.x6.Y.n3 dcell_lv_0.logic_shift_seg2_0.x6.Y 16.5652
R4686 dcell_lv_0.logic_shift_seg2_0.x6.Y.n3 dcell_lv_0.logic_shift_seg2_0.x6.Y 9.03579
R4687 dcell_lv_0.logic_shift_seg2_0.x6.Y.n3 dcell_lv_0.logic_shift_seg2_0.x6.Y.n2 8.8386
R4688 dcell_lv_0.logic_shift_seg2_0.x6.Y dcell_lv_0.logic_shift_seg2_0.x6.Y.n3 1.72748
R4689 a_7046_n1748.t0 a_7046_n1748.t1 49.8467
R4690 a_7130_n1748.t0 a_7130_n1748.t1 60.9236
R4691 DIN6.n0 DIN6.t1 212.081
R4692 DIN6.n1 DIN6.t3 212.081
R4693 DIN6.n2 DIN6.n1 183.185
R4694 DIN6.n0 DIN6.t0 139.78
R4695 DIN6.n1 DIN6.t2 139.78
R4696 DIN6.n1 DIN6.n0 61.346
R4697 DIN6.n3 DIN6.n2 9.30224
R4698 DIN6.n2 DIN6 5.8885
R4699 DIN6.n3 DIN6 5.1005
R4700 DIN6 DIN6.n3 0.0525833
R4701 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t0 227.856
R4702 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n0 152.333
R4703 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t4 140.382
R4704 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t2 114.031
R4705 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t1 83.3993
R4706 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t3 81.5883
R4707 lvsf_7bit_0/lvsf_buff_5/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n1 14.4422
R4708 lvsf_7bit_0/lvsf_buff_5/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n3 7.56882
R4709 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n2 5.08175
R4710 lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_5/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R4711 bb[4].n4 bb[4].n3 863.124
R4712 bb[4].n3 bb[4].n2 585
R4713 bb[4].n1 bb[4].t1 490.913
R4714 bb[4].n7 bb[4].n6 152
R4715 bb[4].n0 bb[4].t0 144.376
R4716 bb[4].n3 bb[4].t1 140.738
R4717 bb[4].n6 bb[4].t2 114.031
R4718 bb[4].n6 bb[4].t3 81.5883
R4719 bb[4] bb[4].n7 16.7132
R4720 bb[4] bb[4].n5 13.7979
R4721 bb[4] bb[4].n0 11.3477
R4722 bb[4] bb[4].n1 11.2054
R4723 bb[4].n2 bb[4] 8.81089
R4724 bb[4] bb[4].n4 7.61955
R4725 bb[4].n5 bb[4] 7.17626
R4726 bb[4].n5 bb[4] 6.59444
R4727 bb[4].n4 bb[4] 4.98751
R4728 bb[4].n2 bb[4] 3.49141
R4729 bb[4].n0 bb[4] 2.94838
R4730 bb[4].n5 bb[4] 2.16154
R4731 bb[4].n7 bb[4] 1.16414
R4732 bb[4].n1 bb[4] 1.09557
R4733 b[4].n4 b[4].n3 863.124
R4734 b[4].n3 b[4].n2 585
R4735 b[4].n1 b[4].t1 490.913
R4736 b[4].n0 b[4].t0 144.376
R4737 b[4].n3 b[4].t1 140.738
R4738 b[4] b[4].n5 14.3755
R4739 b[4].n5 b[4] 13.5763
R4740 b[4] b[4].n0 11.3477
R4741 b[4] b[4].n1 11.2054
R4742 b[4].n2 b[4] 8.81089
R4743 b[4] b[4].n4 7.61955
R4744 b[4].n4 b[4] 4.98751
R4745 b[4].n2 b[4] 3.49141
R4746 b[4].n0 b[4] 2.94838
R4747 b[4].n1 b[4] 1.09557
R4748 b[4].n5 b[4] 0.776258
R4749 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 593.163
R4750 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n3 224.776
R4751 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 132.067
R4752 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n3 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 26.5955
R4753 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n3 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 26.5955
R4754 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 3.76521
R4755 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 2.13158
R4756 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 2.0264
R4757 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 1.17559
R4758 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.921363
R4759 dcell_lv_0.logic_shift_seg2_0.x8.Y.n1 dcell_lv_0.logic_shift_seg2_0.x8.Y.t0 274.793
R4760 dcell_lv_0.logic_shift_seg2_0.x8.Y.n2 dcell_lv_0.logic_shift_seg2_0.x8.Y.t5 232.214
R4761 dcell_lv_0.logic_shift_seg2_0.x8.Y.n1 dcell_lv_0.logic_shift_seg2_0.x8.Y.n0 205.28
R4762 dcell_lv_0.logic_shift_seg2_0.x8.Y dcell_lv_0.logic_shift_seg2_0.x8.Y.t1 169.452
R4763 dcell_lv_0.logic_shift_seg2_0.x8.Y.n2 dcell_lv_0.logic_shift_seg2_0.x8.Y.t4 159.915
R4764 dcell_lv_0.logic_shift_seg2_0.x8.Y.n3 dcell_lv_0.logic_shift_seg2_0.x8.Y.n2 152
R4765 dcell_lv_0.logic_shift_seg2_0.x8.Y.n4 dcell_lv_0.logic_shift_seg2_0.x8.Y.n1 54.4975
R4766 dcell_lv_0.logic_shift_seg2_0.x8.Y.n0 dcell_lv_0.logic_shift_seg2_0.x8.Y.t3 26.5955
R4767 dcell_lv_0.logic_shift_seg2_0.x8.Y.n0 dcell_lv_0.logic_shift_seg2_0.x8.Y.t2 26.5955
R4768 dcell_lv_0.logic_shift_seg2_0.x8.Y.n4 dcell_lv_0.logic_shift_seg2_0.x8.Y.n3 23.9063
R4769 dcell_lv_0.logic_shift_seg2_0.x8.Y dcell_lv_0.logic_shift_seg2_0.x8.Y.n4 12.9887
R4770 dcell_lv_0.logic_shift_seg2_0.x8.Y.n3 dcell_lv_0.logic_shift_seg2_0.x8.Y 0.970197
R4771 a_19324_n1619.t0 a_19324_n1619.t1 114.052
R4772 bb[5].n4 bb[5].n3 863.124
R4773 bb[5].n3 bb[5].n2 585
R4774 bb[5].n1 bb[5].t1 490.913
R4775 bb[5].n7 bb[5].n6 152
R4776 bb[5].n0 bb[5].t0 144.376
R4777 bb[5].n3 bb[5].t1 140.738
R4778 bb[5].n6 bb[5].t2 114.031
R4779 bb[5].n6 bb[5].t3 81.5883
R4780 bb[5] bb[5].n7 16.7132
R4781 bb[5] bb[5].n5 13.7979
R4782 bb[5] bb[5].n0 11.3477
R4783 bb[5] bb[5].n1 11.2054
R4784 bb[5].n2 bb[5] 8.81089
R4785 bb[5] bb[5].n4 7.61955
R4786 bb[5].n5 bb[5] 7.17626
R4787 bb[5].n5 bb[5] 6.59444
R4788 bb[5].n4 bb[5] 4.98751
R4789 bb[5].n2 bb[5] 3.49141
R4790 bb[5].n0 bb[5] 2.94838
R4791 bb[5].n5 bb[5] 2.16154
R4792 bb[5].n7 bb[5] 1.16414
R4793 bb[5].n1 bb[5] 1.09557
R4794 b[5].n4 b[5].n3 863.124
R4795 b[5].n3 b[5].n2 585
R4796 b[5].n1 b[5].t1 490.913
R4797 b[5].n0 b[5].t0 144.376
R4798 b[5].n3 b[5].t1 140.738
R4799 b[5] b[5].n5 14.3755
R4800 b[5].n5 b[5] 13.5763
R4801 b[5] b[5].n0 11.3477
R4802 b[5] b[5].n1 11.2054
R4803 b[5].n2 b[5] 8.81089
R4804 b[5] b[5].n4 7.61955
R4805 b[5].n4 b[5] 4.98751
R4806 b[5].n2 b[5] 3.49141
R4807 b[5].n0 b[5] 2.94838
R4808 b[5].n1 b[5] 1.09557
R4809 b[5].n5 b[5] 0.776258
R4810 dcell_lv_0.bb[9].n5 dcell_lv_0.bb[9].t8 230.155
R4811 dcell_lv_0.bb[9].n9 dcell_lv_0.bb[9].t12 230.155
R4812 dcell_lv_0.bb[9].n8 dcell_lv_0.bb[9].t5 229.369
R4813 dcell_lv_0.bb[9].n2 dcell_lv_0.bb[9].t7 212.081
R4814 dcell_lv_0.bb[9].n3 dcell_lv_0.bb[9].t10 212.081
R4815 dcell_lv_0.bb[9].n1 dcell_lv_0.bb[9].n0 208.965
R4816 dcell_lv_0.bb[9].n4 dcell_lv_0.bb[9].n3 186.001
R4817 dcell_lv_0.bb[9] dcell_lv_0.bb[9].n8 157.927
R4818 dcell_lv_0.bb[9].n5 dcell_lv_0.bb[9].t13 157.856
R4819 dcell_lv_0.bb[9].n9 dcell_lv_0.bb[9].t11 157.856
R4820 dcell_lv_0.bb[9].n8 dcell_lv_0.bb[9].t4 157.07
R4821 dcell_lv_0.bb[9].n6 dcell_lv_0.bb[9].n5 152
R4822 dcell_lv_0.bb[9].n10 dcell_lv_0.bb[9].n9 152
R4823 dcell_lv_0.bb[9].n2 dcell_lv_0.bb[9].t6 139.78
R4824 dcell_lv_0.bb[9].n3 dcell_lv_0.bb[9].t9 139.78
R4825 dcell_lv_0.bb[9] dcell_lv_0.bb[9].n16 96.8352
R4826 dcell_lv_0.bb[9].n3 dcell_lv_0.bb[9].n2 61.346
R4827 dcell_lv_0.bb[9].n12 dcell_lv_0.bb[9].n11 31.3499
R4828 dcell_lv_0.bb[9].n13 dcell_lv_0.bb[9].n12 29.8627
R4829 dcell_lv_0.bb[9].n0 dcell_lv_0.bb[9].t1 26.5955
R4830 dcell_lv_0.bb[9].n0 dcell_lv_0.bb[9].t3 26.5955
R4831 dcell_lv_0.bb[9].n16 dcell_lv_0.bb[9].t0 24.9236
R4832 dcell_lv_0.bb[9].n16 dcell_lv_0.bb[9].t2 24.9236
R4833 dcell_lv_0.bb[9].n7 dcell_lv_0.bb[9].n6 19.1764
R4834 dcell_lv_0.bb[9].n14 dcell_lv_0.bb[9] 12.5445
R4835 dcell_lv_0.bb[9].n15 dcell_lv_0.bb[9] 11.2645
R4836 dcell_lv_0.bb[9].n11 dcell_lv_0.bb[9] 11.0938
R4837 dcell_lv_0.bb[9].n11 dcell_lv_0.bb[9].n10 9.9845
R4838 dcell_lv_0.bb[9].n14 dcell_lv_0.bb[9].n13 9.65467
R4839 dcell_lv_0.bb[9].n13 dcell_lv_0.bb[9].n4 9.30258
R4840 dcell_lv_0.bb[9].n15 dcell_lv_0.bb[9] 6.1445
R4841 dcell_lv_0.bb[9] dcell_lv_0.bb[9].n14 4.8645
R4842 dcell_lv_0.bb[9] dcell_lv_0.bb[9].n15 4.65505
R4843 dcell_lv_0.bb[9].n4 dcell_lv_0.bb[9] 3.0725
R4844 dcell_lv_0.bb[9].n10 dcell_lv_0.bb[9] 2.3045
R4845 dcell_lv_0.bb[9].n12 dcell_lv_0.bb[9].n7 2.24073
R4846 dcell_lv_0.bb[9].n6 dcell_lv_0.bb[9] 2.10199
R4847 dcell_lv_0.bb[9] dcell_lv_0.bb[9].n1 2.0485
R4848 dcell_lv_0.bb[9].n1 dcell_lv_0.bb[9] 1.55202
R4849 dcell_lv_0.bb[9].n7 dcell_lv_0.bb[9] 0.482922
R4850 a_6866_n660.t0 a_6866_n660.t1 49.8467
R4851 dcell_lv_0.b[9].n2 dcell_lv_0.b[9].t9 231.017
R4852 dcell_lv_0.b[9].n15 dcell_lv_0.b[9].t13 230.155
R4853 dcell_lv_0.b[9].n5 dcell_lv_0.b[9].t8 229.369
R4854 dcell_lv_0.b[9].n9 dcell_lv_0.b[9].t12 229.369
R4855 dcell_lv_0.b[9].n14 dcell_lv_0.b[9].t4 229.369
R4856 dcell_lv_0.b[9].n12 dcell_lv_0.b[9].t17 229.369
R4857 dcell_lv_0.b[9].n3 dcell_lv_0.b[9].t7 228.649
R4858 dcell_lv_0.b[9].n22 dcell_lv_0.b[9].n21 208.964
R4859 dcell_lv_0.b[9].n2 dcell_lv_0.b[9].t16 158.716
R4860 dcell_lv_0.b[9] dcell_lv_0.b[9].n14 157.927
R4861 dcell_lv_0.b[9].n15 dcell_lv_0.b[9].t5 157.856
R4862 dcell_lv_0.b[9].n5 dcell_lv_0.b[9].t15 157.07
R4863 dcell_lv_0.b[9].n9 dcell_lv_0.b[9].t11 157.07
R4864 dcell_lv_0.b[9].n14 dcell_lv_0.b[9].t10 157.07
R4865 dcell_lv_0.b[9].n12 dcell_lv_0.b[9].t6 157.07
R4866 dcell_lv_0.b[9].n3 dcell_lv_0.b[9].t14 156.35
R4867 dcell_lv_0.b[9] dcell_lv_0.b[9].n2 156.268
R4868 dcell_lv_0.b[9].n6 dcell_lv_0.b[9].n5 153.423
R4869 dcell_lv_0.b[9].n10 dcell_lv_0.b[9].n9 152
R4870 dcell_lv_0.b[9].n16 dcell_lv_0.b[9].n15 152
R4871 dcell_lv_0.b[9].n13 dcell_lv_0.b[9].n12 152
R4872 dcell_lv_0.b[9].n4 dcell_lv_0.b[9].n3 152
R4873 dcell_lv_0.b[9] dcell_lv_0.b[9].n0 96.8352
R4874 dcell_lv_0.b[9].n4 dcell_lv_0.b[9] 53.8309
R4875 dcell_lv_0.b[9].n20 dcell_lv_0.b[9].n19 43.993
R4876 dcell_lv_0.b[9].n21 dcell_lv_0.b[9].t1 26.5955
R4877 dcell_lv_0.b[9].n21 dcell_lv_0.b[9].t0 26.5955
R4878 dcell_lv_0.b[9].n0 dcell_lv_0.b[9].t3 24.9236
R4879 dcell_lv_0.b[9].n0 dcell_lv_0.b[9].t2 24.9236
R4880 dcell_lv_0.b[9].n11 dcell_lv_0.b[9].n10 18.4368
R4881 dcell_lv_0.b[9].n8 dcell_lv_0.b[9].n4 16.4183
R4882 dcell_lv_0.b[9].n7 dcell_lv_0.b[9].n6 14.4998
R4883 dcell_lv_0.b[9].n17 dcell_lv_0.b[9].n16 13.1513
R4884 dcell_lv_0.b[9] dcell_lv_0.b[9].n20 13.0565
R4885 dcell_lv_0.b[9].n18 dcell_lv_0.b[9].n13 11.8414
R4886 dcell_lv_0.b[9] dcell_lv_0.b[9].n1 11.2645
R4887 dcell_lv_0.b[9].n18 dcell_lv_0.b[9].n17 9.3005
R4888 dcell_lv_0.b[9].n17 dcell_lv_0.b[9] 7.11161
R4889 dcell_lv_0.b[9].n19 dcell_lv_0.b[9].n18 6.60324
R4890 dcell_lv_0.b[9].n1 dcell_lv_0.b[9] 6.1445
R4891 dcell_lv_0.b[9].n10 dcell_lv_0.b[9] 5.92643
R4892 dcell_lv_0.b[9].n1 dcell_lv_0.b[9] 4.65505
R4893 dcell_lv_0.b[9].n6 dcell_lv_0.b[9] 4.5042
R4894 dcell_lv_0.b[9].n13 dcell_lv_0.b[9] 4.39453
R4895 dcell_lv_0.b[9].n20 dcell_lv_0.b[9] 4.3525
R4896 dcell_lv_0.b[9].n16 dcell_lv_0.b[9] 2.3045
R4897 dcell_lv_0.b[9].n22 dcell_lv_0.b[9] 2.0485
R4898 dcell_lv_0.b[9] dcell_lv_0.b[9].n22 1.55202
R4899 dcell_lv_0.b[9].n4 dcell_lv_0.b[9] 1.43334
R4900 dcell_lv_0.b[9].n11 dcell_lv_0.b[9].n8 1.13136
R4901 dcell_lv_0.b[9].n8 dcell_lv_0.b[9].n7 1.10597
R4902 dcell_lv_0.b[9] dcell_lv_0.b[9].n11 0.434094
R4903 dcell_lv_0.b[9].n7 dcell_lv_0.b[9] 0.412609
R4904 dcell_lv_0.b[9].n19 dcell_lv_0.b[9] 0.266125
R4905 dcell_lv_0.logic_shift_seg2_0.x4.B.t0 dcell_lv_0.logic_shift_seg2_0.x4.B 272.038
R4906 dcell_lv_0.logic_shift_seg2_0.x4.B.n4 dcell_lv_0.logic_shift_seg2_0.x4.B.t0 258.846
R4907 dcell_lv_0.logic_shift_seg2_0.x4.B.n1 dcell_lv_0.logic_shift_seg2_0.x4.B.t4 241.536
R4908 dcell_lv_0.logic_shift_seg2_0.x4.B.n3 dcell_lv_0.logic_shift_seg2_0.x4.B.n0 195.704
R4909 dcell_lv_0.logic_shift_seg2_0.x4.B.n1 dcell_lv_0.logic_shift_seg2_0.x4.B.t3 169.237
R4910 dcell_lv_0.logic_shift_seg2_0.x4.B.n2 dcell_lv_0.logic_shift_seg2_0.x4.B.n1 154.514
R4911 dcell_lv_0.logic_shift_seg2_0.x4.B dcell_lv_0.logic_shift_seg2_0.x4.B.n3 29.0733
R4912 dcell_lv_0.logic_shift_seg2_0.x4.B.n0 dcell_lv_0.logic_shift_seg2_0.x4.B.t1 26.5955
R4913 dcell_lv_0.logic_shift_seg2_0.x4.B.n0 dcell_lv_0.logic_shift_seg2_0.x4.B.t2 26.5955
R4914 dcell_lv_0.logic_shift_seg2_0.x4.B.n3 dcell_lv_0.logic_shift_seg2_0.x4.B.n2 25.6543
R4915 dcell_lv_0.logic_shift_seg2_0.x4.B.n5 dcell_lv_0.logic_shift_seg2_0.x4.B 3.76521
R4916 dcell_lv_0.logic_shift_seg2_0.x4.B.n5 dcell_lv_0.logic_shift_seg2_0.x4.B.n4 3.03935
R4917 dcell_lv_0.logic_shift_seg2_0.x4.B.n4 dcell_lv_0.logic_shift_seg2_0.x4.B 2.30266
R4918 dcell_lv_0.logic_shift_seg2_0.x4.B dcell_lv_0.logic_shift_seg2_0.x4.B.n5 0.921363
R4919 dcell_lv_0.logic_shift_seg2_0.x4.B.n2 dcell_lv_0.logic_shift_seg2_0.x4.B 0.229071
R4920 decoder_3_0/decoder_2to4_2.bb[1].n1 decoder_3_0/decoder_2to4_2.bb[1].t3 230.155
R4921 decoder_3_0/decoder_2to4_2.bb[1].n0 decoder_3_0/decoder_2to4_2.bb[1].t5 229.369
R4922 decoder_3_0/decoder_2to4_2.bb[1].n4 decoder_3_0/decoder_2to4_2.bb[1].t1 221.538
R4923 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_2.bb[1].t0 162.351
R4924 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_2.bb[1].n0 157.927
R4925 decoder_3_0/decoder_2to4_2.bb[1].n1 decoder_3_0/decoder_2to4_2.bb[1].t2 157.856
R4926 decoder_3_0/decoder_2to4_2.bb[1].n0 decoder_3_0/decoder_2to4_2.bb[1].t4 157.07
R4927 decoder_3_0/decoder_2to4_2.bb[1].n2 decoder_3_0/decoder_2to4_2.bb[1].n1 152
R4928 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_2.bb[1].n3 24.6592
R4929 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_2.bb[1].n2 19.6746
R4930 decoder_3_0/decoder_2to4_2.bb[1].n4 decoder_3_0/decoder_2to4_2.bb[1] 17.3671
R4931 decoder_3_0/decoder_2to4_2.bb[1].n3 decoder_3_0/decoder_2to4_2.bb[1] 13.8127
R4932 decoder_3_0/decoder_2to4_2.bb[1].n5 decoder_3_0/decoder_2to4_2.bb[1] 11.6875
R4933 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_2.bb[1].n4 8.98055
R4934 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_2.bb[1].n5 7.23528
R4935 decoder_3_0/decoder_2to4_2.bb[1].n5 decoder_3_0/decoder_2to4_2.bb[1] 5.04292
R4936 decoder_3_0/decoder_2to4_2.bb[1].n2 decoder_3_0/decoder_2to4_2.bb[1] 2.13383
R4937 decoder_3_0/decoder_2to4_2.bb[1].n3 decoder_3_0/decoder_2to4_2.bb[1] 0.717167
R4938 a_24288_n1428.t0 a_24288_n1428.t1 49.8467
R4939 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 593.154
R4940 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 272.038
R4941 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 258.846
R4942 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 224.778
R4943 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 26.5955
R4944 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 26.5955
R4945 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 18.824
R4946 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 6.77697
R4947 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n3 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 3.76521
R4948 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n3 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 3.03935
R4949 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 2.30266
R4950 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n3 0.921363
R4951 dec2[2].n3 dec2[2].t1 334.788
R4952 dec2[2].n1 dec2[2].n0 152
R4953 dec2[2].n5 dec2[2].t2 126.27
R4954 dec2[2].n5 dec2[2].t4 125.558
R4955 dec2[2].n4 dec2[2].t5 121.127
R4956 dec2[2].n0 dec2[2].t3 114.031
R4957 dec2[2].n3 dec2[2].t0 87.8063
R4958 dec2[2].n0 dec2[2].t6 81.5883
R4959 dec2[2].n2 dec2[2] 15.1338
R4960 dec2[2] dec2[2].n1 11.4706
R4961 dec2[2].n6 dec2[2].n5 5.73592
R4962 dec2[2] dec2[2].n6 5.388
R4963 dec2[2].n1 dec2[2] 4.48881
R4964 dec2[2] dec2[2].n2 1.02758
R4965 dec2[2].n2 dec2[2] 0.6505
R4966 dec2[2].n4 dec2[2].n3 0.322615
R4967 dec2[2].n6 dec2[2].n4 0.177583
R4968 a_21282_427.t0 a_21282_427.t1 65.941
R4969 a_21282_685.t0 a_21282_685.t1 65.941
R4970 DIN2.n0 DIN2.t3 212.081
R4971 DIN2.n1 DIN2.t1 212.081
R4972 DIN2.n2 DIN2.n1 183.185
R4973 DIN2.n0 DIN2.t2 139.78
R4974 DIN2.n1 DIN2.t0 139.78
R4975 DIN2.n1 DIN2.n0 61.346
R4976 DIN2.n3 DIN2.n2 9.30224
R4977 DIN2.n2 DIN2 5.8885
R4978 DIN2.n3 DIN2 5.1005
R4979 DIN2 DIN2.n3 0.0525833
R4980 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t3 732.662
R4981 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 593.34
R4982 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n7 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 289.24
R4983 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t4 230.576
R4984 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t5 158.275
R4985 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 152
R4986 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n6 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 147.262
R4987 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n7 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n6 29.5774
R4988 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t2 26.5955
R4989 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t1 24.9236
R4990 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t0 24.9236
R4991 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 21.096
R4992 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 18.0633
R4993 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n7 11.3699
R4994 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 10.6891
R4995 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n6 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 10.3005
R4996 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 6.66717
R4997 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.0400833
R4998 a_13384_n1619.t0 a_13384_n1619.t1 114.052
R4999 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 593.154
R5000 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n3 224.776
R5001 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 132.067
R5002 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n3 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 26.5955
R5003 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n3 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 26.5955
R5004 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 18.824
R5005 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 6.77697
R5006 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 4.15748
R5007 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 3.76521
R5008 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 1.17559
R5009 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.921363
R5010 a_22669_n395.t0 a_22669_n395.t1 129.28
R5011 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n4 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t0 268.077
R5012 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n4 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t0 258.846
R5013 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n1 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t4 241.536
R5014 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n3 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n0 227.412
R5015 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n1 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t3 169.237
R5016 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n2 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n1 155.103
R5017 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n3 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n2 30.9223
R5018 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n0 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t1 26.5955
R5019 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n0 dcell_lv_0.seg_selector_logic_0.x2/x4.C.t2 26.5955
R5020 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n5 dcell_lv_0.seg_selector_logic_0.x2/x4.C 16.5652
R5021 dcell_lv_0.seg_selector_logic_0.x2/x4.C dcell_lv_0.seg_selector_logic_0.x2/x4.C.n3 10.1652
R5022 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n5 dcell_lv_0.seg_selector_logic_0.x2/x4.C 9.03579
R5023 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n5 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n4 8.8386
R5024 dcell_lv_0.seg_selector_logic_0.x2/x4.C.n2 dcell_lv_0.seg_selector_logic_0.x2/x4.C 7.75808
R5025 dcell_lv_0.seg_selector_logic_0.x2/x4.C dcell_lv_0.seg_selector_logic_0.x2/x4.C.n5 1.72748
R5026 decoder_3_0/decoder_2to4_1.b[1].n9 decoder_3_0/decoder_2to4_1.b[1].t16 231.017
R5027 decoder_3_0/decoder_2to4_1.b[1].n15 decoder_3_0/decoder_2to4_1.b[1].t4 230.155
R5028 decoder_3_0/decoder_2to4_1.b[1].n3 decoder_3_0/decoder_2to4_1.b[1].t5 230.155
R5029 decoder_3_0/decoder_2to4_1.b[1].n6 decoder_3_0/decoder_2to4_1.b[1].t6 229.369
R5030 decoder_3_0/decoder_2to4_1.b[1].n12 decoder_3_0/decoder_2to4_1.b[1].t10 229.369
R5031 decoder_3_0/decoder_2to4_1.b[1].n18 decoder_3_0/decoder_2to4_1.b[1].t13 229.369
R5032 decoder_3_0/decoder_2to4_1.b[1].n2 decoder_3_0/decoder_2to4_1.b[1].t14 229.369
R5033 decoder_3_0/decoder_2to4_1.b[1].n24 decoder_3_0/decoder_2to4_1.b[1].n23 208.964
R5034 decoder_3_0/decoder_2to4_1.b[1].n9 decoder_3_0/decoder_2to4_1.b[1].t15 158.716
R5035 decoder_3_0/decoder_2to4_1.b[1] decoder_3_0/decoder_2to4_1.b[1].n2 157.927
R5036 decoder_3_0/decoder_2to4_1.b[1].n15 decoder_3_0/decoder_2to4_1.b[1].t11 157.856
R5037 decoder_3_0/decoder_2to4_1.b[1].n3 decoder_3_0/decoder_2to4_1.b[1].t17 157.856
R5038 decoder_3_0/decoder_2to4_1.b[1].n6 decoder_3_0/decoder_2to4_1.b[1].t12 157.07
R5039 decoder_3_0/decoder_2to4_1.b[1].n12 decoder_3_0/decoder_2to4_1.b[1].t9 157.07
R5040 decoder_3_0/decoder_2to4_1.b[1].n18 decoder_3_0/decoder_2to4_1.b[1].t8 157.07
R5041 decoder_3_0/decoder_2to4_1.b[1].n2 decoder_3_0/decoder_2to4_1.b[1].t7 157.07
R5042 decoder_3_0/decoder_2to4_1.b[1].n7 decoder_3_0/decoder_2to4_1.b[1].n6 152.475
R5043 decoder_3_0/decoder_2to4_1.b[1].n19 decoder_3_0/decoder_2to4_1.b[1].n18 152.238
R5044 decoder_3_0/decoder_2to4_1.b[1].n10 decoder_3_0/decoder_2to4_1.b[1].n9 152
R5045 decoder_3_0/decoder_2to4_1.b[1].n13 decoder_3_0/decoder_2to4_1.b[1].n12 152
R5046 decoder_3_0/decoder_2to4_1.b[1].n16 decoder_3_0/decoder_2to4_1.b[1].n15 152
R5047 decoder_3_0/decoder_2to4_1.b[1].n4 decoder_3_0/decoder_2to4_1.b[1].n3 152
R5048 decoder_3_0/decoder_2to4_1.b[1] decoder_3_0/decoder_2to4_1.b[1].n0 96.8352
R5049 decoder_3_0/decoder_2to4_1.b[1].n23 decoder_3_0/decoder_2to4_1.b[1].t1 26.5955
R5050 decoder_3_0/decoder_2to4_1.b[1].n23 decoder_3_0/decoder_2to4_1.b[1].t0 26.5955
R5051 decoder_3_0/decoder_2to4_1.b[1].n21 decoder_3_0/decoder_2to4_1.b[1] 24.9713
R5052 decoder_3_0/decoder_2to4_1.b[1].n0 decoder_3_0/decoder_2to4_1.b[1].t3 24.9236
R5053 decoder_3_0/decoder_2to4_1.b[1].n0 decoder_3_0/decoder_2to4_1.b[1].t2 24.9236
R5054 decoder_3_0/decoder_2to4_1.b[1].n21 decoder_3_0/decoder_2to4_1.b[1].n20 23.8264
R5055 decoder_3_0/decoder_2to4_1.b[1].n22 decoder_3_0/decoder_2to4_1.b[1].n21 21.9086
R5056 decoder_3_0/decoder_2to4_1.b[1].n14 decoder_3_0/decoder_2to4_1.b[1].n13 20.0229
R5057 decoder_3_0/decoder_2to4_1.b[1].n17 decoder_3_0/decoder_2to4_1.b[1].n16 19.8154
R5058 decoder_3_0/decoder_2to4_1.b[1].n8 decoder_3_0/decoder_2to4_1.b[1].n7 17.1938
R5059 decoder_3_0/decoder_2to4_1.b[1].n11 decoder_3_0/decoder_2to4_1.b[1].n10 15.9118
R5060 decoder_3_0/decoder_2to4_1.b[1].n20 decoder_3_0/decoder_2to4_1.b[1].n19 15.7596
R5061 decoder_3_0/decoder_2to4_1.b[1] decoder_3_0/decoder_2to4_1.b[1].n5 14.5363
R5062 decoder_3_0/decoder_2to4_1.b[1] decoder_3_0/decoder_2to4_1.b[1].n22 13.0565
R5063 decoder_3_0/decoder_2to4_1.b[1].n5 decoder_3_0/decoder_2to4_1.b[1].n4 12.5635
R5064 decoder_3_0/decoder_2to4_1.b[1] decoder_3_0/decoder_2to4_1.b[1].n1 11.2645
R5065 decoder_3_0/decoder_2to4_1.b[1].n5 decoder_3_0/decoder_2to4_1.b[1] 7.11161
R5066 decoder_3_0/decoder_2to4_1.b[1].n1 decoder_3_0/decoder_2to4_1.b[1] 6.1445
R5067 decoder_3_0/decoder_2to4_1.b[1].n19 decoder_3_0/decoder_2to4_1.b[1] 5.68939
R5068 decoder_3_0/decoder_2to4_1.b[1].n7 decoder_3_0/decoder_2to4_1.b[1] 5.45235
R5069 decoder_3_0/decoder_2to4_1.b[1].n1 decoder_3_0/decoder_2to4_1.b[1] 4.65505
R5070 decoder_3_0/decoder_2to4_1.b[1].n16 decoder_3_0/decoder_2to4_1.b[1] 4.39453
R5071 decoder_3_0/decoder_2to4_1.b[1].n22 decoder_3_0/decoder_2to4_1.b[1] 4.3525
R5072 decoder_3_0/decoder_2to4_1.b[1].n10 decoder_3_0/decoder_2to4_1.b[1] 4.26717
R5073 decoder_3_0/decoder_2to4_1.b[1].n4 decoder_3_0/decoder_2to4_1.b[1] 2.13383
R5074 decoder_3_0/decoder_2to4_1.b[1].n13 decoder_3_0/decoder_2to4_1.b[1] 2.10199
R5075 decoder_3_0/decoder_2to4_1.b[1].n24 decoder_3_0/decoder_2to4_1.b[1] 2.0485
R5076 decoder_3_0/decoder_2to4_1.b[1] decoder_3_0/decoder_2to4_1.b[1].n24 1.55202
R5077 decoder_3_0/decoder_2to4_1.b[1].n20 decoder_3_0/decoder_2to4_1.b[1].n17 1.38917
R5078 decoder_3_0/decoder_2to4_1.b[1].n11 decoder_3_0/decoder_2to4_1.b[1].n8 1.30714
R5079 decoder_3_0/decoder_2to4_1.b[1].n14 decoder_3_0/decoder_2to4_1.b[1].n11 0.900891
R5080 decoder_3_0/decoder_2to4_1.b[1] decoder_3_0/decoder_2to4_1.b[1].n14 0.764172
R5081 decoder_3_0/decoder_2to4_1.b[1].n17 decoder_3_0/decoder_2to4_1.b[1] 0.15675
R5082 decoder_3_0/decoder_2to4_1.b[1].n8 decoder_3_0/decoder_2to4_1.b[1] 0.111828
R5083 dcell_lv_0.logic_shift_seg2_0.x4.C.n3 dcell_lv_0.logic_shift_seg2_0.x4.C.t4 230.363
R5084 dcell_lv_0.logic_shift_seg2_0.x4.C.n5 dcell_lv_0.logic_shift_seg2_0.x4.C.n2 203.147
R5085 dcell_lv_0.logic_shift_seg2_0.x4.C.n3 dcell_lv_0.logic_shift_seg2_0.x4.C.t3 158.064
R5086 dcell_lv_0.logic_shift_seg2_0.x4.C.n4 dcell_lv_0.logic_shift_seg2_0.x4.C.n3 156.364
R5087 dcell_lv_0.logic_shift_seg2_0.x4.C.n0 dcell_lv_0.logic_shift_seg2_0.x4.C.t1 132.067
R5088 dcell_lv_0.logic_shift_seg2_0.x4.C.n2 dcell_lv_0.logic_shift_seg2_0.x4.C.t0 26.5955
R5089 dcell_lv_0.logic_shift_seg2_0.x4.C.n2 dcell_lv_0.logic_shift_seg2_0.x4.C.t2 26.5955
R5090 dcell_lv_0.logic_shift_seg2_0.x4.C dcell_lv_0.logic_shift_seg2_0.x4.C.n5 21.6304
R5091 dcell_lv_0.logic_shift_seg2_0.x4.C.n5 dcell_lv_0.logic_shift_seg2_0.x4.C.n4 19.7021
R5092 dcell_lv_0.logic_shift_seg2_0.x4.C.n1 dcell_lv_0.logic_shift_seg2_0.x4.C.n0 4.15748
R5093 dcell_lv_0.logic_shift_seg2_0.x4.C dcell_lv_0.logic_shift_seg2_0.x4.C.n1 3.76521
R5094 dcell_lv_0.logic_shift_seg2_0.x4.C.n4 dcell_lv_0.logic_shift_seg2_0.x4.C 2.32777
R5095 dcell_lv_0.logic_shift_seg2_0.x4.C.n0 dcell_lv_0.logic_shift_seg2_0.x4.C 1.17559
R5096 dcell_lv_0.logic_shift_seg2_0.x4.C.n1 dcell_lv_0.logic_shift_seg2_0.x4.C 0.921363
R5097 a_7322_n884.t0 a_7322_n884.t1 49.8467
R5098 a_17078_n709.t0 a_17078_n709.t1 114.052
R5099 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t0 227.856
R5100 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n0 152.333
R5101 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t2 140.382
R5102 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t3 114.031
R5103 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t1 83.3993
R5104 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t4 81.5883
R5105 lvsf_7bit_0/lvsf_buff_7/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n1 14.4422
R5106 lvsf_7bit_0/lvsf_buff_7/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n3 7.56882
R5107 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n2 5.08175
R5108 lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_7/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R5109 a_20444_n199.t0 a_20444_n199.t1 55.3905
R5110 a_19848_n296.t0 a_19848_n296.n0 228.04
R5111 a_19848_n296.n0 a_19848_n296.t2 145.648
R5112 a_19848_n296.n0 a_19848_n296.t1 83.2159
R5113 dec1[2].n0 dec1[2].t1 334.788
R5114 dec1[2].n2 dec1[2].t2 126.27
R5115 dec1[2].n2 dec1[2].t3 125.558
R5116 dec1[2].n1 dec1[2].t4 121.127
R5117 dec1[2].n0 dec1[2].t0 87.8063
R5118 dec1[2].n3 dec1[2].n2 5.73592
R5119 dec1[2] dec1[2].n3 5.37342
R5120 dec1[2].n1 dec1[2].n0 0.322615
R5121 dec1[2].n3 dec1[2].n1 0.177583
R5122 a_22706_427.t0 a_22706_427.t1 65.941
R5123 a_22706_685.t0 a_22706_685.t1 65.941
R5124 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n1 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t0 227.856
R5125 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R5126 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n2 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t3 140.163
R5127 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n0 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t4 114.031
R5128 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n1 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t1 83.3993
R5129 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n0 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t2 81.5883
R5130 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n3 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R5131 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n3 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R5132 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R5133 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n2 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R5134 SH[2].n5 SH[2].n4 863.124
R5135 SH[2].n4 SH[2].n3 585
R5136 SH[2].n2 SH[2].t1 490.913
R5137 SH[2].n0 SH[2].t0 144.376
R5138 SH[2].n4 SH[2].t1 140.738
R5139 SH[2].n1 SH[2] 14.4526
R5140 SH[2].n1 SH[2] 13.9641
R5141 SH[2] SH[2].n0 11.3477
R5142 SH[2] SH[2].n2 11.2054
R5143 SH[2].n3 SH[2] 8.81089
R5144 SH[2] SH[2].n5 7.61955
R5145 SH[2].n5 SH[2] 4.98751
R5146 SH[2].n3 SH[2] 3.49141
R5147 SH[2].n0 SH[2] 2.94838
R5148 SH[2].n2 SH[2] 1.09557
R5149 SH[2] SH[2].n1 0.388379
R5150 a_25116_n1428.t0 a_25116_n1428.t1 49.8467
R5151 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 593.154
R5152 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 224.776
R5153 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 132.067
R5154 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 26.5955
R5155 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 26.5955
R5156 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 18.824
R5157 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 6.77697
R5158 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 4.15748
R5159 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 3.76521
R5160 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 1.17559
R5161 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.921363
R5162 a_14068_n199.t0 a_14068_n199.t1 55.3905
R5163 a_6406_n884.t0 a_6406_n884.t1 49.8467
R5164 dcell_lv_0.logic_shift_seg2_0.x4.A.n3 dcell_lv_0.logic_shift_seg2_0.x4.A.t4 232.214
R5165 dcell_lv_0.logic_shift_seg2_0.x4.A.n5 dcell_lv_0.logic_shift_seg2_0.x4.A.n2 191.1
R5166 dcell_lv_0.logic_shift_seg2_0.x4.A.n3 dcell_lv_0.logic_shift_seg2_0.x4.A.t3 159.915
R5167 dcell_lv_0.logic_shift_seg2_0.x4.A.n4 dcell_lv_0.logic_shift_seg2_0.x4.A.n3 155.097
R5168 dcell_lv_0.logic_shift_seg2_0.x4.A.n0 dcell_lv_0.logic_shift_seg2_0.x4.A.t2 132.067
R5169 dcell_lv_0.logic_shift_seg2_0.x4.A dcell_lv_0.logic_shift_seg2_0.x4.A.n5 33.6787
R5170 dcell_lv_0.logic_shift_seg2_0.x4.A.n5 dcell_lv_0.logic_shift_seg2_0.x4.A.n4 33.6331
R5171 dcell_lv_0.logic_shift_seg2_0.x4.A.n2 dcell_lv_0.logic_shift_seg2_0.x4.A.t1 26.5955
R5172 dcell_lv_0.logic_shift_seg2_0.x4.A.n2 dcell_lv_0.logic_shift_seg2_0.x4.A.t0 26.5955
R5173 dcell_lv_0.logic_shift_seg2_0.x4.A.n1 dcell_lv_0.logic_shift_seg2_0.x4.A.n0 4.15748
R5174 dcell_lv_0.logic_shift_seg2_0.x4.A dcell_lv_0.logic_shift_seg2_0.x4.A.n1 3.76521
R5175 dcell_lv_0.logic_shift_seg2_0.x4.A.n4 dcell_lv_0.logic_shift_seg2_0.x4.A 1.65211
R5176 dcell_lv_0.logic_shift_seg2_0.x4.A.n0 dcell_lv_0.logic_shift_seg2_0.x4.A 1.17559
R5177 dcell_lv_0.logic_shift_seg2_0.x4.A.n1 dcell_lv_0.logic_shift_seg2_0.x4.A 0.921363
R5178 a_21992_n1428.t0 a_21992_n1428.t1 49.8467
R5179 a_12128_n709.t0 a_12128_n709.t1 114.052
R5180 a_12524_n199.t0 a_12524_n199.t1 55.3905
R5181 a_18334_n1619.t0 a_18334_n1619.t1 114.052
R5182 a_17868_n296.t0 a_17868_n296.n0 228.04
R5183 a_17868_n296.n0 a_17868_n296.t2 145.648
R5184 a_17868_n296.n0 a_17868_n296.t1 83.2159
R5185 decoder_3_0/decoder_2to4_2.b[1].n10 decoder_3_0/decoder_2to4_2.b[1].t2 274.793
R5186 decoder_3_0/decoder_2to4_2.b[1].n5 decoder_3_0/decoder_2to4_2.b[1].t8 230.576
R5187 decoder_3_0/decoder_2to4_2.b[1].n1 decoder_3_0/decoder_2to4_2.b[1].t4 230.155
R5188 decoder_3_0/decoder_2to4_2.b[1].n0 decoder_3_0/decoder_2to4_2.b[1].t6 229.369
R5189 decoder_3_0/decoder_2to4_2.b[1].n10 decoder_3_0/decoder_2to4_2.b[1].n9 205.28
R5190 decoder_3_0/decoder_2to4_2.b[1].n5 decoder_3_0/decoder_2to4_2.b[1].t7 158.275
R5191 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_2.b[1].n0 157.927
R5192 decoder_3_0/decoder_2to4_2.b[1].n1 decoder_3_0/decoder_2to4_2.b[1].t9 157.856
R5193 decoder_3_0/decoder_2to4_2.b[1].n0 decoder_3_0/decoder_2to4_2.b[1].t5 157.07
R5194 decoder_3_0/decoder_2to4_2.b[1].n6 decoder_3_0/decoder_2to4_2.b[1].n5 153.067
R5195 decoder_3_0/decoder_2to4_2.b[1].n2 decoder_3_0/decoder_2to4_2.b[1].n1 152
R5196 decoder_3_0/decoder_2to4_2.b[1].n8 decoder_3_0/decoder_2to4_2.b[1].t3 133.124
R5197 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_2.b[1].n10 67.4857
R5198 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_2.b[1].n8 36.3299
R5199 decoder_3_0/decoder_2to4_2.b[1].n9 decoder_3_0/decoder_2to4_2.b[1].t0 26.5955
R5200 decoder_3_0/decoder_2to4_2.b[1].n9 decoder_3_0/decoder_2to4_2.b[1].t1 26.5955
R5201 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_2.b[1].n4 24.8883
R5202 decoder_3_0/decoder_2to4_2.b[1].n4 decoder_3_0/decoder_2to4_2.b[1].n3 13.8092
R5203 decoder_3_0/decoder_2to4_2.b[1].n3 decoder_3_0/decoder_2to4_2.b[1].n2 12.5635
R5204 decoder_3_0/decoder_2to4_2.b[1].n8 decoder_3_0/decoder_2to4_2.b[1].n7 10.6878
R5205 decoder_3_0/decoder_2to4_2.b[1].n7 decoder_3_0/decoder_2to4_2.b[1].n6 9.3005
R5206 decoder_3_0/decoder_2to4_2.b[1].n3 decoder_3_0/decoder_2to4_2.b[1] 7.11161
R5207 decoder_3_0/decoder_2to4_2.b[1].n7 decoder_3_0/decoder_2to4_2.b[1] 5.67507
R5208 decoder_3_0/decoder_2to4_2.b[1].n6 decoder_3_0/decoder_2to4_2.b[1] 5.6005
R5209 decoder_3_0/decoder_2to4_2.b[1].n2 decoder_3_0/decoder_2to4_2.b[1] 2.13383
R5210 decoder_3_0/decoder_2to4_2.b[1].n4 decoder_3_0/decoder_2to4_2.b[1] 0.727583
R5211 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 593.393
R5212 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 224.776
R5213 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 132.067
R5214 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 26.5955
R5215 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 26.5955
R5216 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 18.824
R5217 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 6.77697
R5218 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 4.15748
R5219 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 3.76521
R5220 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 1.17559
R5221 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.921363
R5222 a_12918_n296.t0 a_12918_n296.n0 228.04
R5223 a_12918_n296.n0 a_12918_n296.t2 145.648
R5224 a_12918_n296.n0 a_12918_n296.t1 83.2159
R5225 a_13078_n199.t0 a_13078_n199.t1 55.3905
R5226 a_7690_n1748.t0 a_7690_n1748.t1 49.8467
R5227 a_25142_n983.t0 a_25142_n983.t1 129.28
R5228 dec0[1].n0 dec0[1].t1 334.771
R5229 dec0[1].n3 dec0[1].t2 131.306
R5230 dec0[1].n1 dec0[1].t4 126.278
R5231 dec0[1].n1 dec0[1].t3 125.566
R5232 dec0[1].n0 dec0[1].t0 87.8231
R5233 dec0[1] dec0[1].n3 5.10467
R5234 dec0[1].n2 dec0[1].n1 4.68383
R5235 dec0[1].n2 dec0[1].n0 0.608192
R5236 dec0[1].n3 dec0[1].n2 0.177583
R5237 a_17474_n199.t0 a_17474_n199.t1 55.3905
R5238 dec2[0].n3 dec2[0].t0 334.771
R5239 dec2[0].n1 dec2[0].n0 152
R5240 dec2[0].n4 dec2[0].t3 126.278
R5241 dec2[0].n5 dec2[0].t5 125.566
R5242 dec2[0].n4 dec2[0].t6 125.566
R5243 dec2[0].n0 dec2[0].t2 114.031
R5244 dec2[0].n3 dec2[0].t1 87.8568
R5245 dec2[0].n0 dec2[0].t4 81.5883
R5246 dec2[0].n2 dec2[0] 15.6308
R5247 dec2[0] dec2[0].n1 11.4706
R5248 dec2[0] dec2[0].n6 5.04008
R5249 dec2[0].n6 dec2[0].n5 4.68383
R5250 dec2[0].n1 dec2[0] 4.48881
R5251 dec2[0] dec2[0].n2 1.01508
R5252 dec2[0].n6 dec2[0].n3 0.876942
R5253 dec2[0].n5 dec2[0].n4 0.713
R5254 dec2[0].n2 dec2[0] 0.6505
R5255 dec2b[0].n5 dec2b[0].n4 863.124
R5256 dec2b[0].n4 dec2b[0].n3 585
R5257 dec2b[0].n2 dec2b[0].t1 490.913
R5258 dec2b[0].n0 dec2b[0].t0 144.376
R5259 dec2b[0].n4 dec2b[0].t1 140.738
R5260 dec2b[0].n1 dec2b[0] 14.6401
R5261 dec2b[0].n1 dec2b[0] 13.9641
R5262 dec2b[0] dec2b[0].n0 11.3477
R5263 dec2b[0] dec2b[0].n2 11.2054
R5264 dec2b[0].n3 dec2b[0] 8.81089
R5265 dec2b[0] dec2b[0].n5 7.61955
R5266 dec2b[0].n5 dec2b[0] 4.98751
R5267 dec2b[0].n3 dec2b[0] 3.49141
R5268 dec2b[0].n0 dec2b[0] 2.94838
R5269 dec2b[0].n2 dec2b[0] 1.09557
R5270 dec2b[0] dec2b[0].n1 0.388379
R5271 a_22294_n983.t0 a_22294_n983.t1 129.28
R5272 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t1 227.856
R5273 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n0 152.333
R5274 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t2 140.382
R5275 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t3 114.031
R5276 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n2 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t0 83.3993
R5277 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n0 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t4 81.5883
R5278 lvsf_7bit_0/lvsf_buff_1/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n1 14.4422
R5279 lvsf_7bit_0/lvsf_buff_1/buff_hvl_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n3 7.56882
R5280 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n3 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n2 5.08175
R5281 lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n1 lvsf_7bit_0/lvsf_buff_1/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R5282 a_15494_n199.t0 a_15494_n199.t1 55.3905
R5283 a_14898_n296.n0 a_14898_n296.t1 228.04
R5284 a_14898_n296.n0 a_14898_n296.t2 145.648
R5285 a_14898_n296.t0 a_14898_n296.n0 83.2159
R5286 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n0 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t2 732.662
R5287 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n2 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t0 235.56
R5288 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n1 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t1 133.192
R5289 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n0 20.6511
R5290 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n1 19.6976
R5291 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n1 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 14.2962
R5292 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n2 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 2.22659
R5293 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n2 1.55202
R5294 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n0 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN 0.0400833
R5295 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n5 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n0 258.363
R5296 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n1 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t6 230.155
R5297 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n4 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n3 196.889
R5298 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n1 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t5 157.856
R5299 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n2 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n1 152
R5300 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n6 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t4 132.982
R5301 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n6 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n5 62.4946
R5302 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n3 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t3 32.5055
R5303 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n3 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t0 32.5055
R5304 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n4 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n2 30.2423
R5305 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n0 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t1 26.5955
R5306 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n0 dcell_lv_0.seg_selector_logic_0.x3/x3.A.t2 26.5955
R5307 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n5 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n4 5.2056
R5308 dcell_lv_0.seg_selector_logic_0.x3/x3.A dcell_lv_0.seg_selector_logic_0.x3/x3.A.n6 4.04261
R5309 dcell_lv_0.seg_selector_logic_0.x3/x3.A.n2 dcell_lv_0.seg_selector_logic_0.x3/x3.A 2.3045
R5310 a_7050_n884.t0 a_7050_n884.t1 49.8467
R5311 VBNDEC.n4 VBNDEC.t1 122.656
R5312 VBNDEC.n5 VBNDEC.t5 122.656
R5313 VBNDEC.n6 VBNDEC.t11 122.656
R5314 VBNDEC.n7 VBNDEC.t2 122.656
R5315 VBNDEC.n8 VBNDEC.t7 122.656
R5316 VBNDEC.n9 VBNDEC.t0 122.656
R5317 VBNDEC.n10 VBNDEC.t9 122.656
R5318 VBNDEC.n11 VBNDEC.t8 122.656
R5319 VBNDEC.n3 VBNDEC.t4 122.656
R5320 VBNDEC.n2 VBNDEC.t3 122.656
R5321 VBNDEC.n1 VBNDEC.t10 122.656
R5322 VBNDEC.n0 VBNDEC.t6 122.656
R5323 VBNDEC.n1 VBNDEC.n0 0.742167
R5324 VBNDEC.n2 VBNDEC.n1 0.742167
R5325 VBNDEC.n3 VBNDEC.n2 0.742167
R5326 VBNDEC.n11 VBNDEC.n10 0.742167
R5327 VBNDEC.n10 VBNDEC.n9 0.742167
R5328 VBNDEC.n9 VBNDEC.n8 0.742167
R5329 VBNDEC.n7 VBNDEC.n6 0.742167
R5330 VBNDEC.n6 VBNDEC.n5 0.742167
R5331 VBNDEC.n5 VBNDEC.n4 0.742167
R5332 VBNDEC VBNDEC.n11 0.652583
R5333 VBNDEC VBNDEC.n7 0.652583
R5334 VBNDEC.n0 VBNDEC 0.504667
R5335 VBNDEC VBNDEC.n3 0.0900833
R5336 VBNDEC.n8 VBNDEC 0.0900833
R5337 VBNDEC.n4 VBNDEC 0.0900833
R5338 a_23006_n983.t0 a_23006_n983.t1 129.28
R5339 dec1[1].n0 dec1[1].t1 334.771
R5340 dec1[1].n3 dec1[1].t4 131.306
R5341 dec1[1].n1 dec1[1].t2 126.278
R5342 dec1[1].n1 dec1[1].t3 125.566
R5343 dec1[1].n0 dec1[1].t0 87.8231
R5344 dec1[1] dec1[1].n3 5.10467
R5345 dec1[1].n2 dec1[1].n1 4.68383
R5346 dec1[1].n2 dec1[1].n0 0.608192
R5347 dec1[1].n3 dec1[1].n2 0.177583
R5348 a_18028_n199.t0 a_18028_n199.t1 55.3905
R5349 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n0 dcell_lv_0.seg_selector_logic_0.x4/x3.B.t3 230.363
R5350 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n3 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n2 201.161
R5351 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n0 dcell_lv_0.seg_selector_logic_0.x4/x3.B.t4 158.064
R5352 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n1 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n0 155.328
R5353 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n4 dcell_lv_0.seg_selector_logic_0.x4/x3.B.t2 140.53
R5354 dcell_lv_0.seg_selector_logic_0.x4/x3.B dcell_lv_0.seg_selector_logic_0.x4/x3.B.n3 36.416
R5355 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n3 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n1 29.1319
R5356 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n2 dcell_lv_0.seg_selector_logic_0.x4/x3.B.t1 26.5955
R5357 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n2 dcell_lv_0.seg_selector_logic_0.x4/x3.B.t0 26.5955
R5358 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n4 dcell_lv_0.seg_selector_logic_0.x4/x3.B 16.5652
R5359 dcell_lv_0.seg_selector_logic_0.x4/x3.B dcell_lv_0.seg_selector_logic_0.x4/x3.B.n4 9.03579
R5360 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n1 dcell_lv_0.seg_selector_logic_0.x4/x3.B 3.0725
R5361 dcell_lv_0.seg_selector_logic_0.x4/x3.B.n4 dcell_lv_0.seg_selector_logic_0.x4/x3.B 1.72748
R5362 a_24130_685.t0 a_24130_685.t1 65.941
R5363 a_24130_943.t0 a_24130_943.t1 65.941
R5364 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 593.393
R5365 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 272.038
R5366 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 258.846
R5367 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 224.778
R5368 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 26.5955
R5369 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 26.5955
R5370 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 18.824
R5371 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 6.77697
R5372 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 3.76521
R5373 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 3.03935
R5374 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 2.30266
R5375 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 0.921363
R5376 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 593.393
R5377 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 224.776
R5378 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 132.067
R5379 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 26.5955
R5380 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n3 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 26.5955
R5381 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 18.824
R5382 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 6.77697
R5383 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 4.15748
R5384 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 3.76521
R5385 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 1.17559
R5386 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.921363
R5387 a_21624_943.t0 a_21624_943.t1 65.941
R5388 a_7406_n884.t0 a_7406_n884.t1 60.9236
R5389 a_10414_n1619.t0 a_10414_n1619.t1 114.052
R5390 a_9948_n296.t0 a_9948_n296.n0 228.04
R5391 a_9948_n296.n0 a_9948_n296.t2 145.648
R5392 a_9948_n296.n0 a_9948_n296.t1 83.2159
R5393 dec2[1].n3 dec2[1].t1 334.771
R5394 dec2[1].n1 dec2[1].n0 152
R5395 dec2[1].n6 dec2[1].t4 131.306
R5396 dec2[1].n4 dec2[1].t3 126.278
R5397 dec2[1].n4 dec2[1].t2 125.566
R5398 dec2[1].n0 dec2[1].t5 114.031
R5399 dec2[1].n3 dec2[1].t0 87.8231
R5400 dec2[1].n0 dec2[1].t6 81.5883
R5401 dec2[1].n2 dec2[1] 14.6403
R5402 dec2[1] dec2[1].n1 11.4706
R5403 dec2[1] dec2[1].n6 5.12863
R5404 dec2[1].n5 dec2[1].n4 4.68383
R5405 dec2[1].n1 dec2[1] 4.48881
R5406 dec2[1] dec2[1].n2 1.01821
R5407 dec2[1].n2 dec2[1] 0.6505
R5408 dec2[1].n5 dec2[1].n3 0.608192
R5409 dec2[1].n6 dec2[1].n5 0.177583
R5410 a_21966_427.t0 a_21966_427.t1 65.941
R5411 a_21966_685.t0 a_21966_685.t1 65.941
R5412 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t4 732.773
R5413 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t8 212.081
R5414 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t6 212.081
R5415 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 208.965
R5416 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 186.001
R5417 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t7 139.78
R5418 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t5 139.78
R5419 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 96.8352
R5420 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 61.346
R5421 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t3 26.5955
R5422 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t2 26.5955
R5423 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t0 24.9236
R5424 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t1 24.9236
R5425 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 19.3172
R5426 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 12.5445
R5427 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 11.2645
R5428 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 9.65467
R5429 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 9.30258
R5430 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 6.1445
R5431 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 4.8645
R5432 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 4.65505
R5433 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 3.0725
R5434 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 2.0485
R5435 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 1.55202
R5436 a_16878_n296.t0 a_16878_n296.n0 228.04
R5437 a_16878_n296.n0 a_16878_n296.t2 145.648
R5438 a_16878_n296.n0 a_16878_n296.t1 83.2159
R5439 dec2[3].n3 dec2[3].t0 334.822
R5440 dec2[3].n1 dec2[3].n0 152
R5441 dec2[3].n4 dec2[3].t2 126.27
R5442 dec2[3].n4 dec2[3].t6 125.558
R5443 dec2[3].n5 dec2[3].t3 125.558
R5444 dec2[3].n0 dec2[3].t4 114.031
R5445 dec2[3].n3 dec2[3].t1 87.8063
R5446 dec2[3].n0 dec2[3].t5 81.5883
R5447 dec2[3].n2 dec2[3] 13.9702
R5448 dec2[3] dec2[3].n1 11.4706
R5449 dec2[3].n6 dec2[3].n5 5.73592
R5450 dec2[3] dec2[3].n6 5.66196
R5451 dec2[3].n1 dec2[3] 4.48881
R5452 dec2[3] dec2[3].n2 1.02238
R5453 dec2[3].n5 dec2[3].n4 0.713
R5454 dec2[3].n2 dec2[3] 0.6505
R5455 dec2[3].n6 dec2[3].n3 0.197295
R5456 a_6946_204.t0 a_6946_204.t1 49.8467
R5457 a_14108_n709.t0 a_14108_n709.t1 114.052
R5458 DIN5.n0 DIN5.t1 212.081
R5459 DIN5.n1 DIN5.t3 212.081
R5460 DIN5.n2 DIN5.n1 183.185
R5461 DIN5.n0 DIN5.t0 139.78
R5462 DIN5.n1 DIN5.t2 139.78
R5463 DIN5.n1 DIN5.n0 61.346
R5464 DIN5.n3 DIN5.n2 9.30224
R5465 DIN5.n2 DIN5 5.8885
R5466 DIN5.n3 DIN5 5.1005
R5467 DIN5 DIN5.n3 0.0525833
R5468 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n0 dcell_lv_0.seg_selector_logic_0.x2/x4.B.t4 241.536
R5469 dcell_lv_0.seg_selector_logic_0.x2/x4.B dcell_lv_0.seg_selector_logic_0.x2/x4.B.n3 237.577
R5470 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n0 dcell_lv_0.seg_selector_logic_0.x2/x4.B.t3 169.237
R5471 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n1 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n0 153.032
R5472 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n2 dcell_lv_0.seg_selector_logic_0.x2/x4.B.t2 131.691
R5473 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n2 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n1 32.8186
R5474 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n1 dcell_lv_0.seg_selector_logic_0.x2/x4.B 31.0244
R5475 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n3 dcell_lv_0.seg_selector_logic_0.x2/x4.B.t1 26.5955
R5476 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n3 dcell_lv_0.seg_selector_logic_0.x2/x4.B.t0 26.5955
R5477 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n4 dcell_lv_0.seg_selector_logic_0.x2/x4.B 16.5652
R5478 dcell_lv_0.seg_selector_logic_0.x2/x4.B dcell_lv_0.seg_selector_logic_0.x2/x4.B.n4 9.03579
R5479 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n4 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n2 8.8386
R5480 dcell_lv_0.seg_selector_logic_0.x2/x4.B.n4 dcell_lv_0.seg_selector_logic_0.x2/x4.B 1.72748
R5481 a_7682_n660.t0 a_7682_n660.t1 49.8467
R5482 a_7314_n660.t0 a_7314_n660.t1 60.9236
R5483 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n4 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t2 274.793
R5484 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n0 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t5 231.017
R5485 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n4 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n3 205.28
R5486 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n0 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t4 158.716
R5487 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n1 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n0 152.583
R5488 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n2 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t1 130.49
R5489 dcell_lv_0.seg_selector_logic_0.x2/x5.Y dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n4 67.4857
R5490 dcell_lv_0.seg_selector_logic_0.x2/x5.Y dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n2 38.9629
R5491 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n3 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t3 26.5955
R5492 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n3 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t0 26.5955
R5493 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n2 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n1 22.1046
R5494 dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n1 dcell_lv_0.seg_selector_logic_0.x2/x5.Y 3.68535
R5495 dec1[3].n0 dec1[3].t1 334.822
R5496 dec1[3].n1 dec1[3].t2 126.27
R5497 dec1[3].n1 dec1[3].t3 125.558
R5498 dec1[3].n2 dec1[3].t4 125.558
R5499 dec1[3].n0 dec1[3].t0 87.8063
R5500 dec1[3].n3 dec1[3].n2 5.73592
R5501 dec1[3] dec1[3].n3 5.64217
R5502 dec1[3].n2 dec1[3].n1 0.713
R5503 dec1[3].n3 dec1[3].n0 0.197295
R5504 a_21440_n1428.t0 a_21440_n1428.t1 49.8467
R5505 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 593.154
R5506 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 272.038
R5507 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 258.846
R5508 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 224.778
R5509 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 26.5955
R5510 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 26.5955
R5511 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 18.824
R5512 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 6.77697
R5513 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n3 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 3.76521
R5514 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n3 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 3.03935
R5515 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 2.30266
R5516 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n3 0.921363
R5517 a_15364_n1619.t0 a_15364_n1619.t1 114.052
R5518 bb[0].n4 bb[0].n3 863.124
R5519 bb[0].n3 bb[0].n2 585
R5520 bb[0].n1 bb[0].t1 490.913
R5521 bb[0].n7 bb[0].n6 152
R5522 bb[0].n0 bb[0].t0 144.376
R5523 bb[0].n3 bb[0].t1 140.738
R5524 bb[0].n6 bb[0].t2 114.031
R5525 bb[0].n6 bb[0].t3 81.5883
R5526 bb[0] bb[0].n7 16.7132
R5527 bb[0] bb[0].n5 13.7979
R5528 bb[0] bb[0].n0 11.3477
R5529 bb[0] bb[0].n1 11.2054
R5530 bb[0].n2 bb[0] 8.81089
R5531 bb[0] bb[0].n4 7.61955
R5532 bb[0].n5 bb[0] 7.17626
R5533 bb[0].n5 bb[0] 6.59444
R5534 bb[0].n4 bb[0] 4.98751
R5535 bb[0].n2 bb[0] 3.49141
R5536 bb[0].n0 bb[0] 2.94838
R5537 bb[0].n5 bb[0] 2.16154
R5538 bb[0].n7 bb[0] 1.16414
R5539 bb[0].n1 bb[0] 1.09557
R5540 b[0].n4 b[0].n3 863.124
R5541 b[0].n3 b[0].n2 585
R5542 b[0].n1 b[0].t1 490.913
R5543 b[0].n0 b[0].t0 144.376
R5544 b[0].n3 b[0].t1 140.738
R5545 b[0] b[0].n5 14.3755
R5546 b[0].n5 b[0] 13.5763
R5547 b[0] b[0].n0 11.3477
R5548 b[0] b[0].n1 11.2054
R5549 b[0].n2 b[0] 8.81089
R5550 b[0] b[0].n4 7.61955
R5551 b[0].n4 b[0] 4.98751
R5552 b[0].n2 b[0] 3.49141
R5553 b[0].n0 b[0] 2.94838
R5554 b[0].n1 b[0] 1.09557
R5555 b[0].n5 b[0] 0.776258
R5556 a_10108_n199.t0 a_10108_n199.t1 55.3905
R5557 a_7326_204.t0 a_7326_204.t1 49.8467
R5558 a_22308_685.t0 a_22308_685.t1 65.941
R5559 a_22308_943.t0 a_22308_943.t1 65.941
R5560 bb[1].n4 bb[1].n3 863.124
R5561 bb[1].n3 bb[1].n2 585
R5562 bb[1].n1 bb[1].t1 490.913
R5563 bb[1].n7 bb[1].n6 152
R5564 bb[1].n0 bb[1].t0 144.376
R5565 bb[1].n3 bb[1].t1 140.738
R5566 bb[1].n6 bb[1].t2 114.031
R5567 bb[1].n6 bb[1].t3 81.5883
R5568 bb[1] bb[1].n7 16.7132
R5569 bb[1] bb[1].n5 13.7979
R5570 bb[1] bb[1].n0 11.3477
R5571 bb[1] bb[1].n1 11.2054
R5572 bb[1].n2 bb[1] 8.81089
R5573 bb[1] bb[1].n4 7.61955
R5574 bb[1].n5 bb[1] 7.17626
R5575 bb[1].n5 bb[1] 6.59444
R5576 bb[1].n4 bb[1] 4.98751
R5577 bb[1].n2 bb[1] 3.49141
R5578 bb[1].n0 bb[1] 2.94838
R5579 bb[1].n5 bb[1] 2.16154
R5580 bb[1].n7 bb[1] 1.16414
R5581 bb[1].n1 bb[1] 1.09557
R5582 b[1].n4 b[1].n3 863.124
R5583 b[1].n3 b[1].n2 585
R5584 b[1].n1 b[1].t1 490.913
R5585 b[1].n0 b[1].t0 144.376
R5586 b[1].n3 b[1].t1 140.738
R5587 b[1] b[1].n5 14.3755
R5588 b[1].n5 b[1] 13.5763
R5589 b[1] b[1].n0 11.3477
R5590 b[1] b[1].n1 11.2054
R5591 b[1].n2 b[1] 8.81089
R5592 b[1] b[1].n4 7.61955
R5593 b[1].n4 b[1] 4.98751
R5594 b[1].n2 b[1] 3.49141
R5595 b[1].n0 b[1] 2.94838
R5596 b[1].n1 b[1] 1.09557
R5597 b[1].n5 b[1] 0.776258
R5598 a_23048_427.t0 a_23048_427.t1 65.941
R5599 a_23048_685.t0 a_23048_685.t1 65.941
R5600 a_21245_n395.t0 a_21245_n395.t1 129.28
R5601 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n1 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t0 268.077
R5602 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n1 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t0 258.846
R5603 dcell_lv_0.seg_selector_logic_0.x4/x3.A dcell_lv_0.seg_selector_logic_0.x4/x3.A.n0 237.577
R5604 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n2 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t3 231.835
R5605 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n2 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t4 157.07
R5606 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n3 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n2 152
R5607 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n0 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t1 26.5955
R5608 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n0 dcell_lv_0.seg_selector_logic_0.x4/x3.A.t2 26.5955
R5609 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n4 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n3 22.6473
R5610 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n5 dcell_lv_0.seg_selector_logic_0.x4/x3.A 16.5652
R5611 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n5 dcell_lv_0.seg_selector_logic_0.x4/x3.A 9.03579
R5612 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n5 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n4 8.0259
R5613 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n3 dcell_lv_0.seg_selector_logic_0.x4/x3.A 2.01193
R5614 dcell_lv_0.seg_selector_logic_0.x4/x3.A dcell_lv_0.seg_selector_logic_0.x4/x3.A.n5 1.72748
R5615 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n4 dcell_lv_0.seg_selector_logic_0.x4/x3.A.n1 0.813198
R5616 a_7598_n660.t0 a_7598_n660.t1 49.8467
R5617 a_23390_685.t0 a_23390_685.t1 65.941
R5618 a_23390_943.t0 a_23390_943.t1 65.941
R5619 a_18068_n709.t0 a_18068_n709.t1 114.052
R5620 a_22864_n1428.t0 a_22864_n1428.t1 49.8467
R5621 a_15058_n199.t0 a_15058_n199.t1 55.3905
R5622 a_24430_n983.t0 a_24430_n983.t1 129.28
R5623 a_6862_678.t0 a_6862_678.t1 41.3705
R5624 DIN1.n0 DIN1.t1 212.081
R5625 DIN1.n1 DIN1.t3 212.081
R5626 DIN1.n2 DIN1.n1 183.185
R5627 DIN1.n0 DIN1.t0 139.78
R5628 DIN1.n1 DIN1.t2 139.78
R5629 DIN1.n1 DIN1.n0 61.346
R5630 DIN1.n3 DIN1.n2 9.30224
R5631 DIN1.n2 DIN1 5.8885
R5632 DIN1.n3 DIN1 5.1005
R5633 DIN1 DIN1.n3 0.0525833
R5634 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t6 732.773
R5635 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t8 212.081
R5636 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t5 212.081
R5637 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 208.964
R5638 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 186.001
R5639 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t7 139.78
R5640 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t4 139.78
R5641 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 96.8352
R5642 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 61.346
R5643 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t1 26.5955
R5644 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t0 26.5955
R5645 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t3 24.9236
R5646 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t2 24.9236
R5647 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 24.588
R5648 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 12.5445
R5649 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 11.2645
R5650 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 9.65467
R5651 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 9.30258
R5652 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 6.1445
R5653 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 4.8645
R5654 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 4.65505
R5655 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 3.0725
R5656 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 2.0485
R5657 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 1.55202
R5658 dec0[0].n0 dec0[0].t0 334.771
R5659 dec0[0].n1 dec0[0].t3 126.278
R5660 dec0[0].n2 dec0[0].t4 125.566
R5661 dec0[0].n1 dec0[0].t2 125.566
R5662 dec0[0].n0 dec0[0].t1 87.8568
R5663 dec0[0] dec0[0].n3 5.013
R5664 dec0[0].n3 dec0[0].n2 4.68383
R5665 dec0[0].n3 dec0[0].n0 0.876942
R5666 dec0[0].n2 dec0[0].n1 0.713
R5667 a_24814_685.t0 a_24814_685.t1 65.941
R5668 a_24814_943.t0 a_24814_943.t1 65.941
R5669 a_13514_n199.t0 a_13514_n199.t1 55.3905
R5670 a_7774_n1748.t0 a_7774_n1748.t1 60.9236
R5671 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t2 732.662
R5672 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t0 233.621
R5673 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t1 152.889
R5674 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 26.8833
R5675 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 20.332
R5676 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n2 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 2.22659
R5677 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n2 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 1.93989
R5678 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n2 1.55202
R5679 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.110917
R5680 a_11534_n199.t0 a_11534_n199.t1 55.3905
R5681 a_10938_n296.t0 a_10938_n296.n0 228.04
R5682 a_10938_n296.n0 a_10938_n296.t2 145.648
R5683 a_10938_n296.n0 a_10938_n296.t1 83.2159
R5684 a_6406_n1748.t0 a_6406_n1748.t1 49.8467
R5685 a_21582_n983.t0 a_21582_n983.t1 129.28
R5686 a_23692_n1428.t0 a_23692_n1428.t1 49.8467
R5687 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t4 732.702
R5688 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 208.964
R5689 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 96.8352
R5690 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 30.179
R5691 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t1 26.5955
R5692 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t0 26.5955
R5693 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t3 24.9236
R5694 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t2 24.9236
R5695 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 13.0565
R5696 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 11.2645
R5697 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 6.1445
R5698 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 4.65505
R5699 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 4.3525
R5700 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 2.0485
R5701 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 1.55202
R5702 a_18464_n199.t0 a_18464_n199.t1 55.3905
R5703 dec2b[2].n4 dec2b[2].n3 863.124
R5704 dec2b[2].n3 dec2b[2].n2 585
R5705 dec2b[2].n1 dec2b[2].t1 490.913
R5706 dec2b[2].n0 dec2b[2].t0 144.376
R5707 dec2b[2].n3 dec2b[2].t1 140.738
R5708 dec2b[2] dec2b[2].n0 11.3477
R5709 dec2b[2] dec2b[2].n1 11.2054
R5710 dec2b[2].n2 dec2b[2] 8.81089
R5711 dec2b[2] dec2b[2].n4 7.61955
R5712 dec2b[2].n4 dec2b[2] 4.98751
R5713 dec2b[2].n2 dec2b[2] 3.49141
R5714 dec2b[2].n0 dec2b[2] 2.94838
R5715 dec2b[2].n1 dec2b[2] 1.09557
R5716 a_23732_427.t0 a_23732_427.t1 65.941
R5717 DIN9.n0 DIN9.t3 212.081
R5718 DIN9.n1 DIN9.t1 212.081
R5719 DIN9.n2 DIN9.n1 183.185
R5720 DIN9.n0 DIN9.t2 139.78
R5721 DIN9.n1 DIN9.t0 139.78
R5722 DIN9.n1 DIN9.n0 61.346
R5723 DIN9.n3 DIN9.n2 9.30224
R5724 DIN9.n2 DIN9 5.8885
R5725 DIN9.n3 DIN9 5.1005
R5726 DIN9 DIN9.n3 0.0525833
R5727 a_21624_685.t0 a_21624_685.t1 65.941
R5728 a_19018_n199.t0 a_19018_n199.t1 55.3905
R5729 dec2b[3].n4 dec2b[3].n3 863.124
R5730 dec2b[3].n3 dec2b[3].n2 585
R5731 dec2b[3].n1 dec2b[3].t1 490.913
R5732 dec2b[3].n0 dec2b[3].t0 144.376
R5733 dec2b[3].n3 dec2b[3].t1 140.738
R5734 dec2b[3] dec2b[3].n0 11.3477
R5735 dec2b[3] dec2b[3].n1 11.2054
R5736 dec2b[3].n2 dec2b[3] 8.81089
R5737 dec2b[3] dec2b[3].n4 7.61955
R5738 dec2b[3].n4 dec2b[3] 4.98751
R5739 dec2b[3].n2 dec2b[3] 3.49141
R5740 dec2b[3].n0 dec2b[3] 2.94838
R5741 dec2b[3].n1 dec2b[3] 1.09557
R5742 a_6682_n884.t0 a_6682_n884.t1 49.8467
R5743 a_11404_n1619.t0 a_11404_n1619.t1 114.052
R5744 bb[6].n4 bb[6].n3 863.124
R5745 bb[6].n3 bb[6].n2 585
R5746 bb[6].n1 bb[6].t1 490.913
R5747 bb[6].n7 bb[6].n6 152
R5748 bb[6].n0 bb[6].t0 144.376
R5749 bb[6].n3 bb[6].t1 140.738
R5750 bb[6].n6 bb[6].t2 114.031
R5751 bb[6].n6 bb[6].t3 81.5883
R5752 bb[6] bb[6].n7 16.7132
R5753 bb[6] bb[6].n5 13.7979
R5754 bb[6] bb[6].n0 11.3477
R5755 bb[6] bb[6].n1 11.2054
R5756 bb[6].n2 bb[6] 8.81089
R5757 bb[6] bb[6].n4 7.61955
R5758 bb[6].n5 bb[6] 7.17626
R5759 bb[6].n5 bb[6] 6.59444
R5760 bb[6].n4 bb[6] 4.98751
R5761 bb[6].n2 bb[6] 3.49141
R5762 bb[6].n0 bb[6] 2.94838
R5763 bb[6].n5 bb[6] 2.16154
R5764 bb[6].n7 bb[6] 1.16414
R5765 bb[6].n1 bb[6] 1.09557
R5766 b[6].n4 b[6].n3 863.124
R5767 b[6].n3 b[6].n2 585
R5768 b[6].n1 b[6].t1 490.913
R5769 b[6].n0 b[6].t0 144.376
R5770 b[6].n3 b[6].t1 140.738
R5771 b[6] b[6].n5 14.3755
R5772 b[6].n5 b[6] 13.5763
R5773 b[6] b[6].n0 11.3477
R5774 b[6] b[6].n1 11.2054
R5775 b[6].n2 b[6] 8.81089
R5776 b[6] b[6].n4 7.61955
R5777 b[6].n4 b[6] 4.98751
R5778 b[6].n2 b[6] 3.49141
R5779 b[6].n0 b[6] 2.94838
R5780 b[6].n1 b[6] 1.09557
R5781 b[6].n5 b[6] 0.776258
R5782 a_20314_n1619.t0 a_20314_n1619.t1 114.052
R5783 a_24472_943.t0 a_24472_943.t1 65.941
R5784 a_6590_n660.t0 a_6590_n660.t1 49.8467
R5785 a_16354_n1619.t0 a_16354_n1619.t1 114.052
R5786 a_7230_n660.t0 a_7230_n660.t1 49.8467
R5787 a_23140_n1428.t0 a_23140_n1428.t1 49.8467
R5788 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 593.163
R5789 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 272.038
R5790 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 258.846
R5791 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 224.778
R5792 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 26.5955
R5793 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 26.5955
R5794 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n3 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 3.76521
R5795 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 2.30266
R5796 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n3 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 2.0264
R5797 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n2 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 1.01345
R5798 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n3 0.921363
R5799 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 593.154
R5800 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 224.776
R5801 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 132.067
R5802 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 26.5955
R5803 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n3 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 26.5955
R5804 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 18.824
R5805 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 6.77697
R5806 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 4.15748
R5807 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 3.76521
R5808 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 1.17559
R5809 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.921363
R5810 a_23718_n983.t0 a_23718_n983.t1 129.28
R5811 a_11098_n199.t0 a_11098_n199.t1 55.3905
R5812 a_6590_428.t0 a_6590_428.t1 49.8467
R5813 a_20008_n199.t0 a_20008_n199.t1 55.3905
R5814 DIN8.n0 DIN8.t1 212.081
R5815 DIN8.n1 DIN8.t3 212.081
R5816 DIN8.n2 DIN8.n1 183.185
R5817 DIN8.n0 DIN8.t0 139.78
R5818 DIN8.n1 DIN8.t2 139.78
R5819 DIN8.n1 DIN8.n0 61.346
R5820 DIN8.n3 DIN8.n2 9.30224
R5821 DIN8.n2 DIN8 5.8885
R5822 DIN8.n3 DIN8 5.1005
R5823 DIN8 DIN8.n3 0.0525833
R5824 a_25156_685.t0 a_25156_685.t1 65.941
R5825 a_25156_943.t0 a_25156_943.t1 65.941
R5826 a_8058_678.t0 a_8058_678.t1 41.3705
R5827 a_19058_n709.t0 a_19058_n709.t1 114.052
R5828 a_24093_n395.t0 a_24093_n395.t1 129.28
R5829 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t4 732.702
R5830 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 208.964
R5831 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 96.8352
R5832 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 33.7628
R5833 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t0 26.5955
R5834 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t1 26.5955
R5835 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t2 24.9236
R5836 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t3 24.9236
R5837 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 13.0565
R5838 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 11.2645
R5839 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 6.1445
R5840 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 4.65505
R5841 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 4.3525
R5842 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 2.0485
R5843 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 1.55202
R5844 a_24564_n1428.t0 a_24564_n1428.t1 49.8467
R5845 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n1 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t0 227.856
R5846 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R5847 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n2 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t2 140.163
R5848 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n0 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t3 114.031
R5849 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n1 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t1 83.3993
R5850 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n0 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t4 81.5883
R5851 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n3 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R5852 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n3 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R5853 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R5854 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n2 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R5855 a_11928_n296.t0 a_11928_n296.n0 228.04
R5856 a_11928_n296.n0 a_11928_n296.t2 145.648
R5857 a_11928_n296.n0 a_11928_n296.t1 83.2159
R5858 a_6314_n660.t0 a_6314_n660.t1 49.8467
R5859 a_24130_427.t0 a_24130_427.t1 65.941
R5860 a_24805_n395.t0 a_24805_n395.t1 129.28
R5861 a_10148_n709.t0 a_10148_n709.t1 114.052
R5862 a_6314_428.t0 a_6314_428.t1 49.8467
R5863 a_6862_204.t0 a_6862_204.t1 49.8467
R5864 a_11138_n709.t0 a_11138_n709.t1 114.052
R5865 a_21957_n395.t0 a_21957_n395.t1 129.28
R5866 a_22268_n1428.t0 a_22268_n1428.t1 49.8467
R5867 a_12394_n1619.t0 a_12394_n1619.t1 114.052
R5868 DIN0.n0 DIN0.t3 212.081
R5869 DIN0.n1 DIN0.t1 212.081
R5870 DIN0.n2 DIN0.n1 183.185
R5871 DIN0.n0 DIN0.t2 139.78
R5872 DIN0.n1 DIN0.t0 139.78
R5873 DIN0.n1 DIN0.n0 61.346
R5874 DIN0.n3 DIN0.n2 9.30224
R5875 DIN0.n2 DIN0 5.8885
R5876 DIN0.n3 DIN0 5.1005
R5877 DIN0 DIN0.n3 0.0525833
R5878 a_21716_n1428.t0 a_21716_n1428.t1 49.8467
R5879 DIN4.n0 DIN4.t3 212.081
R5880 DIN4.n1 DIN4.t1 212.081
R5881 DIN4.n2 DIN4.n1 183.185
R5882 DIN4.n0 DIN4.t2 139.78
R5883 DIN4.n1 DIN4.t0 139.78
R5884 DIN4.n1 DIN4.n0 61.346
R5885 DIN4.n3 DIN4.n2 9.30224
R5886 DIN4.n2 DIN4 5.8885
R5887 DIN4.n3 DIN4 5.1005
R5888 DIN4 DIN4.n3 0.0525833
R5889 a_22308_427.t0 a_22308_427.t1 65.941
R5890 a_6478_204.t0 a_6478_204.t1 60.9236
R5891 a_6394_204.t0 a_6394_204.t1 49.8467
R5892 DIN7.n0 DIN7.t1 212.081
R5893 DIN7.n1 DIN7.t3 212.081
R5894 DIN7.n2 DIN7.n1 183.185
R5895 DIN7.n0 DIN7.t0 139.78
R5896 DIN7.n1 DIN7.t2 139.78
R5897 DIN7.n1 DIN7.n0 61.346
R5898 DIN7.n3 DIN7.n2 9.30224
R5899 DIN7.n2 DIN7 5.8885
R5900 DIN7.n3 DIN7 5.1005
R5901 DIN7 DIN7.n3 0.0525833
R5902 a_15098_n709.t0 a_15098_n709.t1 114.052
R5903 a_23390_427.t0 a_23390_427.t1 65.941
R5904 a_23381_n395.t0 a_23381_n395.t1 129.28
R5905 a_12088_n199.t0 a_12088_n199.t1 55.3905
R5906 a_10544_n199.t0 a_10544_n199.t1 55.3905
R5907 a_21282_943.t0 a_21282_943.t1 65.941
R5908 a_24814_427.t0 a_24814_427.t1 65.941
R5909 dec2b[1].n4 dec2b[1].n3 863.124
R5910 dec2b[1].n3 dec2b[1].n2 585
R5911 dec2b[1].n1 dec2b[1].t1 490.913
R5912 dec2b[1].n0 dec2b[1].t0 144.376
R5913 dec2b[1].n3 dec2b[1].t1 140.738
R5914 dec2b[1].n5 dec2b[1] 14.6422
R5915 dec2b[1].n5 dec2b[1] 14.1581
R5916 dec2b[1] dec2b[1].n0 11.3477
R5917 dec2b[1] dec2b[1].n1 11.2054
R5918 dec2b[1].n2 dec2b[1] 8.81089
R5919 dec2b[1] dec2b[1].n4 7.61955
R5920 dec2b[1].n4 dec2b[1] 4.98751
R5921 dec2b[1].n2 dec2b[1] 3.49141
R5922 dec2b[1].n0 dec2b[1] 2.94838
R5923 dec2b[1].n1 dec2b[1] 1.09557
R5924 dec2b[1] dec2b[1].n5 0.194439
R5925 a_6310_204.t0 a_6310_204.t1 49.8467
R5926 a_21966_943.t0 a_21966_943.t1 65.941
R5927 DIN3.n0 DIN3.t1 212.081
R5928 DIN3.n1 DIN3.t3 212.081
R5929 DIN3.n2 DIN3.n1 183.185
R5930 DIN3.n0 DIN3.t0 139.78
R5931 DIN3.n1 DIN3.t2 139.78
R5932 DIN3.n1 DIN3.n0 61.346
R5933 DIN3.n3 DIN3.n2 9.30224
R5934 DIN3.n2 DIN3 5.8885
R5935 DIN3.n3 DIN3 5.06092
R5936 DIN3 DIN3.n3 0.0525833
R5937 a_21624_427.t0 a_21624_427.t1 65.941
R5938 SH[3].n5 SH[3].n4 863.124
R5939 SH[3].n4 SH[3].n3 585
R5940 SH[3].n2 SH[3].t1 490.913
R5941 SH[3].n0 SH[3].t0 144.376
R5942 SH[3].n4 SH[3].t1 140.738
R5943 SH[3].n1 SH[3] 14.4526
R5944 SH[3].n1 SH[3] 13.9641
R5945 SH[3] SH[3].n0 11.3477
R5946 SH[3] SH[3].n2 11.2054
R5947 SH[3].n3 SH[3] 8.81089
R5948 SH[3] SH[3].n5 7.61955
R5949 SH[3].n5 SH[3] 4.98751
R5950 SH[3].n3 SH[3] 3.49141
R5951 SH[3].n0 SH[3] 2.94838
R5952 SH[3].n2 SH[3] 1.09557
R5953 SH[3] SH[3].n1 0.388379
R5954 SH[4].n5 SH[4].n4 863.124
R5955 SH[4].n4 SH[4].n3 585
R5956 SH[4].n2 SH[4].t1 490.913
R5957 SH[4].n0 SH[4].t0 144.376
R5958 SH[4].n4 SH[4].t1 140.738
R5959 SH[4].n1 SH[4] 14.4526
R5960 SH[4].n1 SH[4] 13.9641
R5961 SH[4] SH[4].n0 11.3477
R5962 SH[4] SH[4].n2 11.2054
R5963 SH[4].n3 SH[4] 8.81089
R5964 SH[4] SH[4].n5 7.61955
R5965 SH[4].n5 SH[4] 4.98751
R5966 SH[4].n3 SH[4] 3.49141
R5967 SH[4].n0 SH[4] 2.94838
R5968 SH[4].n2 SH[4] 1.09557
R5969 SH[4] SH[4].n1 0.388379
R5970 a_23048_943.t0 a_23048_943.t1 65.941
R5971 a_23416_n1428.t0 a_23416_n1428.t1 49.8467
C0 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN decoder_3_0/decoder_2to4_1.b[1] 0.07891f
C1 bb[3] b[3] 0.38613f
C2 decoder_3_0/decoder_2to4_2.bb[1] a_7980_n1212# 0.04364f
C3 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/decoder_2to4_1.bb[1] 0.07215f
C4 dcell_lv_0.seg_selector_logic_0.x3/x3.B lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.04268f
C5 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB dcell_lv_0.b[9] 0.09972f
C6 dcell_lv_0.seg_selector_logic_0.x3/x3.A dcell_lv_0.b[9] 0.1894f
C7 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/decoder_2to4_2.bb[0] 0.01833f
C8 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.06023f
C9 DIN4 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.17948f
C10 decoder_3_0/decoder_2to4_1.bb[1] dcell_lv_0.bb[9] 0.22976f
C11 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.07189f
C12 VBNLV lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.01121f
C13 DIN4 VDD 0.1713f
C14 DIN7 dcell_lv_0.b[8] 0.0349f
C15 bb[3] VDDH 0.59451f
C16 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB dcell_lv_0.bb[8] 0.13009f
C17 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB dcell_lv_0.bb[9] 0.4777f
C18 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[0] 0.14521f
C19 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.08402f
C20 DIN3 DIN2 0.0205f
C21 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.0673f
C22 dcell_lv_0.seg_selector_logic_0.x2/x4.A seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.26787f
C23 VDDH dec2b[1] 0.2927f
C24 bb[5] VBPLV 0.02136f
C25 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB decoder_3_0/decoder_2to4_1.b[1] 0.09158f
C26 dcell_lv_0.seg_selector_logic_0.x3/x3.A decoder_3_0/decoder_2to4_1.b[1] 0.01426f
C27 dcell_lv_0.seg_selector_logic_0.x2/x4.B VDD 0.25715f
C28 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.05681f
C29 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[0] 0.04293f
C30 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.06351f
C31 dcell_lv_0.logic_shift_seg2_0.x7.Y dcell_lv_0.b[8] 0.05396f
C32 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.09286f
C33 dcell_lv_0.seg_selector_logic_0.x4/x3.A VDD 0.32055f
C34 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.05086f
C35 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.32075f
C36 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN dcell_lv_0.bb[8] 0.14569f
C37 dcell_lv_0.seg_selector_logic_0.x4/x3.B dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.18203f
C38 dcell_lv_0.seg_selector_logic_0.x2/x4.A decoder_3_0/decoder_2to4_2.b[1] 0.01753f
C39 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN dcell_lv_0.bb[8] 0.04121f
C40 bb[2] VDDH 0.59451f
C41 decoder_3_0/decoder_2to4_2.b[0] lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.13258f
C42 decoder_3_0/decoder_2to4_2.b[0] VDD 1.23994f
C43 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.08793f
C44 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 8.33205f
C45 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN VDD 0.45123f
C46 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.07764f
C47 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.09277f
C48 dec2[0] VBPDEC 0.42415f
C49 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN dcell_lv_0.bb[9] 0.15563f
C50 dcell_lv_0.seg_selector_logic_0.x2/x4.B decoder_3_0/decoder_2to4_1.bb[1] 0.01119f
C51 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_2.bb[1] 0.04706f
C52 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN dcell_lv_0.b[8] 0.096f
C53 DIN5 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.17945f
C54 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 8.86068f
C55 bb[4] VBPLV 0.02136f
C56 dcell_lv_0.seg_selector_logic_0.x2/x4.B lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.02926f
C57 dcell_lv_0.seg_selector_logic_0.x2/x4.A dcell_lv_0.b[9] 0.08478f
C58 VBPLV bb[6] 0.02136f
C59 dcell_lv_0.seg_selector_logic_0.x3/x3.B lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.15193f
C60 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.13831f
C61 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB dcell_lv_0.bb[8] 0.13152f
C62 dcell_lv_0.bb[8] VDD 1.96294f
C63 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN decoder_3_0/decoder_2to4_2.bb[0] 0.0232f
C64 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.17262f
C65 dcell_lv_0.logic_shift_seg2_0.x8.Y VDD 0.41346f
C66 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.09544f
C67 decoder_3_0/decoder_2to4_2.bb[1] VDDH 0.19216f
C68 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.08566f
C69 b[3] VDDH 0.35752f
C70 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN dcell_lv_0.bb[9] 0.31523f
C71 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.08251f
C72 decoder_3_0/decoder_2to4_2.b[0] decoder_3_0/decoder_2to4_1.bb[1] 0.19158f
C73 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN decoder_3_0/decoder_2to4_1.bb[1] 0.08682f
C74 dcell_lv_0.seg_selector_logic_0.x3/x3.B seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 0.0651f
C75 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB dcell_lv_0.bb[9] 0.11469f
C76 dcell_lv_0.seg_selector_logic_0.x2/x4.A dcell_lv_0.logic_shift_seg2_0.x4.B 0.01088f
C77 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 1.70953f
C78 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.01148f
C79 decoder_3_0/decoder_2to4_2.b[0] lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.21931f
C80 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB dcell_lv_0.b[8] 0.09112f
C81 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.09125f
C82 dcell_lv_0.seg_selector_logic_0.x2/x4.A decoder_3_0/decoder_2to4_1.b[1] 0.04529f
C83 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C84 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN VDD 0.26425f
C85 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05095f
C86 dcell_lv_0.logic_shift_seg2_0.x6.Y VDD 0.28031f
C87 decoder_3_0/decoder_2to4_2.bb[0] dcell_lv_0.bb[9] 0.03366f
C88 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.12526f
C89 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN dcell_lv_0.bb[9] 0.02756f
C90 b[1] bb[1] 0.38613f
C91 bb[4] b[4] 0.38613f
C92 bb[3] VBPLV 0.02136f
C93 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.02359f
C94 dcell_lv_0.seg_selector_logic_0.x2/x4.A dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.01642f
C95 decoder_3_0/decoder_2to4_1.bb[1] dcell_lv_0.bb[8] 3.15778f
C96 dec2[3] VDDH 1.34981f
C97 dec2[2] dec2b[3] 0.136f
C98 dcell_lv_0.logic_shift_seg2_0.x8.Y decoder_3_0/decoder_2to4_1.bb[1] 0.18515f
C99 dcell_lv_0.bb[8] lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.60995f
C100 dcell_lv_0.seg_selector_logic_0.x2/x4.A dcell_lv_0.logic_shift_seg2_0.x4.C 0.01056f
C101 DIN9 DIN8 0.0205f
C102 dcell_lv_0.logic_shift_seg2_0.x8.Y lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.1019f
C103 dcell_lv_0.logic_shift_seg2_0.x4.A dcell_lv_0.b[8] 0.05306f
C104 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB VDD 0.31603f
C105 dcell_lv_0.b[8] dcell_lv_0.b[9] 2.90343f
C106 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.19088f
C107 VDD DIN0 0.1713f
C108 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.08636f
C109 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB VDD 0.63919f
C110 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD 0.2275f
C111 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 9.60185f
C112 DIN1 DIN0 0.0205f
C113 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.13238f
C114 DIN5 VDD 0.1713f
C115 dcell_lv_0.bb[9] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01428f
C116 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04786f
C117 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN decoder_3_0/decoder_2to4_1.bb[1] 0.04365f
C118 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/decoder_2to4_2.bb[1] 0.06435f
C119 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN VDD 0.55951f
C120 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.07407f
C121 dcell_lv_0.seg_selector_logic_0.x2/x4.B lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.04138f
C122 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[0] 0.13355f
C123 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.11368f
C124 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.08441f
C125 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 0.09351f
C126 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.04885f
C127 dcell_lv_0.b[8] decoder_3_0/decoder_2to4_1.b[1] 2.979f
C128 dec1[3] VDDH 0.93679f
C129 DIN6 DIN5 0.0205f
C130 bb[2] VBPLV 0.02136f
C131 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB decoder_3_0/decoder_2to4_1.bb[1] 0.06395f
C132 dec1[0] VDDH 0.82965f
C133 SH[4] seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.1675f
C134 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB decoder_3_0/decoder_2to4_1.bb[1] 0.07862f
C135 dcell_lv_0.seg_selector_logic_0.x2/x4.C dcell_lv_0.b[8] 0.0386f
C136 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.11522f
C137 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN dcell_lv_0.bb[8] 0.14193f
C138 dec2[0] dec2[2] 0.63138f
C139 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.08344f
C140 dec1[3] dec2[3] 0.07441f
C141 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.09478f
C142 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.10172f
C143 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.9653f
C144 decoder_3_0/decoder_2to4_2.b[0] lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.16722f
C145 decoder_3_0/decoder_2to4_1.bb[1] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.01978f
C146 VBNDEC dec2[1] 0.067f
C147 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB VDD 0.89562f
C148 DIN5 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.01586f
C149 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN dcell_lv_0.bb[9] 0.10655f
C150 dec1[0] dec2[3] 0.19105f
C151 VBNDEC dec1[1] 0.067f
C152 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.02523f
C153 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN dcell_lv_0.b[8] 0.08345f
C154 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[0] 0.07978f
C155 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB dcell_lv_0.bb[9] 0.10794f
C156 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.15699f
C157 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 8.29955f
C158 a_7980_n1490# dcell_lv_0.bb[8] 0.02963f
C159 VBPLV decoder_3_0/decoder_2to4_2.bb[1] 0.09601f
C160 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.30992f
C161 a_7980_n1490# dcell_lv_0.logic_shift_seg2_0.x8.Y 0.02202f
C162 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.12526f
C163 decoder_3_0/decoder_2to4_2.b[0] decoder_3_0/decoder_2to4_2.bb[0] 9.22813f
C164 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN decoder_3_0/decoder_2to4_2.bb[0] 0.02029f
C165 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[0] 0.0405f
C166 dcell_lv_0.bb[8] lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.23571f
C167 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 8.44169f
C168 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_2.b[0] 0.28496f
C169 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.05086f
C170 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN VDD 0.89921f
C171 VBPLV VDDH 11.3844f
C172 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB dcell_lv_0.bb[8] 0.10707f
C173 VBNLV seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.10895f
C174 VBNLV seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.91327f
C175 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN dcell_lv_0.b[9] 0.10073f
C176 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB dcell_lv_0.bb[9] 0.02209f
C177 dcell_lv_0.seg_selector_logic_0.x2/x5.Y dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.15447f
C178 dcell_lv_0.seg_selector_logic_0.x1/x3.B dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.13753f
C179 decoder_3_0/decoder_2to4_2.b[1] dcell_lv_0.bb[9] 0.01903f
C180 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB dcell_lv_0.bb[9] 0.09997f
C181 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB decoder_3_0/decoder_2to4_1.bb[1] 0.12539f
C182 dec0[0] VDDH 0.83181f
C183 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/decoder_2to4_2.bb[1] 0.05296f
C184 decoder_3_0/decoder_2to4_2.bb[0] dcell_lv_0.bb[8] 0.11989f
C185 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB dcell_lv_0.b[8] 0.09644f
C186 dcell_lv_0.logic_shift_seg2_0.x8.Y decoder_3_0/decoder_2to4_2.bb[0] 0.13705f
C187 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN dcell_lv_0.bb[8] 0.03532f
C188 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN VDD 0.46252f
C189 dcell_lv_0.seg_selector_logic_0.x3/x3.A dcell_lv_0.b[8] 0.19766f
C190 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.13661f
C191 dec1[3] dec1[0] 0.37541f
C192 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 8.31228f
C193 SH[3] seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.1675f
C194 dec0[3] VBNDEC 0.12185f
C195 dcell_lv_0.seg_selector_logic_0.x3/x3.B dcell_lv_0.b[9] 0.0191f
C196 decoder_3_0/decoder_2to4_2.b[0] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.04173f
C197 dcell_lv_0.logic_shift_seg2_0.x6.Y lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.04106f
C198 DIN7 dcell_lv_0.bb[8] 0.01582f
C199 bb[5] b[5] 0.38613f
C200 dcell_lv_0.logic_shift_seg2_0.x7.Y decoder_3_0/decoder_2to4_2.b[0] 0.08193f
C201 VBNDEC dec0[1] 0.067f
C202 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C203 VDDH VBPDEC 3.57436f
C204 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN decoder_3_0/decoder_2to4_1.b[1] 0.46012f
C205 dcell_lv_0.b[9] dcell_lv_0.bb[9] 11.5957f
C206 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN decoder_3_0/decoder_2to4_1.bb[1] 0.14241f
C207 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN decoder_3_0/decoder_2to4_2.bb[0] 0.08972f
C208 dcell_lv_0.seg_selector_logic_0.x2/x4.B seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 0.14577f
C209 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.22059f
C210 dcell_lv_0.bb[8] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01425f
C211 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB VDD 1.19512f
C212 b[4] VDDH 0.35752f
C213 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.08134f
C214 dec2[3] VBPDEC 0.18494f
C215 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.16804f
C216 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB DIN0 0.18007f
C217 VDD DIN1 0.1713f
C218 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN decoder_3_0/decoder_2to4_1.bb[1] 0.05032f
C219 dcell_lv_0.seg_selector_logic_0.x4/x3.B VDD 0.29366f
C220 DIN5 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.03498f
C221 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.09128f
C222 dcell_lv_0.logic_shift_seg2_0.x7.Y dcell_lv_0.logic_shift_seg2_0.x8.Y 0.01028f
C223 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.18829f
C224 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.03612f
C225 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB decoder_3_0/decoder_2to4_2.bb[0] 0.22756f
C226 dec0[2] VDDH 0.85277f
C227 decoder_3_0/decoder_2to4_1.b[1] dcell_lv_0.bb[9] 0.2026f
C228 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.72924f
C229 decoder_3_0/decoder_2to4_2.bb[0] lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.02032f
C230 DIN6 VDD 0.1713f
C231 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.01788f
C232 decoder_3_0/decoder_2to4_2.b[0] lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 0.07957f
C233 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB a_7980_n884# 0.02698f
C234 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB DIN2 0.01828f
C235 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 0.08837f
C236 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09291f
C237 dec1[3] dec0[0] 0.19105f
C238 dec0[3] dec0[1] 0.45254f
C239 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.6007f
C240 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.01851f
C241 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[0] 0.04718f
C242 VBNLV seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C243 dec1[2] dec2[1] 0.05012f
C244 SH[2] seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.1675f
C245 dcell_lv_0.seg_selector_logic_0.x2/x4.C dcell_lv_0.bb[9] 0.56698f
C246 decoder_3_0/decoder_2to4_2.bb[0] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.05346f
C247 dcell_lv_0.bb[9] dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.10418f
C248 dec1[1] dec1[2] 1.23984f
C249 VBNDEC dec1[2] 0.07829f
C250 DIN8 dcell_lv_0.bb[9] 0.01582f
C251 dcell_lv_0.logic_shift_seg2_0.x7.Y dcell_lv_0.logic_shift_seg2_0.x6.Y 0.29614f
C252 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB decoder_3_0/decoder_2to4_1.bb[1] 0.12627f
C253 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.09312f
C254 decoder_3_0/decoder_2to4_1.bb[1] VDD 2.59454f
C255 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.13636f
C256 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN dcell_lv_0.bb[8] 0.0975f
C257 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB VDD 3.59356f
C258 b[6] bb[6] 0.38613f
C259 dec1[3] VBPDEC 0.18454f
C260 dcell_lv_0.seg_selector_logic_0.x2/x4.A dcell_lv_0.b[8] 0.02039f
C261 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB dcell_lv_0.bb[8] 0.06022f
C262 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.47318f
C263 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[0] 0.04315f
C264 dcell_lv_0.seg_selector_logic_0.x2/x4.B dcell_lv_0.b[9] 0.01333f
C265 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 8.34443f
C266 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN dcell_lv_0.bb[9] 0.09511f
C267 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_2.b[0] 0.26566f
C268 dcell_lv_0.seg_selector_logic_0.x4/x3.A dcell_lv_0.b[9] 0.06751f
C269 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[0] 0.05752f
C270 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 0.09386f
C271 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 9.33133f
C272 DIN6 decoder_3_0/decoder_2to4_1.bb[1] 0.01584f
C273 dec1[0] VBPDEC 0.42417f
C274 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.09111f
C275 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD 0.23151f
C276 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01002f
C277 DIN6 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.17939f
C278 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 4.7892f
C279 b[0] VDDH 0.35752f
C280 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.06435f
C281 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB decoder_3_0/decoder_2to4_2.bb[0] 0.06296f
C282 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB 1.89276f
C283 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB dcell_lv_0.bb[8] 0.02716f
C284 dec0[3] dec1[2] 0.04526f
C285 dec1[3] dec0[2] 0.05726f
C286 dcell_lv_0.seg_selector_logic_0.x3/x3.B dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.28615f
C287 decoder_3_0/decoder_2to4_2.bb[1] dcell_lv_0.bb[9] 0.02906f
C288 decoder_3_0/decoder_2to4_2.b[1] dcell_lv_0.bb[8] 0.01841f
C289 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.15349f
C290 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB dcell_lv_0.bb[8] 0.09249f
C291 dcell_lv_0.seg_selector_logic_0.x2/x4.B decoder_3_0/decoder_2to4_1.b[1] 0.05972f
C292 decoder_3_0/decoder_2to4_2.b[0] dcell_lv_0.b[9] 0.2354f
C293 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN dcell_lv_0.b[9] 0.09202f
C294 decoder_3_0/decoder_2to4_1.bb[1] lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 4.05461f
C295 dcell_lv_0.seg_selector_logic_0.x4/x3.A decoder_3_0/decoder_2to4_1.b[1] 0.05552f
C296 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.09061f
C297 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB dcell_lv_0.bb[9] 0.11132f
C298 SH[1] seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.1675f
C299 dcell_lv_0.seg_selector_logic_0.x2/x4.A dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.0249f
C300 dcell_lv_0.seg_selector_logic_0.x2/x4.B dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.60657f
C301 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN VDD 0.7775f
C302 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 9.82456f
C303 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.09259f
C304 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.22947f
C305 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN decoder_3_0/decoder_2to4_2.bb[0] 0.07603f
C306 VBNLV seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C307 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB 1.2419f
C308 dec2[2] VDDH 1.28195f
C309 dcell_lv_0.bb[8] dcell_lv_0.b[9] 10.4407f
C310 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[1] 0.25101f
C311 dec0[0] VBPDEC 0.42417f
C312 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.09312f
C313 decoder_3_0/decoder_2to4_2.b[0] decoder_3_0/decoder_2to4_1.b[1] 0.1334f
C314 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN decoder_3_0/decoder_2to4_1.b[1] 0.08642f
C315 a_7980_n1490# VDD 0.03791f
C316 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN decoder_3_0/decoder_2to4_2.bb[0] 0.15048f
C317 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 0.02913f
C318 dec2[2] dec2[3] 1.06719f
C319 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.82224f
C320 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.13075f
C321 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN VDD 3.53121f
C322 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[1] 0.03899f
C323 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB DIN0 0.01622f
C324 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.0897f
C325 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C326 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.09111f
C327 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB VDD 0.66813f
C328 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.29968f
C329 dcell_lv_0.bb[8] decoder_3_0/decoder_2to4_1.b[1] 0.28897f
C330 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05095f
C331 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN decoder_3_0/decoder_2to4_1.bb[1] 0.13686f
C332 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.13238f
C333 dec0[0] dec0[2] 0.63006f
C334 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.1591f
C335 decoder_3_0/decoder_2to4_2.bb[0] lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.08388f
C336 decoder_3_0/decoder_2to4_2.b[0] lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09062f
C337 decoder_3_0/decoder_2to4_2.b[1] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.05677f
C338 decoder_3_0/decoder_2to4_2.bb[0] VDD 1.04528f
C339 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.0848f
C340 VDDH dec2b[2] 0.29298f
C341 VDD DIN2 0.1713f
C342 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN VDD 0.36208f
C343 dcell_lv_0.seg_selector_logic_0.x2/x4.C dcell_lv_0.bb[8] 0.01151f
C344 dcell_lv_0.bb[8] dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.06718f
C345 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 0.08957f
C346 dcell_lv_0.seg_selector_logic_0.x2/x5.Y dcell_lv_0.b[8] 0.10246f
C347 DIN8 dcell_lv_0.bb[8] 0.17935f
C348 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD 0.23023f
C349 DIN2 DIN1 0.0205f
C350 DIN7 VDD 0.1713f
C351 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB dcell_lv_0.b[9] 0.08386f
C352 a_7980_n1490# lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.01008f
C353 dec2[0] dec2[1] 1.3432f
C354 dec1[3] dec2[2] 0.04526f
C355 dec0[2] VBPDEC 0.19485f
C356 decoder_3_0/decoder_2to4_1.bb[1] lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.54465f
C357 dcell_lv_0.logic_shift_seg2_0.x6.Y decoder_3_0/decoder_2to4_1.b[1] 0.06271f
C358 decoder_3_0/decoder_2to4_2.bb[1] a_7980_n884# 0.01759f
C359 dec1[1] dec2[0] 0.05039f
C360 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN dcell_lv_0.bb[8] 0.08499f
C361 VBNDEC dec2[0] 0.06769f
C362 dcell_lv_0.seg_selector_logic_0.x2/x4.A dcell_lv_0.bb[9] 0.09623f
C363 b[5] VDDH 0.35752f
C364 decoder_3_0/decoder_2to4_2.b[0] decoder_3_0/decoder_2to4_2.bb[1] 0.21776f
C365 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 12.0047f
C366 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN dcell_lv_0.b[9] 0.01121f
C367 VBNLV seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C368 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB decoder_3_0/decoder_2to4_1.bb[1] 0.46395f
C369 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 0.0973f
C370 DIN9 dcell_lv_0.bb[9] 0.17935f
C371 VDD seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 1.25889f
C372 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.09009f
C373 DIN7 DIN6 0.0205f
C374 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[0] 0.10618f
C375 b[6] VDDH 0.21782f
C376 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 0.17015f
C377 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_1.bb[1] 0.11902f
C378 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[1] 0.01273f
C379 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.08118f
C380 dcell_lv_0.logic_shift_seg2_0.x7.Y VDD 0.33964f
C381 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN decoder_3_0/decoder_2to4_1.bb[1] 0.68564f
C382 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB decoder_3_0/decoder_2to4_1.b[1] 0.07852f
C383 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.28823f
C384 decoder_3_0/decoder_2to4_2.bb[0] lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.31211f
C385 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y decoder_3_0/decoder_2to4_1.b[1] 0.15076f
C386 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN dcell_lv_0.b[8] 0.09946f
C387 decoder_3_0/decoder_2to4_2.bb[1] dcell_lv_0.bb[8] 0.02834f
C388 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.07926f
C389 DIN7 decoder_3_0/decoder_2to4_1.bb[1] 0.17937f
C390 SH[4] VDDH 0.3346f
C391 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN 0.72875f
C392 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.09211f
C393 VBNLV lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.01349f
C394 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB dcell_lv_0.bb[8] 0.09836f
C395 dcell_lv_0.seg_selector_logic_0.x3/x3.B dcell_lv_0.b[8] 0.06214f
C396 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.02163f
C397 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[1] 0.01393f
C398 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB dcell_lv_0.b[9] 0.13022f
C399 VDDH bb[1] 0.59451f
C400 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.0888f
C401 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.10475f
C402 VBNLV decoder_3_0/decoder_2to4_2.bb[0] 0.01501f
C403 decoder_3_0/decoder_2to4_1.bb[1] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01445f
C404 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN decoder_3_0/decoder_2to4_2.bb[1] 0.0256f
C405 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 9.82232f
C406 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.11249f
C407 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.048f
C408 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN VDD 0.44141f
C409 dcell_lv_0.b[8] dcell_lv_0.bb[9] 0.10646f
C410 VBNDEC decoder_3_0/decoder_2to4_2.b[1] 0.01209f
C411 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.14053f
C412 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB 0.6219f
C413 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB VDD 0.51982f
C414 decoder_3_0/decoder_2to4_2.b[0] decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.18005f
C415 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[1] 0.14159f
C416 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB 0.09079f
C417 dcell_lv_0.seg_selector_logic_0.x2/x4.B dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.77374f
C418 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN DIN1 0.03521f
C419 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN dcell_lv_0.b[9] 0.14582f
C420 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB decoder_3_0/decoder_2to4_1.b[1] 0.12612f
C421 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB decoder_3_0/decoder_2to4_2.bb[1] 0.03132f
C422 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN decoder_3_0/decoder_2to4_2.bb[0] 0.08602f
C423 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD 0.21864f
C424 VBNLV seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01401f
C425 dec2[2] VBPDEC 0.19525f
C426 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05297f
C427 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB VDD 0.32717f
C428 decoder_3_0/decoder_2to4_2.b[1] lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.01895f
C429 decoder_3_0/decoder_2to4_2.b[1] VDD 1.57888f
C430 VDDH bb[0] 0.5944f
C431 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.09515f
C432 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.08961f
C433 decoder_3_0/decoder_2to4_2.bb[1] seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C434 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB VDD 0.64867f
C435 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD 0.23151f
C436 decoder_3_0/decoder_2to4_2.bb[1] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.26447f
C437 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN decoder_3_0/decoder_2to4_1.bb[1] 0.09178f
C438 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.09058f
C439 dec2[1] dec2b[1] 0.43405f
C440 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB decoder_3_0/decoder_2to4_1.bb[1] 0.07479f
C441 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN decoder_3_0/decoder_2to4_1.b[1] 0.14083f
C442 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.0962f
C443 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB DIN1 0.17975f
C444 dcell_lv_0.seg_selector_logic_0.x2/x5.Y dcell_lv_0.bb[9] 0.0184f
C445 dcell_lv_0.bb[9] dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.24146f
C446 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.18193f
C447 decoder_3_0/decoder_2to4_2.bb[0] lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.10438f
C448 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A VDDH 0.8236f
C449 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.07731f
C450 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN VDDH 0.19611f
C451 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB decoder_3_0/decoder_2to4_2.bb[0] 0.02445f
C452 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB dcell_lv_0.b[9] 0.13166f
C453 dcell_lv_0.logic_shift_seg2_0.x4.A VDD 1.0548f
C454 DIN4 DIN3 0.0205f
C455 dcell_lv_0.seg_selector_logic_0.x2/x4.A dcell_lv_0.bb[8] 0.18669f
C456 dcell_lv_0.b[9] VDD 1.60376f
C457 dcell_lv_0.seg_selector_logic_0.x2/x4.B dcell_lv_0.b[8] 0.01469f
C458 dcell_lv_0.seg_selector_logic_0.x4/x3.A dcell_lv_0.b[8] 0.15687f
C459 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB decoder_3_0/decoder_2to4_1.bb[1] 0.03508f
C460 a_7980_n1212# VDD 0.02571f
C461 dcell_lv_0.seg_selector_logic_0.x4/x3.B dcell_lv_0.b[9] 0.04039f
C462 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.1319f
C463 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN decoder_3_0/decoder_2to4_2.bb[0] 0.05327f
C464 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_1.bb[1] 0.02891f
C465 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB decoder_3_0/decoder_2to4_1.bb[1] 0.08705f
C466 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.16815f
C467 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.08451f
C468 a_7980_n1756# decoder_3_0/decoder_2to4_2.b[0] 0.01631f
C469 decoder_3_0/decoder_2to4_2.b[1] lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.04741f
C470 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.10315f
C471 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.06351f
C472 dcell_lv_0.logic_shift_seg2_0.x4.B VDD 0.36582f
C473 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 0.09845f
C474 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN dcell_lv_0.bb[9] 0.11097f
C475 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB decoder_3_0/decoder_2to4_1.b[1] 0.12629f
C476 decoder_3_0/decoder_2to4_1.b[1] VDD 1.81275f
C477 dcell_lv_0.logic_shift_seg2_0.x7.Y lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.20923f
C478 decoder_3_0/decoder_2to4_2.b[0] dcell_lv_0.b[8] 0.12874f
C479 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN dcell_lv_0.b[8] 0.09083f
C480 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 0.20842f
C481 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.05434f
C482 decoder_3_0/decoder_2to4_1.bb[1] dcell_lv_0.b[9] 0.11542f
C483 dcell_lv_0.seg_selector_logic_0.x4/x3.B decoder_3_0/decoder_2to4_1.b[1] 0.0979f
C484 VBPLV bb[1] 0.02136f
C485 decoder_3_0/decoder_2to4_2.bb[0] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.05506f
C486 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 2.40873f
C487 VBNLV decoder_3_0/decoder_2to4_2.b[1] 0.03924f
C488 dcell_lv_0.seg_selector_logic_0.x2/x4.C VDD 0.26021f
C489 a_7980_n1756# dcell_lv_0.logic_shift_seg2_0.x8.Y 0.01335f
C490 VDD dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.33616f
C491 SH[3] VDDH 0.33127f
C492 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB dcell_lv_0.b[9] 0.24589f
C493 DIN8 VDD 0.1713f
C494 decoder_3_0/decoder_2to4_2.bb[1] seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C495 dcell_lv_0.seg_selector_logic_0.x2/x4.B dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.04842f
C496 DIN6 decoder_3_0/decoder_2to4_1.b[1] 0.03492f
C497 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 0.16266f
C498 dcell_lv_0.logic_shift_seg2_0.x4.C VDD 0.33515f
C499 dcell_lv_0.bb[8] dcell_lv_0.b[8] 11.8247f
C500 VBNDEC decoder_3_0/decoder_2to4_2.bb[1] 0.06649f
C501 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN decoder_3_0/decoder_2to4_2.bb[1] 0.0811f
C502 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A VDDH 0.90722f
C503 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.15627f
C504 dec2[1] VDDH 1.2541f
C505 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN VDD 0.43649f
C506 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.09372f
C507 decoder_3_0/decoder_2to4_1.bb[1] decoder_3_0/decoder_2to4_1.b[1] 11.41f
C508 dec1[1] VDDH 0.82606f
C509 VBNDEC VDDH 0.33564f
C510 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[1] 0.0288f
C511 dcell_lv_0.logic_shift_seg2_0.x4.B lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.01229f
C512 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.08933f
C513 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.28825f
C514 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 0.09237f
C515 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB decoder_3_0/decoder_2to4_1.b[1] 10.545f
C516 dec2[0] dec2b[0] 0.43405f
C517 dec2[1] dec2[3] 0.45257f
C518 dcell_lv_0.seg_selector_logic_0.x2/x4.C decoder_3_0/decoder_2to4_1.bb[1] 0.02737f
C519 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.19474f
C520 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD 0.21766f
C521 decoder_3_0/decoder_2to4_1.bb[1] dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.14095f
C522 dcell_lv_0.logic_shift_seg2_0.x6.Y dcell_lv_0.b[8] 0.15123f
C523 VBPLV bb[0] 0.02136f
C524 decoder_3_0/decoder_2to4_2.bb[0] lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 0.02187f
C525 dec1[1] dec2[3] 0.05747f
C526 VBNDEC dec2[3] 0.12185f
C527 decoder_3_0/decoder_2to4_2.bb[1] VDD 0.48049f
C528 dcell_lv_0.seg_selector_logic_0.x2/x4.C lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.04593f
C529 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB decoder_3_0/decoder_2to4_2.bb[0] 0.12942f
C530 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.07209f
C531 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.48789f
C532 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_1.b[1] 0.10472f
C533 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 0.01148f
C534 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.21135f
C535 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN dcell_lv_0.b[9] 0.14205f
C536 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB VDD 0.64104f
C537 decoder_3_0/decoder_2to4_2.b[1] lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.02885f
C538 VBPLV seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.29407f
C539 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.2707f
C540 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN decoder_3_0/decoder_2to4_1.bb[1] 0.07915f
C541 dcell_lv_0.seg_selector_logic_0.x2/x5.Y dcell_lv_0.bb[8] 0.0239f
C542 dcell_lv_0.seg_selector_logic_0.x3/x3.A VDD 0.58965f
C543 VBPLV seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.02638f
C544 dcell_lv_0.bb[8] dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.09248f
C545 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB DIN1 0.01607f
C546 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.2094f
C547 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.08365f
C548 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB 0.09657f
C549 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB dcell_lv_0.b[8] 0.08269f
C550 dec0[3] VDDH 0.90345f
C551 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB decoder_3_0/decoder_2to4_2.bb[0] 0.05782f
C552 decoder_3_0/decoder_2to4_2.bb[1] seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C553 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 2.66992f
C554 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_2.bb[0] 2.8803f
C555 dec0[1] VDDH 0.82847f
C556 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB decoder_3_0/decoder_2to4_2.bb[0] 0.02029f
C557 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.02001f
C558 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.09702f
C559 dcell_lv_0.seg_selector_logic_0.x2/x4.B dcell_lv_0.bb[9] 0.22399f
C560 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[0] 0.07179f
C561 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[1] 0.18208f
C562 dec2[2] dec2b[2] 0.43405f
C563 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y decoder_3_0/decoder_2to4_2.b[1] 0.17953f
C564 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN decoder_3_0/decoder_2to4_1.b[1] 0.13647f
C565 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_1.bb[1] 0.02873f
C566 dcell_lv_0.logic_shift_seg2_0.x4.A lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.10863f
C567 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN dcell_lv_0.b[9] 0.69542f
C568 dec1[3] dec1[1] 0.45254f
C569 decoder_3_0/decoder_2to4_2.b[0] decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.16197f
C570 dec1[3] VBNDEC 0.12185f
C571 DIN3 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.17953f
C572 VBNLV lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.01074f
C573 decoder_3_0/decoder_2to4_2.bb[1] lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.04259f
C574 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A VDDH 0.90722f
C575 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB dcell_lv_0.b[9] 0.10397f
C576 b[1] VDDH 0.35752f
C577 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB decoder_3_0/decoder_2to4_1.bb[1] 0.09197f
C578 dec1[1] dec1[0] 1.25358f
C579 VBNDEC dec1[0] 0.06769f
C580 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN dcell_lv_0.bb[8] 0.10061f
C581 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.09623f
C582 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD 0.21618f
C583 dcell_lv_0.seg_selector_logic_0.x3/x3.A lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.63463f
C584 decoder_3_0/decoder_2to4_2.b[1] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.07455f
C585 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.04792f
C586 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.14368f
C587 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN dcell_lv_0.bb[9] 0.09979f
C588 decoder_3_0/decoder_2to4_2.b[0] dcell_lv_0.bb[9] 0.33687f
C589 dcell_lv_0.logic_shift_seg2_0.x4.B lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.17656f
C590 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN decoder_3_0/decoder_2to4_1.b[1] 3.75653f
C591 VBNLV decoder_3_0/decoder_2to4_2.bb[1] 0.47152f
C592 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y VDD 0.21864f
C593 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.0897f
C594 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB dcell_lv_0.b[8] 0.12894f
C595 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.06017f
C596 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD 0.21631f
C597 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB decoder_3_0/decoder_2to4_1.b[1] 0.0852f
C598 VBNLV lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 0.01579f
C599 dec1[3] dec0[3] 0.07441f
C600 dcell_lv_0.seg_selector_logic_0.x2/x4.C lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.20013f
C601 VBNLV VDDH 0.18205f
C602 VBPLV seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.30237f
C603 dec1[2] VDDH 0.85004f
C604 dcell_lv_0.bb[8] dcell_lv_0.bb[9] 3.28115f
C605 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_1.b[1] 0.07012f
C606 SH[2] VDDH 0.33127f
C607 dcell_lv_0.seg_selector_logic_0.x2/x4.A VDD 0.35618f
C608 dec1[3] dec0[1] 0.05747f
C609 DIN9 VDD 0.1675f
C610 dcell_lv_0.logic_shift_seg2_0.x7.Y dcell_lv_0.b[9] 0.0152f
C611 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN dcell_lv_0.b[8] 0.14448f
C612 dec1[2] dec2[3] 0.05726f
C613 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.08134f
C614 dec1[0] dec0[1] 0.05039f
C615 decoder_3_0/decoder_2to4_2.bb[1] seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C616 VBNDEC dec0[0] 0.06769f
C617 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.15073f
C618 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB 0.31321f
C619 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 0.08827f
C620 b[0] bb[0] 0.38613f
C621 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09099f
C622 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 8.31336f
C623 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_1.bb[1] 0.13195f
C624 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.09354f
C625 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[1] 0.11776f
C626 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN dcell_lv_0.bb[9] 0.26076f
C627 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.19477f
C628 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A VDDH 0.90535f
C629 DIN8 DIN7 0.0205f
C630 dec2[1] VBPDEC 0.26925f
C631 decoder_3_0/decoder_2to4_2.bb[0] lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.02298f
C632 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN DIN2 0.03543f
C633 dec1[1] VBPDEC 0.26885f
C634 VBNDEC VBPDEC 0.03783f
C635 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04695f
C636 dec2[0] dec2b[1] 0.14127f
C637 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.09312f
C638 dcell_lv_0.seg_selector_logic_0.x1/x3.A seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.01021f
C639 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN dcell_lv_0.b[9] 0.09778f
C640 dcell_lv_0.seg_selector_logic_0.x2/x4.A lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.03886f
C641 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB dcell_lv_0.bb[9] 0.0765f
C642 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.0938f
C643 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[1] 0.42728f
C644 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB dcell_lv_0.bb[9] 0.09135f
C645 dcell_lv_0.seg_selector_logic_0.x3/x3.A lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.1268f
C646 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y decoder_3_0/decoder_2to4_2.bb[0] 0.0203f
C647 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB dcell_lv_0.b[8] 0.13028f
C648 dec0[3] dec0[0] 0.37541f
C649 dec1[3] dec1[2] 0.9809f
C650 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.05433f
C651 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 0.09195f
C652 dcell_lv_0.b[8] VDD 1.73108f
C653 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_2.bb[1] 0.36098f
C654 dcell_lv_0.seg_selector_logic_0.x2/x4.B dcell_lv_0.bb[8] 0.02488f
C655 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN decoder_3_0/decoder_2to4_2.bb[1] 0.47364f
C656 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.09474f
C657 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD 0.2275f
C658 dcell_lv_0.seg_selector_logic_0.x4/x3.B dcell_lv_0.b[8] 0.0151f
C659 dec1[1] dec0[2] 0.05012f
C660 dec1[0] dec1[2] 0.63006f
C661 dec0[1] dec0[0] 1.25358f
C662 VBNDEC dec0[2] 0.07829f
C663 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB decoder_3_0/decoder_2to4_2.bb[0] 0.02583f
C664 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[0] 0.05356f
C665 VBPLV seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.30237f
C666 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB DIN2 0.17961f
C667 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.0935f
C668 VDDH dec2b[3] 0.28782f
C669 dcell_lv_0.seg_selector_logic_0.x3/x3.A seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN 0.21439f
C670 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN decoder_3_0/decoder_2to4_1.b[1] 0.09148f
C671 DIN3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.01594f
C672 DIN3 VDD 0.1713f
C673 dec0[3] VBPDEC 0.1594f
C674 bb[2] b[2] 0.38613f
C675 dcell_lv_0.logic_shift_seg2_0.x4.A decoder_3_0/decoder_2to4_2.b[1] 0.24855f
C676 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB dcell_lv_0.b[9] 0.0923f
C677 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.17257f
C678 dec2b[0] VDDH 0.2239f
C679 decoder_3_0/decoder_2to4_2.b[1] a_7980_n1212# 0.02083f
C680 dec0[1] VBPDEC 0.26885f
C681 decoder_3_0/decoder_2to4_2.bb[1] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB 0.56413f
C682 dec2[3] dec2b[3] 0.43443f
C683 decoder_3_0/decoder_2to4_2.b[0] dcell_lv_0.bb[8] 0.22605f
C684 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN dcell_lv_0.bb[8] 0.0923f
C685 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.05438f
C686 dcell_lv_0.logic_shift_seg2_0.x8.Y decoder_3_0/decoder_2to4_2.b[0] 0.54094f
C687 decoder_3_0/decoder_2to4_1.bb[1] dcell_lv_0.b[8] 10.3939f
C688 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN 0.09276f
C689 DIN5 DIN4 0.0205f
C690 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB dcell_lv_0.b[8] 0.37742f
C691 dcell_lv_0.seg_selector_logic_0.x2/x5.Y VDD 0.49553f
C692 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB dcell_lv_0.bb[9] 0.14375f
C693 VDD dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.25878f
C694 dcell_lv_0.logic_shift_seg2_0.x4.B decoder_3_0/decoder_2to4_2.b[1] 0.21283f
C695 dcell_lv_0.logic_shift_seg2_0.x4.A dcell_lv_0.b[9] 0.13531f
C696 VBNLV VBPLV 0.03932f
C697 dec0[3] dec0[2] 0.9809f
C698 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09485f
C699 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_1.b[1] 0.02113f
C700 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB decoder_3_0/decoder_2to4_1.b[1] 0.08675f
C701 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.06014f
C702 dcell_lv_0.logic_shift_seg2_0.x8.Y dcell_lv_0.bb[8] 0.20641f
C703 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN decoder_3_0/decoder_2to4_2.b[0] 0.041f
C704 dec0[1] dec0[2] 1.23984f
C705 dcell_lv_0.logic_shift_seg2_0.x6.Y decoder_3_0/decoder_2to4_2.b[0] 0.21387f
C706 bb[5] VDDH 0.59451f
C707 dec2[0] VDDH 1.28361f
C708 decoder_3_0/decoder_2to4_2.bb[0] decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.0203f
C709 dcell_lv_0.seg_selector_logic_0.x2/x4.A lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN 0.02611f
C710 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN dcell_lv_0.bb[9] 0.15936f
C711 b[2] VDDH 0.35752f
C712 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.17721f
C713 SH[1] VDDH 0.29652f
C714 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y decoder_3_0/decoder_2to4_2.bb[0] 0.01148f
C715 dcell_lv_0.logic_shift_seg2_0.x4.C decoder_3_0/decoder_2to4_2.b[1] 0.09522f
C716 dcell_lv_0.logic_shift_seg2_0.x4.B dcell_lv_0.logic_shift_seg2_0.x4.A 0.61284f
C717 dcell_lv_0.logic_shift_seg2_0.x4.B dcell_lv_0.b[9] 0.13356f
C718 dcell_lv_0.logic_shift_seg2_0.x4.A decoder_3_0/decoder_2to4_1.b[1] 0.0421f
C719 decoder_3_0/decoder_2to4_1.b[1] dcell_lv_0.b[9] 1.04351f
C720 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB decoder_3_0/decoder_2to4_2.bb[1] 0.22936f
C721 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[0] 0.0761f
C722 VBPLV seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.29848f
C723 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN dcell_lv_0.bb[8] 0.03981f
C724 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN DIN0 0.03542f
C725 dcell_lv_0.seg_selector_logic_0.x2/x5.Y decoder_3_0/decoder_2to4_1.bb[1] 0.22293f
C726 DIN4 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB 0.01591f
C727 dec1[2] VBPDEC 0.19485f
C728 decoder_3_0/decoder_2to4_1.bb[1] dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.02024f
C729 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB 0.09346f
C730 decoder_3_0/decoder_2to4_2.b[0] lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.07676f
C731 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN 9.1182f
C732 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN 0.09039f
C733 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB 0.08478f
C734 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN VDD 6.72553f
C735 dec2[1] dec2[2] 1.32719f
C736 dec2[0] dec2[3] 0.37544f
C737 dcell_lv_0.logic_shift_seg2_0.x6.Y dcell_lv_0.logic_shift_seg2_0.x8.Y 0.10297f
C738 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN dcell_lv_0.bb[9] 0.03731f
C739 dcell_lv_0.seg_selector_logic_0.x2/x4.A decoder_3_0/decoder_2to4_2.bb[0] 0.02308f
C740 dcell_lv_0.seg_selector_logic_0.x2/x5.Y lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.26098f
C741 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.01836f
C742 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y VDD 0.2275f
C743 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN dcell_lv_0.b[8] 0.14066f
C744 VBNDEC dec2[2] 0.07829f
C745 DIN8 dcell_lv_0.b[9] 0.0349f
C746 decoder_3_0/decoder_2to4_2.b[0] seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN 0.04022f
C747 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.38434f
C748 dcell_lv_0.logic_shift_seg2_0.x4.C dcell_lv_0.b[9] 0.05883f
C749 dcell_lv_0.logic_shift_seg2_0.x4.C dcell_lv_0.logic_shift_seg2_0.x4.A 0.01808f
C750 dcell_lv_0.seg_selector_logic_0.x3/x3.B VDD 0.4727f
C751 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.168f
C752 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB dcell_lv_0.bb[8] 0.0543f
C753 dcell_lv_0.logic_shift_seg2_0.x4.B decoder_3_0/decoder_2to4_1.b[1] 0.04684f
C754 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.05001f
C755 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB decoder_3_0/decoder_2to4_2.bb[1] 0.05423f
C756 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y VDD 0.21631f
C757 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB dcell_lv_0.bb[8] 0.08389f
C758 DIN4 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN 0.03501f
C759 decoder_3_0/decoder_2to4_2.b[1] decoder_3_0/decoder_2to4_2.bb[1] 9.03926f
C760 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN dcell_lv_0.b[9] 0.08564f
C761 bb[4] VDDH 0.59451f
C762 decoder_3_0/decoder_2to4_2.bb[1] decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.04783f
C763 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB dcell_lv_0.bb[9] 0.14522f
C764 DIN3 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN 0.03505f
C765 VDD dcell_lv_0.bb[9] 3.68003f
C766 bb[6] VDDH 0.58536f
C767 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB dcell_lv_0.seg_selector_logic_0.x3/x3.A 0.01335f
C768 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB 0.09437f
C769 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN decoder_3_0/decoder_2to4_1.bb[1] 0.11466f
C770 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN dcell_lv_0.b[8] 1.85904f
C771 dcell_lv_0.logic_shift_seg2_0.x4.C dcell_lv_0.logic_shift_seg2_0.x4.B 0.2455f
C772 a_7980_n1756# decoder_3_0/decoder_2to4_2.bb[0] 0.01719f
C773 dec2[1] dec2b[2] 0.13828f
C774 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB 0.4978f
C775 dcell_lv_0.logic_shift_seg2_0.x4.C decoder_3_0/decoder_2to4_1.b[1] 0.26559f
C776 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB 0.25253f
C777 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB dcell_lv_0.b[8] 0.2781f
C778 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB decoder_3_0/decoder_2to4_2.b[0] 0.13975f
C779 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN 0.38843f
C780 dcell_lv_0.seg_selector_logic_0.x3/x3.B decoder_3_0/decoder_2to4_1.bb[1] 0.3076f
C781 DIN0 GND 0.48489f
C782 DIN1 GND 0.46476f
C783 DIN2 GND 0.46241f
C784 DIN3 GND 0.46476f
C785 DIN4 GND 0.46476f
C786 DIN5 GND 0.46465f
C787 DIN6 GND 0.46476f
C788 DIN7 GND 0.46476f
C789 DIN8 GND 0.46476f
C790 DIN9 GND 0.52961f
C791 VBNLV GND 12.5986f
C792 VBNDEC GND 4.28087f
C793 VBPLV GND 5.97493f
C794 dec0[3] GND 0.97496f
C795 dec1[3] GND 0.69193f
C796 dec0[2] GND 0.60586f
C797 dec1[2] GND 0.55796f
C798 dec0[0] GND 0.66499f
C799 dec0[1] GND 0.63592f
C800 dec1[0] GND 0.61627f
C801 dec1[1] GND 0.5825f
C802 b[6] GND 0.38537f
C803 b[5] GND 0.29772f
C804 b[4] GND 0.29772f
C805 b[3] GND 0.29772f
C806 b[2] GND 0.29772f
C807 b[1] GND 0.29772f
C808 b[0] GND 0.29772f
C809 SH[4] GND 0.37966f
C810 SH[3] GND 0.38628f
C811 SH[2] GND 0.38628f
C812 SH[1] GND 0.41932f
C813 bb[6] GND 0.70622f
C814 bb[5] GND 0.69825f
C815 bb[4] GND 0.69825f
C816 bb[3] GND 0.69825f
C817 bb[2] GND 0.69825f
C818 bb[1] GND 0.69825f
C819 bb[0] GND 0.69918f
C820 VBPDEC GND 2.11322f
C821 dec2b[3] GND 0.30107f
C822 dec2b[2] GND 0.2952f
C823 dec2b[1] GND 0.29487f
C824 dec2b[0] GND 0.47474f
C825 dec2[3] GND 1.39381f
C826 dec2[2] GND 1.11364f
C827 dec2[1] GND 1.1383f
C828 dec2[0] GND 1.3096f
C829 VDD GND 45.74228f
C830 VDDH GND 66.16795f
C831 a_7980_n1756# GND 0.02142f $ **FLOATING
C832 decoder_3_0/decoder_2to4_2.bb[0] GND 7.03885f
C833 decoder_3_0/decoder_2to4_2.b[0] GND 8.72121f
C834 dcell_lv_0.logic_shift_seg2_0.x8.Y GND 0.33897f
C835 dcell_lv_0.logic_shift_seg2_0.x6.Y GND 0.70838f
C836 dcell_lv_0.logic_shift_seg2_0.x7.Y GND 0.3768f
C837 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN GND 5.74515f
C838 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB GND 5.93355f
C839 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN GND 6.43251f
C840 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB GND 6.75175f
C841 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN GND 14.46599f
C842 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB GND 12.28317f
C843 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN GND 13.7811f
C844 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB GND 11.73549f
C845 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN GND 13.42611f
C846 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB GND 11.54015f
C847 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN GND 12.12019f
C848 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB GND 11.21747f
C849 a_7980_n884# GND 0.02172f $ **FLOATING
C850 decoder_3_0/decoder_2to4_2.bb[1] GND 7.28464f
C851 decoder_3_0/decoder_2to4_2.b[1] GND 7.20068f
C852 dcell_lv_0.logic_shift_seg2_0.x4.A GND 0.3291f
C853 dcell_lv_0.logic_shift_seg2_0.x4.B GND 0.31137f
C854 dcell_lv_0.logic_shift_seg2_0.x4.C GND 0.33203f
C855 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.75381f
C856 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.63305f
C857 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.66383f
C858 decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.61845f
C859 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.61568f
C860 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.64256f
C861 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.67288f
C862 decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.65617f
C863 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.61395f
C864 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.643f
C865 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.67704f
C866 decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.79418f
C867 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN GND 1.66631f
C868 seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB GND 2.14419f
C869 dcell_lv_0.seg_selector_logic_0.x2/x4.A GND 0.73454f
C870 dcell_lv_0.seg_selector_logic_0.x2/x4.B GND 0.42992f
C871 dcell_lv_0.seg_selector_logic_0.x2/x4.C GND 0.41678f
C872 dcell_lv_0.seg_selector_logic_0.x2/x5.Y GND 0.45218f
C873 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN GND 1.2336f
C874 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB GND 2.40462f
C875 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN GND 3.91072f
C876 dcell_lv_0.seg_selector_logic_0.x3/x3.A GND 0.25661f
C877 dcell_lv_0.seg_selector_logic_0.x3/x3.B GND 0.32574f
C878 seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB GND 1.4861f
C879 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB GND 4.86469f
C880 dcell_lv_0.seg_selector_logic_0.x1/x3.A GND 0.49953f
C881 dcell_lv_0.seg_selector_logic_0.x1/x3.B GND 0.44411f
C882 dcell_lv_0.bb[9] GND 8.03862f
C883 dcell_lv_0.bb[8] GND 3.7934f
C884 decoder_3_0/decoder_2to4_1.bb[1] GND 10.78501f
C885 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB GND 7.92904f
C886 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN GND 4.44299f
C887 dcell_lv_0.seg_selector_logic_0.x4/x3.A GND 0.68096f
C888 dcell_lv_0.seg_selector_logic_0.x4/x3.B GND 0.39649f
C889 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN GND 10.31874f
C890 decoder_3_0/decoder_2to4_1.b[1] GND 9.25869f
C891 dcell_lv_0.b[8] GND 4.70431f
C892 dcell_lv_0.b[9] GND 4.35781f
C893 seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A GND 0.77236f
C894 seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A GND 0.77369f
C895 seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A GND 0.77369f
C896 seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A GND 0.97473f
C897 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t2 GND 0.02802f
C898 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t3 GND 0.02802f
C899 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 GND 0.06156f
C900 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 GND 0.03979f
C901 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t4 GND 0.25825f
C902 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 GND 5.07183f
C903 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t0 GND 0.04311f
C904 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t1 GND 0.04311f
C905 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 GND 0.09914f
C906 lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 GND 0.20106f
C907 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t3 GND 0.02762f
C908 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t2 GND 0.02762f
C909 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 GND 0.06068f
C910 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 GND 0.03922f
C911 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t4 GND 0.25452f
C912 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 GND 4.59489f
C913 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t1 GND 0.04249f
C914 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t0 GND 0.04249f
C915 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 GND 0.09771f
C916 lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 GND 0.19816f
C917 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t1 GND 0.08716f
C918 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t0 GND 0.13242f
C919 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t2 GND 0.21115f
C920 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 GND 3.23299f
C921 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 GND 0.36852f
C922 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n2 GND 0.01016f
C923 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t3 GND 0.02696f
C924 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t2 GND 0.02696f
C925 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 GND 0.05922f
C926 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 GND 0.03828f
C927 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t5 GND 0.06451f
C928 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t4 GND 0.03801f
C929 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t8 GND 0.06451f
C930 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t7 GND 0.03801f
C931 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 GND 0.10824f
C932 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 GND 0.16058f
C933 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 GND 0.04842f
C934 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t6 GND 0.24843f
C935 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 GND 6.79023f
C936 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 GND 0.02983f
C937 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t1 GND 0.04147f
C938 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t0 GND 0.04147f
C939 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 GND 0.09536f
C940 lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 GND 0.1934f
C941 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t3 GND 0.04265f
C942 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t2 GND 0.04265f
C943 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 GND 0.09807f
C944 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 GND 0.19889f
C945 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t6 GND 0.06634f
C946 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t5 GND 0.03909f
C947 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t8 GND 0.06634f
C948 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t7 GND 0.03909f
C949 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 GND 0.11131f
C950 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 GND 0.16514f
C951 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 GND 0.0498f
C952 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t4 GND 0.25549f
C953 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 GND 6.491f
C954 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 GND 0.03068f
C955 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 GND 0.03936f
C956 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t0 GND 0.02772f
C957 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t1 GND 0.02772f
C958 lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 GND 0.0609f
C959 decoder_3_0/decoder_2to4_2.b[1].t3 GND 0.0523f
C960 decoder_3_0/decoder_2to4_2.b[1].t5 GND 0.02729f
C961 decoder_3_0/decoder_2to4_2.b[1].t6 GND 0.04372f
C962 decoder_3_0/decoder_2to4_2.b[1].n0 GND 0.08693f
C963 decoder_3_0/decoder_2to4_2.b[1].t9 GND 0.02734f
C964 decoder_3_0/decoder_2to4_2.b[1].t4 GND 0.04378f
C965 decoder_3_0/decoder_2to4_2.b[1].n1 GND 0.08334f
C966 decoder_3_0/decoder_2to4_2.b[1].n2 GND 0.0164f
C967 decoder_3_0/decoder_2to4_2.b[1].n3 GND 0.03575f
C968 decoder_3_0/decoder_2to4_2.b[1].n4 GND 5.86971f
C969 decoder_3_0/decoder_2to4_2.b[1].t7 GND 0.02736f
C970 decoder_3_0/decoder_2to4_2.b[1].t8 GND 0.04381f
C971 decoder_3_0/decoder_2to4_2.b[1].n5 GND 0.0821f
C972 decoder_3_0/decoder_2to4_2.b[1].n6 GND 0.02222f
C973 decoder_3_0/decoder_2to4_2.b[1].n7 GND 0.29951f
C974 decoder_3_0/decoder_2to4_2.b[1].n8 GND 0.13901f
C975 decoder_3_0/decoder_2to4_2.b[1].t2 GND 0.12153f
C976 decoder_3_0/decoder_2to4_2.b[1].t0 GND 0.02645f
C977 decoder_3_0/decoder_2to4_2.b[1].t1 GND 0.02645f
C978 decoder_3_0/decoder_2to4_2.b[1].n9 GND 0.05879f
C979 decoder_3_0/decoder_2to4_2.b[1].n10 GND 0.29329f
C980 decoder_3_0/decoder_2to4_1.b[1].t3 GND 0.02821f
C981 decoder_3_0/decoder_2to4_1.b[1].t2 GND 0.02821f
C982 decoder_3_0/decoder_2to4_1.b[1].n0 GND 0.06198f
C983 decoder_3_0/decoder_2to4_1.b[1].n1 GND 0.04006f
C984 decoder_3_0/decoder_2to4_1.b[1].t7 GND 0.04479f
C985 decoder_3_0/decoder_2to4_1.b[1].t14 GND 0.07176f
C986 decoder_3_0/decoder_2to4_1.b[1].n2 GND 0.14268f
C987 decoder_3_0/decoder_2to4_1.b[1].t17 GND 0.04486f
C988 decoder_3_0/decoder_2to4_1.b[1].t5 GND 0.07186f
C989 decoder_3_0/decoder_2to4_1.b[1].n3 GND 0.13678f
C990 decoder_3_0/decoder_2to4_1.b[1].n4 GND 0.02691f
C991 decoder_3_0/decoder_2to4_1.b[1].n5 GND 0.07118f
C992 decoder_3_0/decoder_2to4_1.b[1].t6 GND 0.07176f
C993 decoder_3_0/decoder_2to4_1.b[1].t12 GND 0.04479f
C994 decoder_3_0/decoder_2to4_1.b[1].n6 GND 0.14129f
C995 decoder_3_0/decoder_2to4_1.b[1].n7 GND 0.19929f
C996 decoder_3_0/decoder_2to4_1.b[1].n8 GND 0.66039f
C997 decoder_3_0/decoder_2to4_1.b[1].t15 GND 0.04495f
C998 decoder_3_0/decoder_2to4_1.b[1].t16 GND 0.07196f
C999 decoder_3_0/decoder_2to4_1.b[1].n9 GND 0.13234f
C1000 decoder_3_0/decoder_2to4_1.b[1].n10 GND 0.12631f
C1001 decoder_3_0/decoder_2to4_1.b[1].n11 GND 0.75951f
C1002 decoder_3_0/decoder_2to4_1.b[1].t10 GND 0.07176f
C1003 decoder_3_0/decoder_2to4_1.b[1].t9 GND 0.04479f
C1004 decoder_3_0/decoder_2to4_1.b[1].n12 GND 0.14119f
C1005 decoder_3_0/decoder_2to4_1.b[1].n13 GND 0.16454f
C1006 decoder_3_0/decoder_2to4_1.b[1].n14 GND 0.73818f
C1007 decoder_3_0/decoder_2to4_1.b[1].t11 GND 0.04486f
C1008 decoder_3_0/decoder_2to4_1.b[1].t4 GND 0.07186f
C1009 decoder_3_0/decoder_2to4_1.b[1].n15 GND 0.13678f
C1010 decoder_3_0/decoder_2to4_1.b[1].n16 GND 0.29422f
C1011 decoder_3_0/decoder_2to4_1.b[1].n17 GND 0.83984f
C1012 decoder_3_0/decoder_2to4_1.b[1].t13 GND 0.07176f
C1013 decoder_3_0/decoder_2to4_1.b[1].t8 GND 0.04479f
C1014 decoder_3_0/decoder_2to4_1.b[1].n18 GND 0.14124f
C1015 decoder_3_0/decoder_2to4_1.b[1].n19 GND 0.13864f
C1016 decoder_3_0/decoder_2to4_1.b[1].n20 GND 4.55762f
C1017 decoder_3_0/decoder_2to4_1.b[1].n21 GND 11.9797f
C1018 decoder_3_0/decoder_2to4_1.b[1].n22 GND 0.56248f
C1019 decoder_3_0/decoder_2to4_1.b[1].t1 GND 0.04341f
C1020 decoder_3_0/decoder_2to4_1.b[1].t0 GND 0.04341f
C1021 decoder_3_0/decoder_2to4_1.b[1].n23 GND 0.09981f
C1022 decoder_3_0/decoder_2to4_1.b[1].n24 GND 0.20243f
C1023 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t2 GND 0.0216f
C1024 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 GND 0.06193f
C1025 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t3 GND 0.12939f
C1026 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 GND 2.05067f
C1027 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t4 GND 0.03579f
C1028 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t5 GND 0.02235f
C1029 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 GND 0.06697f
C1030 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 GND 0.01708f
C1031 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 GND 0.30063f
C1032 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t1 GND 0.01404f
C1033 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t0 GND 0.01404f
C1034 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 GND 0.05778f
C1035 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n6 GND 0.09765f
C1036 seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n7 GND 0.04153f
C1037 decoder_3_0/decoder_2to4_2.bb[1].t1 GND 0.07759f
C1038 decoder_3_0/decoder_2to4_2.bb[1].t4 GND 0.02253f
C1039 decoder_3_0/decoder_2to4_2.bb[1].t5 GND 0.03611f
C1040 decoder_3_0/decoder_2to4_2.bb[1].n0 GND 0.07179f
C1041 decoder_3_0/decoder_2to4_2.bb[1].t2 GND 0.02257f
C1042 decoder_3_0/decoder_2to4_2.bb[1].t3 GND 0.03615f
C1043 decoder_3_0/decoder_2to4_2.bb[1].n1 GND 0.06882f
C1044 decoder_3_0/decoder_2to4_2.bb[1].n2 GND 0.02009f
C1045 decoder_3_0/decoder_2to4_2.bb[1].n3 GND 4.71088f
C1046 decoder_3_0/decoder_2to4_2.bb[1].n4 GND 0.0984f
C1047 decoder_3_0/decoder_2to4_2.bb[1].t0 GND 0.05929f
C1048 decoder_3_0/decoder_2to4_2.bb[1].n5 GND 0.01959f
C1049 dcell_lv_0.b[9].t3 GND 0.02605f
C1050 dcell_lv_0.b[9].t2 GND 0.02605f
C1051 dcell_lv_0.b[9].n0 GND 0.05724f
C1052 dcell_lv_0.b[9].n1 GND 0.03699f
C1053 dcell_lv_0.b[9].t16 GND 0.04151f
C1054 dcell_lv_0.b[9].t9 GND 0.06645f
C1055 dcell_lv_0.b[9].n2 GND 0.12322f
C1056 dcell_lv_0.b[9].t14 GND 0.04129f
C1057 dcell_lv_0.b[9].t7 GND 0.06618f
C1058 dcell_lv_0.b[9].n3 GND 0.13445f
C1059 dcell_lv_0.b[9].n4 GND 0.15582f
C1060 dcell_lv_0.b[9].t8 GND 0.06626f
C1061 dcell_lv_0.b[9].t15 GND 0.04136f
C1062 dcell_lv_0.b[9].n5 GND 0.13065f
C1063 dcell_lv_0.b[9].n6 GND 0.08905f
C1064 dcell_lv_0.b[9].n7 GND 0.47105f
C1065 dcell_lv_0.b[9].n8 GND 0.84298f
C1066 dcell_lv_0.b[9].t12 GND 0.06626f
C1067 dcell_lv_0.b[9].t11 GND 0.04136f
C1068 dcell_lv_0.b[9].n9 GND 0.13038f
C1069 dcell_lv_0.b[9].n10 GND 0.08233f
C1070 dcell_lv_0.b[9].n11 GND 0.52215f
C1071 dcell_lv_0.b[9].t6 GND 0.04136f
C1072 dcell_lv_0.b[9].t17 GND 0.06626f
C1073 dcell_lv_0.b[9].n12 GND 0.13038f
C1074 dcell_lv_0.b[9].n13 GND 0.05268f
C1075 dcell_lv_0.b[9].t10 GND 0.04136f
C1076 dcell_lv_0.b[9].t4 GND 0.06626f
C1077 dcell_lv_0.b[9].n14 GND 0.13175f
C1078 dcell_lv_0.b[9].t5 GND 0.04143f
C1079 dcell_lv_0.b[9].t13 GND 0.06635f
C1080 dcell_lv_0.b[9].n15 GND 0.1263f
C1081 dcell_lv_0.b[9].n16 GND 0.0229f
C1082 dcell_lv_0.b[9].n17 GND 0.03311f
C1083 dcell_lv_0.b[9].n18 GND 0.46401f
C1084 dcell_lv_0.b[9].n19 GND 11.2596f
C1085 dcell_lv_0.b[9].n20 GND 7.93634f
C1086 dcell_lv_0.b[9].t1 GND 0.04008f
C1087 dcell_lv_0.b[9].t0 GND 0.04008f
C1088 dcell_lv_0.b[9].n21 GND 0.09217f
C1089 dcell_lv_0.b[9].n22 GND 0.18693f
C1090 dcell_lv_0.bb[9].t1 GND 0.0303f
C1091 dcell_lv_0.bb[9].t3 GND 0.0303f
C1092 dcell_lv_0.bb[9].n0 GND 0.06968f
C1093 dcell_lv_0.bb[9].n1 GND 0.14132f
C1094 dcell_lv_0.bb[9].t10 GND 0.04714f
C1095 dcell_lv_0.bb[9].t9 GND 0.02778f
C1096 dcell_lv_0.bb[9].t7 GND 0.04714f
C1097 dcell_lv_0.bb[9].t6 GND 0.02778f
C1098 dcell_lv_0.bb[9].n2 GND 0.07909f
C1099 dcell_lv_0.bb[9].n3 GND 0.11734f
C1100 dcell_lv_0.bb[9].n4 GND 0.03538f
C1101 dcell_lv_0.bb[9].t8 GND 0.05016f
C1102 dcell_lv_0.bb[9].t13 GND 0.03132f
C1103 dcell_lv_0.bb[9].n5 GND 0.09549f
C1104 dcell_lv_0.bb[9].n6 GND 0.14952f
C1105 dcell_lv_0.bb[9].n7 GND 0.74352f
C1106 dcell_lv_0.bb[9].t5 GND 0.0501f
C1107 dcell_lv_0.bb[9].t4 GND 0.03127f
C1108 dcell_lv_0.bb[9].n8 GND 0.09961f
C1109 dcell_lv_0.bb[9].t12 GND 0.05016f
C1110 dcell_lv_0.bb[9].t11 GND 0.03132f
C1111 dcell_lv_0.bb[9].n9 GND 0.09549f
C1112 dcell_lv_0.bb[9].n10 GND 0.01347f
C1113 dcell_lv_0.bb[9].n11 GND 0.34791f
C1114 dcell_lv_0.bb[9].n12 GND 8.73398f
C1115 dcell_lv_0.bb[9].n13 GND 6.92778f
C1116 dcell_lv_0.bb[9].n14 GND 0.0218f
C1117 dcell_lv_0.bb[9].n15 GND 0.02797f
C1118 dcell_lv_0.bb[9].t0 GND 0.0197f
C1119 dcell_lv_0.bb[9].t2 GND 0.0197f
C1120 dcell_lv_0.bb[9].n16 GND 0.04327f
C1121 decoder_3_0/decoder_2to4_2.b[0].t1 GND 0.04115f
C1122 decoder_3_0/decoder_2to4_2.b[0].t6 GND 0.02091f
C1123 decoder_3_0/decoder_2to4_2.b[0].t7 GND 0.0335f
C1124 decoder_3_0/decoder_2to4_2.b[0].n0 GND 0.06386f
C1125 decoder_3_0/decoder_2to4_2.b[0].n1 GND 0.04019f
C1126 decoder_3_0/decoder_2to4_2.b[0].t8 GND 0.02091f
C1127 decoder_3_0/decoder_2to4_2.b[0].t5 GND 0.0335f
C1128 decoder_3_0/decoder_2to4_2.b[0].n2 GND 0.06388f
C1129 decoder_3_0/decoder_2to4_2.b[0].n3 GND 0.01644f
C1130 decoder_3_0/decoder_2to4_2.b[0].n4 GND 0.35374f
C1131 decoder_3_0/decoder_2to4_2.b[0].n5 GND 4.3969f
C1132 decoder_3_0/decoder_2to4_2.b[0].n6 GND 0.1846f
C1133 decoder_3_0/decoder_2to4_2.b[0].t2 GND 0.07487f
C1134 decoder_3_0/decoder_2to4_2.b[0].t4 GND 0.03352f
C1135 decoder_3_0/decoder_2to4_2.b[0].t9 GND 0.02093f
C1136 decoder_3_0/decoder_2to4_2.b[0].n7 GND 0.06281f
C1137 decoder_3_0/decoder_2to4_2.b[0].n8 GND 0.05263f
C1138 decoder_3_0/decoder_2to4_2.b[0].n9 GND 0.14854f
C1139 decoder_3_0/decoder_2to4_2.b[0].t3 GND 0.02023f
C1140 decoder_3_0/decoder_2to4_2.b[0].t0 GND 0.02023f
C1141 decoder_3_0/decoder_2to4_2.b[0].n10 GND 0.04498f
C1142 decoder_3_0/decoder_2to4_2.b[0].n11 GND 0.1296f
C1143 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t1 GND 0.04581f
C1144 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t2 GND 0.10108f
C1145 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 GND 1.41141f
C1146 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n1 GND 0.05865f
C1147 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t0 GND 0.06238f
C1148 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t1 GND 0.05659f
C1149 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 GND 0.02236f
C1150 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t3 GND 0.02938f
C1151 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t5 GND 0.04704f
C1152 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 GND 0.08812f
C1153 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 GND 0.02461f
C1154 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t4 GND 0.17007f
C1155 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 GND 1.97543f
C1156 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 GND 0.32067f
C1157 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 GND 0.04489f
C1158 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 GND 0.01926f
C1159 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t2 GND 0.02839f
C1160 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t0 GND 0.02839f
C1161 seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n8 GND 0.07479f
C1162 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t3 GND 0.03811f
C1163 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t1 GND 0.03811f
C1164 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 GND 0.08764f
C1165 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 GND 0.17775f
C1166 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t11 GND 0.05929f
C1167 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t10 GND 0.03494f
C1168 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t8 GND 0.05929f
C1169 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t7 GND 0.03494f
C1170 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 GND 0.09948f
C1171 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 GND 0.14758f
C1172 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 GND 0.04451f
C1173 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t12 GND 0.03932f
C1174 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t4 GND 0.06301f
C1175 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 GND 0.12528f
C1176 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t5 GND 0.03939f
C1177 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t6 GND 0.06309f
C1178 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 GND 0.1201f
C1179 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 GND 0.03507f
C1180 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t9 GND 0.22833f
C1181 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 GND 8.91454f
C1182 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 GND 3.73702f
C1183 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 GND 0.02742f
C1184 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 GND 0.03518f
C1185 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t2 GND 0.02477f
C1186 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t0 GND 0.02477f
C1187 lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 GND 0.05443f
C1188 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t2 GND 0.02429f
C1189 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t3 GND 0.02429f
C1190 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 GND 0.05336f
C1191 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 GND 0.03449f
C1192 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t11 GND 0.03862f
C1193 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t18 GND 0.06186f
C1194 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 GND 0.11795f
C1195 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 GND 0.07422f
C1196 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t9 GND 0.03862f
C1197 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t17 GND 0.06186f
C1198 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 GND 0.11797f
C1199 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 GND 0.03036f
C1200 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 GND 0.66261f
C1201 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t15 GND 0.22384f
C1202 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 GND 4.3675f
C1203 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t5 GND 0.06186f
C1204 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t10 GND 0.03862f
C1205 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 GND 0.11775f
C1206 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 GND 0.20519f
C1207 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 GND 0.6122f
C1208 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t6 GND 0.03954f
C1209 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t12 GND 0.06298f
C1210 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 GND 0.09489f
C1211 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 GND 0.89543f
C1212 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t14 GND 0.06186f
C1213 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t13 GND 0.03862f
C1214 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 GND 0.11775f
C1215 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 GND 0.22505f
C1216 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 GND 0.81877f
C1217 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t16 GND 0.03862f
C1218 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t8 GND 0.06186f
C1219 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 GND 0.11817f
C1220 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 GND 0.20828f
C1221 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 GND 0.60056f
C1222 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t7 GND 0.06186f
C1223 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t4 GND 0.03862f
C1224 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 GND 0.11775f
C1225 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 GND 0.19927f
C1226 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 GND 4.37812f
C1227 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 GND 8.088f
C1228 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 GND 0.43693f
C1229 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t0 GND 0.03737f
C1230 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t1 GND 0.03737f
C1231 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 GND 0.08593f
C1232 lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 GND 0.17427f
C1233 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t3 GND 0.04058f
C1234 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t1 GND 0.04058f
C1235 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 GND 0.0933f
C1236 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 GND 0.18923f
C1237 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t8 GND 0.06312f
C1238 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t7 GND 0.03719f
C1239 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t6 GND 0.06312f
C1240 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t5 GND 0.03719f
C1241 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 GND 0.1059f
C1242 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 GND 0.15711f
C1243 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 GND 0.04738f
C1244 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t4 GND 0.24308f
C1245 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 GND 6.54065f
C1246 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 GND 0.02919f
C1247 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 GND 0.03745f
C1248 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t2 GND 0.02637f
C1249 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t0 GND 0.02637f
C1250 lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 GND 0.05794f
C1251 decoder_3_0/decoder_2to4_1.bb[1].t1 GND 0.04693f
C1252 decoder_3_0/decoder_2to4_1.bb[1].t3 GND 0.04693f
C1253 decoder_3_0/decoder_2to4_1.bb[1].n0 GND 0.10791f
C1254 decoder_3_0/decoder_2to4_1.bb[1].n1 GND 0.21886f
C1255 decoder_3_0/decoder_2to4_1.bb[1].t9 GND 0.073f
C1256 decoder_3_0/decoder_2to4_1.bb[1].t8 GND 0.04302f
C1257 decoder_3_0/decoder_2to4_1.bb[1].t7 GND 0.073f
C1258 decoder_3_0/decoder_2to4_1.bb[1].t6 GND 0.04302f
C1259 decoder_3_0/decoder_2to4_1.bb[1].n2 GND 0.12249f
C1260 decoder_3_0/decoder_2to4_1.bb[1].n3 GND 0.18172f
C1261 decoder_3_0/decoder_2to4_1.bb[1].n4 GND 0.0548f
C1262 decoder_3_0/decoder_2to4_1.bb[1].t16 GND 0.04842f
C1263 decoder_3_0/decoder_2to4_1.bb[1].t19 GND 0.07759f
C1264 decoder_3_0/decoder_2to4_1.bb[1].n5 GND 0.15426f
C1265 decoder_3_0/decoder_2to4_1.bb[1].t14 GND 0.04851f
C1266 decoder_3_0/decoder_2to4_1.bb[1].t18 GND 0.07769f
C1267 decoder_3_0/decoder_2to4_1.bb[1].n6 GND 0.14788f
C1268 decoder_3_0/decoder_2to4_1.bb[1].n7 GND 0.04318f
C1269 decoder_3_0/decoder_2to4_1.bb[1].t17 GND 0.07769f
C1270 decoder_3_0/decoder_2to4_1.bb[1].t5 GND 0.04851f
C1271 decoder_3_0/decoder_2to4_1.bb[1].n8 GND 0.14788f
C1272 decoder_3_0/decoder_2to4_1.bb[1].n9 GND 0.24277f
C1273 decoder_3_0/decoder_2to4_1.bb[1].n10 GND 0.71242f
C1274 decoder_3_0/decoder_2to4_1.bb[1].t4 GND 0.04834f
C1275 decoder_3_0/decoder_2to4_1.bb[1].t11 GND 0.07749f
C1276 decoder_3_0/decoder_2to4_1.bb[1].n11 GND 0.15742f
C1277 decoder_3_0/decoder_2to4_1.bb[1].n12 GND 0.27042f
C1278 decoder_3_0/decoder_2to4_1.bb[1].n13 GND 1.14249f
C1279 decoder_3_0/decoder_2to4_1.bb[1].t13 GND 0.07909f
C1280 decoder_3_0/decoder_2to4_1.bb[1].t12 GND 0.04966f
C1281 decoder_3_0/decoder_2to4_1.bb[1].n14 GND 0.10732f
C1282 decoder_3_0/decoder_2to4_1.bb[1].n15 GND 1.03162f
C1283 decoder_3_0/decoder_2to4_1.bb[1].t15 GND 0.07909f
C1284 decoder_3_0/decoder_2to4_1.bb[1].t10 GND 0.04966f
C1285 decoder_3_0/decoder_2to4_1.bb[1].n16 GND 0.10732f
C1286 decoder_3_0/decoder_2to4_1.bb[1].n17 GND 5.48586f
C1287 decoder_3_0/decoder_2to4_1.bb[1].n18 GND 11.8351f
C1288 decoder_3_0/decoder_2to4_1.bb[1].n19 GND 1.20346f
C1289 decoder_3_0/decoder_2to4_1.bb[1].n20 GND 0.03376f
C1290 decoder_3_0/decoder_2to4_1.bb[1].n21 GND 0.04331f
C1291 decoder_3_0/decoder_2to4_1.bb[1].t0 GND 0.0305f
C1292 decoder_3_0/decoder_2to4_1.bb[1].t2 GND 0.0305f
C1293 decoder_3_0/decoder_2to4_1.bb[1].n22 GND 0.06701f
C1294 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t3 GND 0.0257f
C1295 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t1 GND 0.0257f
C1296 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 GND 0.05646f
C1297 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 GND 0.03649f
C1298 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t8 GND 0.04079f
C1299 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t4 GND 0.06536f
C1300 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 GND 0.12995f
C1301 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t6 GND 0.04086f
C1302 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t7 GND 0.06545f
C1303 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 GND 0.12458f
C1304 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 GND 0.02451f
C1305 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 GND 0.06483f
C1306 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t5 GND 0.23682f
C1307 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 GND 10.4403f
C1308 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 GND 2.61648f
C1309 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t0 GND 0.03954f
C1310 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t2 GND 0.03954f
C1311 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 GND 0.09091f
C1312 lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 GND 0.18438f
C1313 dcell_lv_0.b[8].t2 GND 0.02814f
C1314 dcell_lv_0.b[8].t3 GND 0.02814f
C1315 dcell_lv_0.b[8].n0 GND 0.06181f
C1316 dcell_lv_0.b[8].n1 GND 0.03995f
C1317 dcell_lv_0.b[8].t5 GND 0.07165f
C1318 dcell_lv_0.b[8].t9 GND 0.04474f
C1319 dcell_lv_0.b[8].n2 GND 0.1364f
C1320 dcell_lv_0.b[8].n3 GND 0.1423f
C1321 dcell_lv_0.b[8].n4 GND 0.50819f
C1322 dcell_lv_0.b[8].t10 GND 0.04581f
C1323 dcell_lv_0.b[8].t14 GND 0.07295f
C1324 dcell_lv_0.b[8].n5 GND 0.09982f
C1325 dcell_lv_0.b[8].n6 GND 0.12298f
C1326 dcell_lv_0.b[8].t13 GND 0.04581f
C1327 dcell_lv_0.b[8].t7 GND 0.07295f
C1328 dcell_lv_0.b[8].n7 GND 0.10991f
C1329 dcell_lv_0.b[8].n8 GND 0.51631f
C1330 dcell_lv_0.b[8].n9 GND 0.64061f
C1331 dcell_lv_0.b[8].t17 GND 0.07168f
C1332 dcell_lv_0.b[8].t16 GND 0.04476f
C1333 dcell_lv_0.b[8].n10 GND 0.13526f
C1334 dcell_lv_0.b[8].n11 GND 0.37535f
C1335 dcell_lv_0.b[8].n12 GND 1.17047f
C1336 dcell_lv_0.b[8].t8 GND 0.04466f
C1337 dcell_lv_0.b[8].t12 GND 0.07156f
C1338 dcell_lv_0.b[8].n13 GND 0.14109f
C1339 dcell_lv_0.b[8].n14 GND 0.12405f
C1340 dcell_lv_0.b[8].n15 GND 0.53513f
C1341 dcell_lv_0.b[8].t4 GND 0.07156f
C1342 dcell_lv_0.b[8].t15 GND 0.04466f
C1343 dcell_lv_0.b[8].n16 GND 0.14228f
C1344 dcell_lv_0.b[8].t11 GND 0.07165f
C1345 dcell_lv_0.b[8].t6 GND 0.04474f
C1346 dcell_lv_0.b[8].n17 GND 0.1364f
C1347 dcell_lv_0.b[8].n18 GND 0.01603f
C1348 dcell_lv_0.b[8].n19 GND 0.16255f
C1349 dcell_lv_0.b[8].n20 GND 12.0678f
C1350 dcell_lv_0.b[8].n21 GND 8.45354f
C1351 dcell_lv_0.b[8].t0 GND 0.04329f
C1352 dcell_lv_0.b[8].t1 GND 0.04329f
C1353 dcell_lv_0.b[8].n22 GND 0.09953f
C1354 dcell_lv_0.b[8].n23 GND 0.20187f
C1355 dcell_lv_0.bb[8].t1 GND 0.04539f
C1356 dcell_lv_0.bb[8].t3 GND 0.04539f
C1357 dcell_lv_0.bb[8].n0 GND 0.10436f
C1358 dcell_lv_0.bb[8].n1 GND 0.21166f
C1359 dcell_lv_0.bb[8].t5 GND 0.0706f
C1360 dcell_lv_0.bb[8].t4 GND 0.0416f
C1361 dcell_lv_0.bb[8].t9 GND 0.0706f
C1362 dcell_lv_0.bb[8].t8 GND 0.0416f
C1363 dcell_lv_0.bb[8].n2 GND 0.11846f
C1364 dcell_lv_0.bb[8].n3 GND 0.17574f
C1365 dcell_lv_0.bb[8].n4 GND 0.053f
C1366 dcell_lv_0.bb[8].t11 GND 0.07503f
C1367 dcell_lv_0.bb[8].t6 GND 0.04683f
C1368 dcell_lv_0.bb[8].n5 GND 0.14763f
C1369 dcell_lv_0.bb[8].n6 GND 0.23929f
C1370 dcell_lv_0.bb[8].n7 GND 1.10227f
C1371 dcell_lv_0.bb[8].t13 GND 0.07513f
C1372 dcell_lv_0.bb[8].t12 GND 0.04691f
C1373 dcell_lv_0.bb[8].n8 GND 0.14301f
C1374 dcell_lv_0.bb[8].n9 GND 0.58286f
C1375 dcell_lv_0.bb[8].n10 GND 1.67264f
C1376 dcell_lv_0.bb[8].t10 GND 0.07516f
C1377 dcell_lv_0.bb[8].t7 GND 0.04693f
C1378 dcell_lv_0.bb[8].n11 GND 0.14182f
C1379 dcell_lv_0.bb[8].n12 GND 0.20135f
C1380 dcell_lv_0.bb[8].n13 GND 11.9265f
C1381 dcell_lv_0.bb[8].n14 GND 9.97149f
C1382 dcell_lv_0.bb[8].n15 GND 0.03265f
C1383 dcell_lv_0.bb[8].n16 GND 0.04189f
C1384 dcell_lv_0.bb[8].t0 GND 0.0295f
C1385 dcell_lv_0.bb[8].t2 GND 0.0295f
C1386 dcell_lv_0.bb[8].n17 GND 0.06481f
C1387 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t1 GND 0.02867f
C1388 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t3 GND 0.02867f
C1389 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 GND 0.06298f
C1390 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 GND 0.04071f
C1391 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t4 GND 0.2642f
C1392 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 GND 4.5886f
C1393 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t2 GND 0.04411f
C1394 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t0 GND 0.04411f
C1395 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 GND 0.10142f
C1396 lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 GND 0.2057f
C1397 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t2 GND 0.02722f
C1398 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t1 GND 0.02722f
C1399 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 GND 0.05979f
C1400 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 GND 0.03864f
C1401 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t13 GND 0.06513f
C1402 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t12 GND 0.03838f
C1403 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t15 GND 0.06513f
C1404 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t14 GND 0.03838f
C1405 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 GND 0.10928f
C1406 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 GND 0.16212f
C1407 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 GND 0.04889f
C1408 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t20 GND 0.0432f
C1409 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t9 GND 0.06922f
C1410 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 GND 0.13633f
C1411 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 GND 0.06254f
C1412 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t10 GND 0.0432f
C1413 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t16 GND 0.06922f
C1414 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 GND 0.13628f
C1415 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 GND 0.04622f
C1416 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 GND 0.71921f
C1417 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t4 GND 0.25083f
C1418 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 GND 4.87592f
C1419 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t19 GND 0.06922f
C1420 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t5 GND 0.0432f
C1421 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 GND 0.1362f
C1422 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 GND 0.12925f
C1423 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 GND 0.86687f
C1424 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t18 GND 0.04431f
C1425 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t6 GND 0.07056f
C1426 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 GND 0.09554f
C1427 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 GND 0.41761f
C1428 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 GND 1.1481f
C1429 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t8 GND 0.06955f
C1430 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t7 GND 0.04347f
C1431 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 GND 0.12226f
C1432 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 GND 0.19214f
C1433 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 GND 0.71521f
C1434 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t17 GND 0.06955f
C1435 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t11 GND 0.04347f
C1436 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 GND 0.12226f
C1437 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 GND 0.11352f
C1438 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 GND 5.23653f
C1439 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 GND 8.0809f
C1440 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 GND 0.99181f
C1441 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 GND 0.03012f
C1442 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t3 GND 0.04187f
C1443 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t0 GND 0.04187f
C1444 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 GND 0.09628f
C1445 lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 GND 0.19526f
C1446 VDD.n0 GND 0.0104f
C1447 VDD.n1 GND 0.01755f
C1448 VDD.t73 GND 0.01283f
C1449 VDD.t3 GND 0.01283f
C1450 VDD.t1 GND 0.01283f
C1451 VDD.n3 GND 0.01499f
C1452 VDD.n4 GND 0.15307f
C1453 VDD.t167 GND 0.01284f
C1454 VDD.n5 GND 0.01789f
C1455 VDD.t59 GND 0.01284f
C1456 VDD.n6 GND 0.01906f
C1457 VDD.t179 GND 0.01284f
C1458 VDD.t165 GND 0.01284f
C1459 VDD.t220 GND 0.01284f
C1460 VDD.t109 GND 0.01284f
C1461 VDD.n11 GND 0.01906f
C1462 VDD.t197 GND 0.01284f
C1463 VDD.t111 GND 0.01284f
C1464 VDD.t51 GND 0.01284f
C1465 VDD.t108 GND 0.02947f
C1466 VDD.t194 GND 0.03942f
C1467 VDD.t196 GND 0.02947f
C1468 VDD.t200 GND 0.03942f
C1469 VDD.t110 GND 0.02947f
C1470 VDD.t34 GND 0.03942f
C1471 VDD.t50 GND 0.02947f
C1472 VDD.t182 GND 0.06986f
C1473 VDD.n16 GND 0.06751f
C1474 VDD.t183 GND 0.01284f
C1475 VDD.n18 GND 0.01789f
C1476 VDD.n20 GND 0.01053f
C1477 VDD.n22 GND 0.01906f
C1478 VDD.t35 GND 0.01284f
C1479 VDD.n23 GND 0.01789f
C1480 VDD.n25 GND 0.01053f
C1481 VDD.n27 GND 0.01906f
C1482 VDD.t201 GND 0.01284f
C1483 VDD.n28 GND 0.01789f
C1484 VDD.n30 GND 0.01053f
C1485 VDD.n32 GND 0.01906f
C1486 VDD.t195 GND 0.01284f
C1487 VDD.n33 GND 0.01789f
C1488 VDD.n35 GND 0.01053f
C1489 VDD.n40 GND 0.06148f
C1490 VDD.t58 GND 0.02947f
C1491 VDD.t176 GND 0.03942f
C1492 VDD.t178 GND 0.02947f
C1493 VDD.t76 GND 0.03942f
C1494 VDD.t164 GND 0.02947f
C1495 VDD.t44 GND 0.03942f
C1496 VDD.t219 GND 0.02947f
C1497 VDD.t81 GND 0.04287f
C1498 VDD.n41 GND 0.07043f
C1499 VDD.t82 GND 0.01284f
C1500 VDD.n46 GND 0.01789f
C1501 VDD.n48 GND 0.01053f
C1502 VDD.n50 GND 0.01906f
C1503 VDD.t45 GND 0.01284f
C1504 VDD.n51 GND 0.01789f
C1505 VDD.n53 GND 0.01053f
C1506 VDD.n55 GND 0.01906f
C1507 VDD.t77 GND 0.01284f
C1508 VDD.n56 GND 0.01789f
C1509 VDD.n58 GND 0.01053f
C1510 VDD.n60 GND 0.01906f
C1511 VDD.t177 GND 0.01284f
C1512 VDD.n61 GND 0.01789f
C1513 VDD.n63 GND 0.01053f
C1514 VDD.n69 GND 0.0578f
C1515 VDD.t155 GND 0.01284f
C1516 VDD.n70 GND 0.01906f
C1517 VDD.t181 GND 0.01284f
C1518 VDD.t157 GND 0.01284f
C1519 VDD.t57 GND 0.01284f
C1520 VDD.n76 GND 0.01053f
C1521 VDD.n78 GND 0.01906f
C1522 VDD.t88 GND 0.01284f
C1523 VDD.n79 GND 0.01789f
C1524 VDD.n81 GND 0.01053f
C1525 VDD.n83 GND 0.01906f
C1526 VDD.t169 GND 0.01284f
C1527 VDD.n84 GND 0.01789f
C1528 VDD.n86 GND 0.01053f
C1529 VDD.n88 GND 0.01906f
C1530 VDD.t235 GND 0.01284f
C1531 VDD.n89 GND 0.01789f
C1532 VDD.n91 GND 0.01053f
C1533 VDD.n96 GND 0.08199f
C1534 VDD.t154 GND 0.02947f
C1535 VDD.t234 GND 0.03942f
C1536 VDD.t180 GND 0.02947f
C1537 VDD.t168 GND 0.03942f
C1538 VDD.t156 GND 0.02947f
C1539 VDD.t87 GND 0.03942f
C1540 VDD.t56 GND 0.02947f
C1541 VDD.t166 GND 0.04287f
C1542 VDD.n97 GND 0.07043f
C1543 VDD.n102 GND 0.12929f
C1544 VDD.n103 GND 0.84719f
C1545 VDD.n104 GND 0.02153f
C1546 VDD.n105 GND 0.02153f
C1547 VDD.n106 GND 0.02153f
C1548 VDD.n107 GND 0.02153f
C1549 VDD.n108 GND 0.02153f
C1550 VDD.n109 GND 0.02153f
C1551 VDD.n110 GND 0.02153f
C1552 VDD.n111 GND 0.02153f
C1553 VDD.t203 GND 0.01283f
C1554 VDD.n112 GND 0.01499f
C1555 VDD.t113 GND 0.01283f
C1556 VDD.n113 GND 0.01615f
C1557 VDD.n114 GND 0.01316f
C1558 VDD.t21 GND 0.01283f
C1559 VDD.n115 GND 0.0104f
C1560 VDD.t47 GND 0.01283f
C1561 VDD.t222 GND 0.01283f
C1562 VDD.n116 GND 0.01499f
C1563 VDD.n117 GND 0.01755f
C1564 VDD.t151 GND 0.01283f
C1565 VDD.n118 GND 0.01316f
C1566 VDD.t15 GND 0.01283f
C1567 VDD.n119 GND 0.0104f
C1568 VDD.t37 GND 0.01283f
C1569 VDD.t137 GND 0.01283f
C1570 VDD.n120 GND 0.01499f
C1571 VDD.n121 GND 0.01755f
C1572 VDD.t11 GND 0.01283f
C1573 VDD.n122 GND 0.01316f
C1574 VDD.t213 GND 0.01283f
C1575 VDD.n123 GND 0.0104f
C1576 VDD.t69 GND 0.01283f
C1577 VDD.t65 GND 0.01283f
C1578 VDD.n124 GND 0.01499f
C1579 VDD.n125 GND 0.01755f
C1580 VDD.t71 GND 0.01283f
C1581 VDD.n126 GND 0.01316f
C1582 VDD.t237 GND 0.01283f
C1583 VDD.n127 GND 0.0104f
C1584 VDD.t209 GND 0.01283f
C1585 VDD.t175 GND 0.01283f
C1586 VDD.n128 GND 0.01499f
C1587 VDD.n129 GND 0.01755f
C1588 VDD.t187 GND 0.01283f
C1589 VDD.n130 GND 0.01316f
C1590 VDD.t33 GND 0.01283f
C1591 VDD.n131 GND 0.0104f
C1592 VDD.t161 GND 0.01283f
C1593 VDD.t159 GND 0.01283f
C1594 VDD.n132 GND 0.01499f
C1595 VDD.n133 GND 0.01755f
C1596 VDD.t79 GND 0.01283f
C1597 VDD.n134 GND 0.01316f
C1598 VDD.t239 GND 0.01283f
C1599 VDD.n135 GND 0.0104f
C1600 VDD.t25 GND 0.01283f
C1601 VDD.t67 GND 0.01283f
C1602 VDD.n136 GND 0.01499f
C1603 VDD.n137 GND 0.01755f
C1604 VDD.t117 GND 0.01283f
C1605 VDD.n138 GND 0.01316f
C1606 VDD.t147 GND 0.01283f
C1607 VDD.n139 GND 0.0104f
C1608 VDD.t55 GND 0.01283f
C1609 VDD.t130 GND 0.01283f
C1610 VDD.n140 GND 0.01499f
C1611 VDD.n141 GND 0.01755f
C1612 VDD.t27 GND 0.01283f
C1613 VDD.n142 GND 0.01316f
C1614 VDD.t139 GND 0.01283f
C1615 VDD.n143 GND 0.0104f
C1616 VDD.t29 GND 0.01283f
C1617 VDD.t92 GND 0.01283f
C1618 VDD.n144 GND 0.01499f
C1619 VDD.t75 GND 0.01283f
C1620 VDD.n145 GND 0.01615f
C1621 VDD.n146 GND 0.0104f
C1622 VDD.n148 GND 0.01316f
C1623 VDD.n149 GND 0.01755f
C1624 VDD.n151 GND 0.01639f
C1625 VDD.n152 GND 0.01515f
C1626 VDD.n154 GND 0.01615f
C1627 VDD.n155 GND 0.0104f
C1628 VDD.n157 GND 0.01316f
C1629 VDD.n158 GND 0.01755f
C1630 VDD.n160 GND 0.01639f
C1631 VDD.n161 GND 0.01515f
C1632 VDD.n163 GND 0.01615f
C1633 VDD.n164 GND 0.0104f
C1634 VDD.n166 GND 0.01316f
C1635 VDD.n167 GND 0.01755f
C1636 VDD.n169 GND 0.01639f
C1637 VDD.n170 GND 0.01515f
C1638 VDD.n172 GND 0.01615f
C1639 VDD.n173 GND 0.0104f
C1640 VDD.n175 GND 0.01316f
C1641 VDD.n176 GND 0.01755f
C1642 VDD.n178 GND 0.01639f
C1643 VDD.n179 GND 0.01515f
C1644 VDD.n181 GND 0.01615f
C1645 VDD.n182 GND 0.0104f
C1646 VDD.n184 GND 0.01316f
C1647 VDD.n185 GND 0.01755f
C1648 VDD.n187 GND 0.01639f
C1649 VDD.n188 GND 0.01515f
C1650 VDD.n190 GND 0.01615f
C1651 VDD.n191 GND 0.0104f
C1652 VDD.n193 GND 0.01316f
C1653 VDD.n194 GND 0.01755f
C1654 VDD.n196 GND 0.01639f
C1655 VDD.n197 GND 0.01515f
C1656 VDD.n199 GND 0.01615f
C1657 VDD.n200 GND 0.0104f
C1658 VDD.n202 GND 0.01316f
C1659 VDD.n203 GND 0.01755f
C1660 VDD.n205 GND 0.01639f
C1661 VDD.n206 GND 0.01515f
C1662 VDD.n208 GND 0.01615f
C1663 VDD.n209 GND 0.0104f
C1664 VDD.n211 GND 0.01316f
C1665 VDD.n212 GND 0.01755f
C1666 VDD.n214 GND 0.01639f
C1667 VDD.n215 GND 0.01515f
C1668 VDD.n217 GND 0.01755f
C1669 VDD.n218 GND 0.0104f
C1670 VDD.n219 GND 0.0104f
C1671 VDD.n221 GND 0.30168f
C1672 VDD.n224 GND 0.01153f
C1673 VDD.t53 GND 0.01283f
C1674 VDD.n225 GND 0.01316f
C1675 VDD.t60 GND 0.05939f
C1676 VDD.t52 GND 0.03239f
C1677 VDD.t89 GND 0.03577f
C1678 VDD.t223 GND 0.02531f
C1679 VDD.n227 GND 0.02741f
C1680 VDD.t224 GND 0.01281f
C1681 VDD.t43 GND 0.0126f
C1682 VDD.n229 GND 0.01524f
C1683 VDD.t7 GND 0.01284f
C1684 VDD.n230 GND 0.01053f
C1685 VDD.n232 GND 0.03851f
C1686 VDD.t189 GND 0.01284f
C1687 VDD.n233 GND 0.01053f
C1688 VDD.t133 GND 0.01284f
C1689 VDD.t39 GND 0.01284f
C1690 VDD.n234 GND 0.03159f
C1691 VDD.t63 GND 0.01284f
C1692 VDD.t232 GND 0.0577f
C1693 VDD.t198 GND 0.03239f
C1694 VDD.t210 GND 0.03577f
C1695 VDD.t6 GND 0.03071f
C1696 VDD.t123 GND 0.04184f
C1697 VDD.t42 GND 0.03239f
C1698 VDD.t227 GND 0.02834f
C1699 VDD.t188 GND 0.02834f
C1700 VDD.t125 GND 0.02295f
C1701 VDD.n236 GND 0.08384f
C1702 VDD.t40 GND 0.07559f
C1703 VDD.t62 GND 0.05197f
C1704 VDD.t38 GND 0.06951f
C1705 VDD.t190 GND 0.05197f
C1706 VDD.n237 GND 0.11745f
C1707 VDD.t143 GND 0.01284f
C1708 VDD.n238 GND 0.01906f
C1709 VDD.t17 GND 0.01284f
C1710 VDD.n240 GND 0.01906f
C1711 VDD.t128 GND 0.01284f
C1712 VDD.t226 GND 0.01284f
C1713 VDD.t205 GND 0.01284f
C1714 VDD.n243 GND 0.01848f
C1715 VDD.n244 GND 0.01053f
C1716 VDD.t149 GND 0.01285f
C1717 VDD.t16 GND 0.02947f
C1718 VDD.t127 GND 0.03942f
C1719 VDD.t225 GND 0.02947f
C1720 VDD.t204 GND 0.03981f
C1721 VDD.t80 GND 0.02603f
C1722 VDD.t148 GND 0.06505f
C1723 VDD.n246 GND 0.08608f
C1724 VDD.n247 GND 0.06619f
C1725 VDD.n248 GND 0.02197f
C1726 VDD.n253 GND 0.01053f
C1727 VDD.n255 GND 0.01906f
C1728 VDD.n256 GND 0.01789f
C1729 VDD.n258 GND 0.01053f
C1730 VDD.n265 GND 0.01053f
C1731 VDD.t122 GND 0.01284f
C1732 VDD.n267 GND 0.01789f
C1733 VDD.t215 GND 0.01284f
C1734 VDD.n268 GND 0.01906f
C1735 VDD.n270 GND 0.01053f
C1736 VDD.t103 GND 0.01284f
C1737 VDD.n272 GND 0.01848f
C1738 VDD.n275 GND 0.01053f
C1739 VDD.t5 GND 0.01285f
C1740 VDD.n277 GND 0.02256f
C1741 VDD.t145 GND 0.01283f
C1742 VDD.n279 GND 0.01371f
C1743 VDD.n281 GND 0.01053f
C1744 VDD.n284 GND 0.02171f
C1745 VDD.n285 GND 0.05576f
C1746 VDD.t144 GND 0.05607f
C1747 VDD.t4 GND 0.04038f
C1748 VDD.t171 GND 0.02603f
C1749 VDD.t102 GND 0.03981f
C1750 VDD.t214 GND 0.02947f
C1751 VDD.t121 GND 0.03942f
C1752 VDD.t142 GND 0.02947f
C1753 VDD.n286 GND 0.04616f
C1754 VDD.n288 GND 0.11784f
C1755 VDD.t107 GND 0.01282f
C1756 VDD.t132 GND 0.01284f
C1757 VDD.n289 GND 0.03277f
C1758 VDD.t185 GND 0.01282f
C1759 VDD.t9 GND 0.01284f
C1760 VDD.n290 GND 0.03277f
C1761 VDD.t141 GND 0.01402f
C1762 VDD.n291 GND 0.01471f
C1763 VDD.t230 GND 0.01282f
C1764 VDD.t153 GND 0.0126f
C1765 VDD.t49 GND 0.01402f
C1766 VDD.t84 GND 0.01282f
C1767 VDD.n294 GND 0.02811f
C1768 VDD.t184 GND 0.02295f
C1769 VDD.t8 GND 0.02834f
C1770 VDD.t192 GND 0.02834f
C1771 VDD.t152 GND 0.02834f
C1772 VDD.t22 GND 0.04724f
C1773 VDD.n295 GND 0.03821f
C1774 VDD.n296 GND 0.01053f
C1775 VDD.t13 GND 0.01284f
C1776 VDD.t231 GND 0.01284f
C1777 VDD.t217 GND 0.0126f
C1778 VDD.t98 GND 0.01259f
C1779 VDD.n299 GND 0.01309f
C1780 VDD.t48 GND 0.02565f
C1781 VDD.t83 GND 0.03037f
C1782 VDD.t18 GND 0.02362f
C1783 VDD.t12 GND 0.03239f
C1784 VDD.t162 GND 0.06985f
C1785 VDD.t216 GND 0.03543f
C1786 VDD.t97 GND 0.02834f
C1787 VDD.t206 GND 0.04285f
C1788 VDD.t114 GND 0.04859f
C1789 VDD.n302 GND 0.03821f
C1790 VDD.t119 GND 0.01388f
C1791 VDD.t135 GND 0.01283f
C1792 VDD.t170 GND 0.01283f
C1793 VDD.n308 GND 0.0247f
C1794 VDD.n310 GND 0.01053f
C1795 VDD.n312 GND 0.05867f
C1796 VDD.n313 GND 0.13584f
C1797 VDD.t134 GND 0.13218f
C1798 VDD.t118 GND 0.03104f
C1799 VDD.n314 GND 0.0497f
C1800 VDD.n315 GND 0.01964f
C1801 VDD.n316 GND 0.01239f
C1802 VDD.n317 GND 0.02224f
C1803 VDD.n321 GND 0.01053f
C1804 VDD.n324 GND 0.01522f
C1805 VDD.n325 GND 0.01804f
C1806 VDD.n326 GND 0.01181f
C1807 VDD.n327 GND 0.01859f
C1808 VDD.n331 GND 0.02161f
C1809 VDD.n332 GND 0.01522f
C1810 VDD.n336 GND 0.01053f
C1811 VDD.t173 GND 0.01284f
C1812 VDD.t101 GND 0.0126f
C1813 VDD.n342 GND 0.01053f
C1814 VDD.n345 GND 0.01522f
C1815 VDD.n346 GND 0.01896f
C1816 VDD.n350 GND 0.03492f
C1817 VDD.n351 GND 0.04698f
C1818 VDD.t229 GND 0.04454f
C1819 VDD.t172 GND 0.03374f
C1820 VDD.t140 GND 0.02362f
C1821 VDD.t30 GND 0.04117f
C1822 VDD.t100 GND 0.02834f
C1823 VDD.t85 GND 0.02834f
C1824 VDD.t131 GND 0.02834f
C1825 VDD.t106 GND 0.02295f
C1826 VDD.n352 GND 0.08735f
C1827 VDD.n354 GND 0.16127f
C1828 VDD.n355 GND 0.45062f
C1829 VDD.n356 GND 0.0506f
C1830 VDD.n358 GND 0.03851f
C1831 VDD.t191 GND 0.01284f
C1832 VDD.t218 GND 0.01284f
C1833 VDD.n359 GND 0.03384f
C1834 VDD.n361 GND 0.01053f
C1835 VDD.t120 GND 0.01284f
C1836 VDD.n364 GND 0.03384f
C1837 VDD.t41 GND 0.01284f
C1838 VDD.t99 GND 0.01284f
C1839 VDD.n366 GND 0.03159f
C1840 VDD.t126 GND 0.01282f
C1841 VDD.n370 GND 0.0325f
C1842 VDD.n372 GND 0.01016f
C1843 VDD.n376 GND 0.01813f
C1844 VDD.t199 GND 0.01283f
C1845 VDD.n378 GND 0.01316f
C1846 VDD.n380 GND 0.01153f
C1847 VDD.n381 GND 0.01053f
C1848 VDD.n384 GND 0.03575f
C1849 VDD.n387 GND 0.01053f
C1850 VDD.n392 GND 0.01053f
C1851 VDD.n393 GND 0.01007f
C1852 VDD.n395 GND 0.06069f
C1853 VDD.n396 GND 0.13869f
C1854 VDD.n397 GND 0.74816f
C1855 VDD.t105 GND 0.01283f
C1856 VDD.n398 GND 0.01428f
C1857 VDD.n399 GND 0.0104f
C1858 VDD.n400 GND 0.01755f
C1859 VDD.n401 GND 0.01316f
C1860 VDD.t96 GND 0.01283f
C1861 VDD.n402 GND 0.01515f
C1862 VDD.t94 GND 0.01283f
C1863 VDD.n403 GND 0.01639f
C1864 VDD.n405 GND 0.01755f
C1865 VDD.n406 GND 0.01316f
C1866 VDD.n408 GND 0.02153f
C1867 VDD.t104 GND 0.0289f
C1868 VDD.t95 GND 0.04f
C1869 VDD.t93 GND 0.0289f
C1870 VDD.t202 GND 0.04325f
C1871 VDD.n409 GND 0.04734f
C1872 VDD.t112 GND 0.0289f
C1873 VDD.t20 GND 0.04f
C1874 VDD.t46 GND 0.0289f
C1875 VDD.t221 GND 0.04325f
C1876 VDD.n410 GND 0.04734f
C1877 VDD.t150 GND 0.0289f
C1878 VDD.t14 GND 0.04f
C1879 VDD.t36 GND 0.0289f
C1880 VDD.t136 GND 0.04325f
C1881 VDD.n411 GND 0.04734f
C1882 VDD.t10 GND 0.0289f
C1883 VDD.t212 GND 0.04f
C1884 VDD.t68 GND 0.0289f
C1885 VDD.t64 GND 0.04325f
C1886 VDD.n412 GND 0.04734f
C1887 VDD.t70 GND 0.0289f
C1888 VDD.t236 GND 0.04f
C1889 VDD.t208 GND 0.0289f
C1890 VDD.t174 GND 0.04325f
C1891 VDD.n413 GND 0.04734f
C1892 VDD.t186 GND 0.0289f
C1893 VDD.t32 GND 0.04f
C1894 VDD.t160 GND 0.0289f
C1895 VDD.t158 GND 0.04325f
C1896 VDD.n414 GND 0.04734f
C1897 VDD.t78 GND 0.0289f
C1898 VDD.t238 GND 0.04f
C1899 VDD.t24 GND 0.0289f
C1900 VDD.t66 GND 0.04325f
C1901 VDD.n415 GND 0.04734f
C1902 VDD.t116 GND 0.0289f
C1903 VDD.t146 GND 0.04f
C1904 VDD.t54 GND 0.0289f
C1905 VDD.t129 GND 0.04325f
C1906 VDD.n416 GND 0.04734f
C1907 VDD.t26 GND 0.0289f
C1908 VDD.t138 GND 0.04f
C1909 VDD.t28 GND 0.0289f
C1910 VDD.t91 GND 0.04325f
C1911 VDD.n417 GND 0.04734f
C1912 VDD.t74 GND 0.0289f
C1913 VDD.t72 GND 0.04f
C1914 VDD.t2 GND 0.0289f
C1915 VDD.t0 GND 0.06517f
C1916 VDD.n418 GND 0.06321f
C1917 VDD.n419 GND 0.34083f
C1918 VDD.n420 GND 0.01316f
C1919 VDD.n421 GND 0.01755f
C1920 VDD.n423 GND 0.01639f
C1921 VDD.n424 GND 0.01515f
C1922 VDD.n425 GND 0.01316f
C1923 VBPDEC.t5 GND 0.17088f
C1924 VBPDEC.n0 GND 0.11518f
C1925 VBPDEC.t7 GND 0.17088f
C1926 VBPDEC.n1 GND 0.12568f
C1927 VBPDEC.t4 GND 0.17088f
C1928 VBPDEC.n2 GND 0.12568f
C1929 VBPDEC.t10 GND 0.17088f
C1930 VBPDEC.n3 GND 0.09212f
C1931 VBPDEC.t11 GND 0.17088f
C1932 VBPDEC.n4 GND 0.09212f
C1933 VBPDEC.t2 GND 0.17088f
C1934 VBPDEC.n5 GND 0.12568f
C1935 VBPDEC.t8 GND 0.17088f
C1936 VBPDEC.n6 GND 0.12568f
C1937 VBPDEC.t3 GND 0.17088f
C1938 VBPDEC.n7 GND 0.12434f
C1939 VBPDEC.t0 GND 0.17088f
C1940 VBPDEC.n8 GND 0.09212f
C1941 VBPDEC.t9 GND 0.17088f
C1942 VBPDEC.n9 GND 0.12568f
C1943 VBPDEC.t6 GND 0.17088f
C1944 VBPDEC.n10 GND 0.12568f
C1945 VBPDEC.t1 GND 0.17088f
C1946 VBPDEC.n11 GND 0.12434f
C1947 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t2 GND 0.038f
C1948 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t3 GND 0.038f
C1949 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 GND 0.08737f
C1950 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 GND 0.1772f
C1951 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t4 GND 0.2276f
C1952 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 GND 4.74263f
C1953 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 GND 0.03507f
C1954 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t0 GND 0.0247f
C1955 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t1 GND 0.0247f
C1956 lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 GND 0.05426f
C1957 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t2 GND 0.04021f
C1958 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t3 GND 0.04021f
C1959 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 GND 0.09246f
C1960 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 GND 0.18752f
C1961 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t5 GND 0.06255f
C1962 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t4 GND 0.03686f
C1963 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t8 GND 0.06255f
C1964 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t7 GND 0.03686f
C1965 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 GND 0.10495f
C1966 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 GND 0.1557f
C1967 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 GND 0.04695f
C1968 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t6 GND 0.24088f
C1969 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 GND 6.85844f
C1970 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 GND 0.02892f
C1971 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 GND 0.03711f
C1972 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t1 GND 0.02614f
C1973 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t0 GND 0.02614f
C1974 lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 GND 0.05742f
C1975 VDDH.n0 GND 0.02048f
C1976 VDDH.n3 GND 0.11759f
C1977 VDDH.n4 GND 0.02048f
C1978 VDDH.n7 GND 0.10372f
C1979 VDDH.n8 GND 0.05756f
C1980 VDDH.n9 GND 0.04638f
C1981 VDDH.n10 GND 0.02628f
C1982 VDDH.n11 GND 0.02048f
C1983 VDDH.t8 GND 0.04775f
C1984 VDDH.n17 GND 0.05094f
C1985 VDDH.t28 GND 0.31875f
C1986 VDDH.t27 GND 0.21407f
C1987 VDDH.t47 GND 0.01232f
C1988 VDDH.n18 GND 0.05083f
C1989 VDDH.n21 GND 0.18813f
C1990 VDDH.t11 GND 0.2419f
C1991 VDDH.t1 GND 0.18968f
C1992 VDDH.n22 GND 0.15349f
C1993 VDDH.t35 GND 0.21407f
C1994 VDDH.t2 GND 0.2912f
C1995 VDDH.t3 GND 0.2912f
C1996 VDDH.t39 GND 0.18968f
C1997 VDDH.n23 GND 0.20533f
C1998 VDDH.n24 GND 0.04638f
C1999 VDDH.n25 GND 0.02628f
C2000 VDDH.n27 GND 0.02602f
C2001 VDDH.n28 GND 0.02905f
C2002 VDDH.n29 GND 0.02717f
C2003 VDDH.n30 GND 0.02824f
C2004 VDDH.n32 GND 0.02602f
C2005 VDDH.n33 GND 0.02905f
C2006 VDDH.n35 GND 0.02273f
C2007 VDDH.n38 GND 0.02048f
C2008 VDDH.n43 GND 0.02273f
C2009 VDDH.n48 GND 0.11759f
C2010 VDDH.n49 GND 0.12991f
C2011 VDDH.t17 GND 0.04775f
C2012 VDDH.n50 GND 0.05083f
C2013 VDDH.n59 GND 0.02273f
C2014 VDDH.n62 GND 0.02628f
C2015 VDDH.n63 GND 0.04638f
C2016 VDDH.n64 GND 0.14777f
C2017 VDDH.n65 GND 0.06316f
C2018 VDDH.t9 GND 0.04775f
C2019 VDDH.n66 GND 0.05083f
C2020 VDDH.n73 GND 0.02273f
C2021 VDDH.n78 GND 0.12632f
C2022 VDDH.n79 GND 0.05083f
C2023 VDDH.t22 GND 0.1108f
C2024 VDDH.n80 GND 0.01529f
C2025 VDDH.n83 GND 0.19122f
C2026 VDDH.t62 GND 0.07959f
C2027 VDDH.n87 GND 0.02577f
C2028 VDDH.n93 GND 0.0333f
C2029 VDDH.n94 GND 0.02926f
C2030 VDDH.t102 GND 0.02496f
C2031 VDDH.t18 GND 0.09933f
C2032 VDDH.t84 GND 0.02577f
C2033 VDDH.t132 GND 0.02577f
C2034 VDDH.n100 GND 0.04858f
C2035 VDDH.n103 GND 0.05704f
C2036 VDDH.n104 GND 0.02273f
C2037 VDDH.n109 GND 0.02657f
C2038 VDDH.t0 GND 0.07982f
C2039 VDDH.n110 GND 0.04885f
C2040 VDDH.n115 GND 0.02273f
C2041 VDDH.n118 GND 0.01f
C2042 VDDH.n121 GND 0.02926f
C2043 VDDH.n122 GND 0.02577f
C2044 VDDH.n123 GND 0.03313f
C2045 VDDH.n124 GND 0.03313f
C2046 VDDH.n126 GND 0.0333f
C2047 VDDH.n127 GND 0.02926f
C2048 VDDH.t116 GND 0.02496f
C2049 VDDH.n132 GND 0.02926f
C2050 VDDH.t106 GND 0.02496f
C2051 VDDH.n133 GND 0.02657f
C2052 VDDH.n136 GND 0.01f
C2053 VDDH.n139 GND 0.02273f
C2054 VDDH.n144 GND 0.04885f
C2055 VDDH.t4 GND 0.07982f
C2056 VDDH.t38 GND 0.07959f
C2057 VDDH.t108 GND 0.02577f
C2058 VDDH.t15 GND 0.02577f
C2059 VDDH.n146 GND 0.04858f
C2060 VDDH.n149 GND 0.02446f
C2061 VDDH.n152 GND 0.02273f
C2062 VDDH.n158 GND 0.02446f
C2063 VDDH.n159 GND 0.19122f
C2064 VDDH.n163 GND 0.02657f
C2065 VDDH.t130 GND 0.02577f
C2066 VDDH.n168 GND 0.02657f
C2067 VDDH.n171 GND 0.04885f
C2068 VDDH.t25 GND 0.07982f
C2069 VDDH.t57 GND 0.07959f
C2070 VDDH.n172 GND 0.04858f
C2071 VDDH.n177 GND 0.0333f
C2072 VDDH.n179 GND 0.02273f
C2073 VDDH.t118 GND 0.02577f
C2074 VDDH.n185 GND 0.02926f
C2075 VDDH.n186 GND 0.02577f
C2076 VDDH.t124 GND 0.02496f
C2077 VDDH.n187 GND 0.02926f
C2078 VDDH.n190 GND 0.01f
C2079 VDDH.n193 GND 0.02273f
C2080 VDDH.n198 GND 0.04885f
C2081 VDDH.t10 GND 0.07982f
C2082 VDDH.t69 GND 0.07959f
C2083 VDDH.n199 GND 0.02577f
C2084 VDDH.n204 GND 0.03313f
C2085 VDDH.n206 GND 0.0333f
C2086 VDDH.n207 GND 0.02926f
C2087 VDDH.t112 GND 0.02496f
C2088 VDDH.n212 GND 0.02926f
C2089 VDDH.t100 GND 0.02496f
C2090 VDDH.n213 GND 0.02657f
C2091 VDDH.n216 GND 0.01f
C2092 VDDH.n219 GND 0.02273f
C2093 VDDH.n224 GND 0.04885f
C2094 VDDH.t70 GND 0.07982f
C2095 VDDH.t76 GND 0.07959f
C2096 VDDH.t92 GND 0.02577f
C2097 VDDH.t55 GND 0.02577f
C2098 VDDH.n226 GND 0.04858f
C2099 VDDH.n229 GND 0.02446f
C2100 VDDH.n232 GND 0.02273f
C2101 VDDH.n238 GND 0.02446f
C2102 VDDH.n239 GND 0.19122f
C2103 VDDH.n241 GND 0.03927f
C2104 VDDH.t128 GND 0.07443f
C2105 VDDH.n244 GND 0.02657f
C2106 VDDH.t65 GND 0.02577f
C2107 VDDH.n249 GND 0.02657f
C2108 VDDH.n252 GND 0.04885f
C2109 VDDH.t83 GND 0.07982f
C2110 VDDH.t49 GND 0.07959f
C2111 VDDH.n253 GND 0.04858f
C2112 VDDH.n258 GND 0.0333f
C2113 VDDH.n260 GND 0.02273f
C2114 VDDH.t98 GND 0.02577f
C2115 VDDH.n266 GND 0.02926f
C2116 VDDH.n267 GND 0.02577f
C2117 VDDH.t122 GND 0.02496f
C2118 VDDH.n268 GND 0.02926f
C2119 VDDH.n271 GND 0.01f
C2120 VDDH.n274 GND 0.02273f
C2121 VDDH.n279 GND 0.04885f
C2122 VDDH.t21 GND 0.08204f
C2123 VDDH.t29 GND 0.07989f
C2124 VDDH.t110 GND 0.04854f
C2125 VDDH.n280 GND 0.03293f
C2126 VDDH.n283 GND 0.03927f
C2127 VDDH.t53 GND 0.07443f
C2128 VDDH.t88 GND 0.04854f
C2129 VDDH.t34 GND 0.08224f
C2130 VDDH.t52 GND 0.08224f
C2131 VDDH.t120 GND 0.04854f
C2132 VDDH.n286 GND 0.03293f
C2133 VDDH.n288 GND 0.03439f
C2134 VDDH.n290 GND 0.03927f
C2135 VDDH.t79 GND 0.07443f
C2136 VDDH.t94 GND 0.04854f
C2137 VDDH.n293 GND 0.03313f
C2138 VDDH.n294 GND 0.03313f
C2139 VDDH.n296 GND 0.03927f
C2140 VDDH.t74 GND 0.07443f
C2141 VDDH.n300 GND 0.02273f
C2142 VDDH.n307 GND 0.02576f
C2143 VDDH.t96 GND 0.04854f
C2144 VDDH.t40 GND 0.08224f
C2145 VDDH.t73 GND 0.08224f
C2146 VDDH.t86 GND 0.04854f
C2147 VDDH.t5 GND 0.08224f
C2148 VDDH.t26 GND 0.08224f
C2149 VDDH.t104 GND 0.04854f
C2150 VDDH.n308 GND 0.03293f
C2151 VDDH.n309 GND 0.03313f
C2152 VDDH.n310 GND 0.03313f
C2153 VDDH.t14 GND 0.10184f
C2154 VDDH.t114 GND 0.04854f
C2155 VDDH.n311 GND 0.03293f
C2156 VDDH.n313 GND 0.02273f
C2157 VDDH.n318 GND 0.02576f
C2158 VDDH.n321 GND 0.03439f
C2159 VDDH.n322 GND 0.18644f
C2160 VDDH.n323 GND 0.02273f
C2161 VDDH.n328 GND 0.02576f
C2162 VDDH.n331 GND 0.03439f
C2163 VDDH.n332 GND 0.02273f
C2164 VDDH.n337 GND 0.02576f
C2165 VDDH.n340 GND 0.03439f
C2166 VDDH.n341 GND 0.19122f
C2167 VDDH.n342 GND 0.19122f
C2168 VDDH.n344 GND 0.02273f
C2169 VDDH.n347 GND 0.01f
C2170 VDDH.n350 GND 0.02926f
C2171 VDDH.n351 GND 0.02577f
C2172 VDDH.n352 GND 0.03313f
C2173 VDDH.n353 GND 0.03313f
C2174 VDDH.n354 GND 0.0333f
C2175 VDDH.n355 GND 0.02273f
C2176 VDDH.n360 GND 0.02926f
C2177 VDDH.t126 GND 0.02577f
C2178 VDDH.t58 GND 0.02577f
C2179 VDDH.n362 GND 0.04858f
C2180 VDDH.n365 GND 0.02446f
C2181 VDDH.n366 GND 0.19122f
C2182 VDDH.n367 GND 0.19122f
C2183 VDDH.n369 GND 0.02273f
C2184 VDDH.n372 GND 0.01f
C2185 VDDH.n375 GND 0.02926f
C2186 VDDH.n376 GND 0.02577f
C2187 VDDH.n377 GND 0.03313f
C2188 VDDH.n378 GND 0.03313f
C2189 VDDH.n379 GND 0.0333f
C2190 VDDH.n380 GND 0.02273f
C2191 VDDH.n385 GND 0.02926f
C2192 VDDH.t90 GND 0.02577f
C2193 VDDH.t32 GND 0.02577f
C2194 VDDH.n387 GND 0.04858f
C2195 VDDH.n390 GND 0.02446f
C2196 VDDH.n391 GND 0.21225f
C2197 VBPLV.t21 GND 0.23663f
C2198 VBPLV.n0 GND 0.19708f
C2199 VBPLV.t12 GND 0.23663f
C2200 VBPLV.n1 GND 0.20844f
C2201 VBPLV.t6 GND 0.23663f
C2202 VBPLV.n2 GND 0.20844f
C2203 VBPLV.t16 GND 0.23663f
C2204 VBPLV.n3 GND 0.20844f
C2205 VBPLV.t11 GND 0.23663f
C2206 VBPLV.n4 GND 0.20844f
C2207 VBPLV.t20 GND 0.23663f
C2208 VBPLV.n5 GND 0.20844f
C2209 VBPLV.t15 GND 0.23663f
C2210 VBPLV.n6 GND 0.20844f
C2211 VBPLV.t3 GND 0.23663f
C2212 VBPLV.n7 GND 0.20844f
C2213 VBPLV.t19 GND 0.23663f
C2214 VBPLV.n8 GND 0.20844f
C2215 VBPLV.t8 GND 0.23663f
C2216 VBPLV.n9 GND 0.20844f
C2217 VBPLV.t2 GND 0.23663f
C2218 VBPLV.n10 GND 0.20844f
C2219 VBPLV.t14 GND 0.23663f
C2220 VBPLV.n11 GND 0.20844f
C2221 VBPLV.t7 GND 0.23663f
C2222 VBPLV.n12 GND 0.20844f
C2223 VBPLV.t17 GND 0.23663f
C2224 VBPLV.n13 GND 0.20844f
C2225 VBPLV.t13 GND 0.23663f
C2226 VBPLV.n14 GND 0.20844f
C2227 VBPLV.t0 GND 0.23663f
C2228 VBPLV.n15 GND 0.20844f
C2229 VBPLV.t1 GND 0.23663f
C2230 VBPLV.n16 GND 0.20844f
C2231 VBPLV.t4 GND 0.23663f
C2232 VBPLV.n17 GND 0.20844f
C2233 VBPLV.t5 GND 0.23663f
C2234 VBPLV.n18 GND 0.20844f
C2235 VBPLV.t9 GND 0.23663f
C2236 VBPLV.n19 GND 0.20844f
C2237 VBPLV.t10 GND 0.23663f
C2238 VBPLV.n20 GND 0.20844f
C2239 VBPLV.t18 GND 0.23663f
C2240 VBPLV.n21 GND 0.20844f
C2241 decoder_3_0/decoder_2to4_2.bb[0].t1 GND 0.10871f
C2242 decoder_3_0/decoder_2to4_2.bb[0].n0 GND 0.1436f
C2243 decoder_3_0/decoder_2to4_2.bb[0].t2 GND 0.02955f
C2244 decoder_3_0/decoder_2to4_2.bb[0].t4 GND 0.04735f
C2245 decoder_3_0/decoder_2to4_2.bb[0].n1 GND 0.09326f
C2246 decoder_3_0/decoder_2to4_2.bb[0].n2 GND 0.04278f
C2247 decoder_3_0/decoder_2to4_2.bb[0].t3 GND 0.02955f
C2248 decoder_3_0/decoder_2to4_2.bb[0].t5 GND 0.04735f
C2249 decoder_3_0/decoder_2to4_2.bb[0].n3 GND 0.09323f
C2250 decoder_3_0/decoder_2to4_2.bb[0].n4 GND 0.03162f
C2251 decoder_3_0/decoder_2to4_2.bb[0].n5 GND 0.48141f
C2252 decoder_3_0/decoder_2to4_2.bb[0].n6 GND 6.01399f
C2253 decoder_3_0/decoder_2to4_2.bb[0].n7 GND 0.14712f
C2254 decoder_3_0/decoder_2to4_2.bb[0].t0 GND 0.07082f
C2255 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t2 GND 0.03812f
C2256 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t3 GND 0.03812f
C2257 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 GND 0.08766f
C2258 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 GND 0.1778f
C2259 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t6 GND 0.0394f
C2260 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t8 GND 0.06311f
C2261 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 GND 0.12033f
C2262 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 GND 0.07572f
C2263 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t7 GND 0.0394f
C2264 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t4 GND 0.06311f
C2265 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 GND 0.12036f
C2266 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 GND 0.03098f
C2267 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 GND 0.676f
C2268 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t5 GND 0.22836f
C2269 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 GND 10.4354f
C2270 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 GND 1.68228f
C2271 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 GND 0.03519f
C2272 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t0 GND 0.02478f
C2273 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t1 GND 0.02478f
C2274 lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 GND 0.05444f
C2275 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t1 GND 0.02431f
C2276 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t3 GND 0.02431f
C2277 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 GND 0.0534f
C2278 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 GND 0.03452f
C2279 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t5 GND 0.05817f
C2280 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t4 GND 0.03428f
C2281 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t8 GND 0.05817f
C2282 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t7 GND 0.03428f
C2283 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 GND 0.09761f
C2284 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 GND 0.1448f
C2285 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 GND 0.04367f
C2286 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t6 GND 0.03858f
C2287 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t10 GND 0.06183f
C2288 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 GND 0.12177f
C2289 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 GND 0.05586f
C2290 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t9 GND 0.03858f
C2291 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t12 GND 0.06183f
C2292 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 GND 0.12173f
C2293 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 GND 0.04128f
C2294 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 GND 0.64238f
C2295 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t11 GND 0.22403f
C2296 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 GND 9.2905f
C2297 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 GND 2.62797f
C2298 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 GND 0.0269f
C2299 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t0 GND 0.0374f
C2300 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t2 GND 0.0374f
C2301 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 GND 0.08599f
C2302 lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 GND 0.1744f
.ends

