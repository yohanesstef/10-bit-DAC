magic
tech sky130A
magscale 1 2
timestamp 1749005012
<< pwell >>
rect -307 -1083 307 1083
<< psubdiff >>
rect -271 1013 -175 1047
rect 175 1013 271 1047
rect -271 951 -237 1013
rect 237 951 271 1013
rect -271 -1013 -237 -951
rect 237 -1013 271 -951
rect -271 -1047 -175 -1013
rect 175 -1047 271 -1013
<< psubdiffcont >>
rect -175 1013 175 1047
rect -271 -951 -237 951
rect 237 -951 271 951
rect -175 -1047 175 -1013
<< xpolycontact >>
rect -141 485 141 917
rect -141 -917 141 -485
<< xpolyres >>
rect -141 -485 141 485
<< locali >>
rect -271 1013 -175 1047
rect 175 1013 271 1047
rect -271 951 -237 1013
rect 237 951 271 1013
rect -271 -1013 -237 -951
rect 237 -1013 271 -951
rect -271 -1047 -175 -1013
rect 175 -1047 271 -1013
<< viali >>
rect -125 502 125 899
rect -125 -899 125 -502
<< metal1 >>
rect -131 899 131 911
rect -131 502 -125 899
rect 125 502 131 899
rect -131 490 131 502
rect -131 -502 131 -490
rect -131 -899 -125 -502
rect 125 -899 131 -502
rect -131 -911 131 -899
<< properties >>
string FIXED_BBOX -254 -1030 254 1030
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 5.013 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 7.377k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
