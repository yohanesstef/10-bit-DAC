magic
tech sky130A
magscale 1 2
timestamp 1750003173
<< error_s >>
rect -440 1373 1250 1439
rect -440 -62 -374 1373
rect -314 1247 1124 1313
rect -314 -62 -248 1247
rect -220 1043 -214 1049
rect -226 1037 -220 1043
rect -7 0 23 1082
rect 59 60 89 1016
rect 721 60 751 1016
rect 59 56 375 60
rect 435 56 751 60
rect 787 0 817 1082
rect 0 -10 817 -6
rect -440 -128 -248 -62
rect 1058 -62 1124 1247
rect 1184 -62 1250 1373
rect 1058 -128 1250 -62
<< mvnsubdiff >>
rect -374 1313 1184 1373
rect -374 -62 -314 1313
rect 1124 -62 1184 1313
<< poly >>
rect -16 30 44 1113
rect 766 30 826 1113
<< locali >>
rect -361 1326 1171 1360
rect -361 -62 -327 1326
rect 1137 -62 1171 1326
<< metal1 >>
rect -280 1103 -220 1109
rect 148 1043 154 1103
rect 280 1043 286 1103
rect 323 1016 369 1126
rect 441 1016 487 1126
rect 524 1043 530 1103
rect 656 1043 662 1103
<< via1 >>
rect -280 1043 -220 1103
rect 154 1043 280 1103
rect 530 1043 656 1103
<< metal2 >>
rect -286 1043 -280 1103
rect -220 1043 154 1103
rect 280 1043 530 1103
rect 656 1043 662 1103
use sky130_fd_pr__pfet_g5v0d10v5_X66K38  sky130_fd_pr__pfet_g5v0d10v5_X66K38_0
timestamp 1749990477
transform 1 0 217 0 1 572
box -224 -582 224 544
use sky130_fd_pr__pfet_g5v0d10v5_X66K38  sky130_fd_pr__pfet_g5v0d10v5_X66K38_1
timestamp 1749990477
transform 1 0 593 0 1 572
box -224 -582 224 544
<< end >>
