* PEX produced on Fri Jun 27 22:11:25 WIB 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from top_rseg_n_dcell.ext - technology: sky130A

.subckt top_rseg_n_dcell DIN0 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 DIN9 ROUT VS1
+ VL2 VH2 VL3 VH3 VS4 SH[1] SH[2] SH[3] SH[4] VDD VDDH GND
X0 GND.t425 GND.t426 GND.t279 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X1 a_42781_10934.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t0 GND.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 top_segment_1_0.rseg_1_v3_1.v19.t0 top_segment_2_0.DEC2[1].t2 a_26719_5238.t0 GND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t3 VDD.t168 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_13061_17684.t0 top_segment_3_0.b[5].t2 a_15695_17684.t1 VDDH.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X5 a_18769_7938.t2 top_segment_4_1.bb3.t2 a_15714_6674.t4 VDDH.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X6 GND.t587 GND.t588 GND.t72 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X7 top_segment_2_0.rseg_2_v3_0.v42.t2 top_segment_2_0.rseg_2_v3_0.v41.t2 GND.t181 sky130_fd_pr__res_xhigh_po_1p41 l=5.32
X8 a_41787_17118.t1 top_segment_2_0.DEC2[2].t2 a_41529_17118.t1 VDDH.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X9 a_41714_2150.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t4 GND.t530 GND.t529 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 top_segment_2_0.rseg_2_v3_0.v4.t0 top_segment_2_0.rseg_2_v3_0.v5.t1 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=7.88
X11 top_segment_1_0.rseg_1_v3_1.v9.t1 top_segment_2_0.DEC2[0].t2 a_28603_6674.t4 GND.t352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X12 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X13 top_segment_2_0.rseg_2_v3_0.v10.t2 top_segment_2_0.DEC0[0].t2 a_19094_19162.t2 GND.t250 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X14 a_42781_13270.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t4 GND.t590 GND.t589 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X15 a_42245_11724.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t2 a_42271_12320.t0 VDDH.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X16 a_42781_9310.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t3 GND.t502 GND.t501 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X17 top_segment_1_0.rseg_1_v3_1.v56.t1 top_segment_2_0.DEC2[3].t2 a_28327_6674.t4 GND.t608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X18 VDDH.t23 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t6 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t3 VDDH.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X19 a_32181_7938.t2 top_segment_4_1.bb3.t3 a_26167_5238.t2 GND.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X20 top_segment_1_0.rseg_1_v3_1.v39.t1 top_segment_1_0.rseg_1_v3_1.v38.t0 GND.t72 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X21 a_43570_17828.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t4 GND.t528 GND.t527 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 VDD.t201 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t3 VDD.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t3 GND.t173 GND.t172 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_15143_17684.t1 top_segment_3_0.bb[6].t2 top_segment_3_0.rseg_3_v3_0.v2.t0 VDDH.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X25 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X26 VDD.t5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t1 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t5 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X28 top_segment_3_0.bb[4].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t2 GND.t459 GND.t458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X29 a_34580_9019.t2 top_segment_4_1.bb2.t2 a_31905_7938.t1 GND.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X30 GND.t368 GND.t369 GND.t122 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X31 top_segment_1_0.rseg_1_v3_1.v47.t0 top_segment_1_0.rseg_1_v3_1.v46.t0 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X32 GND.t461 GND.t462 GND.t21 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X33 a_13588_5238.t2 top_segment_4_1.DEC2.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t0 VDDH.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X34 a_34580_9019.t1 top_segment_4_1.b2.t2 a_32851_7938.t1 GND.t286 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X35 a_21596_17121.t5 top_segment_2_0.DEC2[2].t3 VL2.t1 GND.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X36 a_42271_15290.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t6 VDDH.t271 VDDH.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X37 a_35435_18538.t1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t4 GND.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X38 VDD.t118 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 VDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X39 a_19479_9019.t2 top_segment_4_1.bb2.t3 a_18217_7938.t1 VDDH.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X40 top_segment_1_0.rseg_1_v3_1.v49.t2 top_segment_1_0.rseg_1_v3_1.v50.t2 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X41 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t7 VDDH.t18 VDDH.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X42 VH3.t0 top_segment_4_1.b3.t2 a_16555_17684.t1 VDDH.t176 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X43 GND.t519 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 a_42609_17081.t0 GND.t518 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X44 top_segment_2_0.rseg_2_v3_0.v16.t1 top_segment_2_0.DEC0[0].t3 a_19922_19162.t2 GND.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X45 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t2 a_35957_18086.t1 GND.t429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X46 a_33724_9019.t0 top_segment_4_1.b2.t3 a_33679_7938.t0 GND.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X47 top_segment_1_0.rseg_1_v3_1.v27.t0 top_segment_2_0.DEC2[1].t3 a_29155_6674.t0 GND.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X48 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t4 VDD.t73 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X49 GND.t189 GND.t190 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X50 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t0 GND.t48 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X51 a_42271_14854.t1 a_42245_14694.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t1 VDDH.t274 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X52 a_18623_9019.t2 top_segment_4_1.bb2.t4 a_19045_7938.t1 VDDH.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X53 VDD.t180 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X54 GND.t353 top_segment_2_0.DEC2[0].t3 top_segment_4_1.DEC0.t0 GND.t339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X55 a_41529_17118.t0 top_segment_2_0.DEC2[1].t4 a_41271_17118.t0 VDDH.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X56 a_34000_9019.t1 top_segment_4_1.b1.t2 a_33420_9019.t2 GND.t403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X57 top_segment_1_0.rseg_1_v3_1.v9.t2 top_segment_1_0.rseg_1_v3_1.v10.t2 GND.t40 sky130_fd_pr__res_xhigh_po_1p41 l=2.19
X58 GND.t145 GND.t146 GND.t86 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X59 a_14416_5238.t3 top_segment_4_1.DEC1.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t1 VDDH.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X60 top_segment_3_0.b[5].t1 top_segment_3_0.bb[5].t2 GND.t276 GND.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X61 GND.t440 GND.t441 GND.t49 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X62 top_segment_1_0.rseg_1_v3_1.v35.t0 top_segment_1_0.rseg_1_v3_1.v36.t1 GND.t72 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X63 top_segment_1_0.rseg_1_v3_1.v19.t2 top_segment_1_0.rseg_1_v3_1.v18.t1 GND.t49 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X64 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t2 VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X65 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t0 top_segment_4_1.DEC1.t3 a_13900_6674.t1 VDDH.t124 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X66 a_42245_13704.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t7 a_42781_14260.t1 GND.t591 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X67 top_segment_4_1.bb2.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t3 VDDH.t4 VDDH.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X68 GND.t620 GND.t621 GND.t72 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X69 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t1 GND.t48 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X70 top_segment_2_0.rseg_2_v3_0.v6.t0 top_segment_2_0.rseg_2_v3_0.v5.t0 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=7.42
X71 VDD.t36 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t1 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X72 a_16831_17684.t0 top_segment_3_0.b[4].t2 a_13613_17684.t1 VDDH.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X73 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t4 a_43570_18104.t1 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X74 a_15714_6674.t0 top_segment_4_1.DEC0.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t1 VDDH.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X75 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t5 VDD.t185 VDD.t184 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X76 top_segment_1_0.rseg_1_v3_1.v25.t2 top_segment_1_0.rseg_1_v3_1.v26.t2 GND.t188 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X77 VDD.t222 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 VDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X78 VDD.t87 DIN7.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t3 VDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X79 top_segment_2_0.rseg_2_v3_0.v39.t2 top_segment_2_0.DEC0[2].t2 a_23510_19162.t2 GND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X80 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t4 VDD.t51 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X81 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t2 top_segment_4_1.DEC3.t2 a_13900_6674.t3 VDDH.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X82 top_segment_1_0.rseg_1_v3_1.v33.t1 top_segment_1_0.rseg_1_v3_1.v34.t0 GND.t72 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X83 top_segment_2_0.rseg_2_v3_0.v12.t2 top_segment_2_0.rseg_2_v3_0.v13.t2 GND.t21 sky130_fd_pr__res_xhigh_po_1p41 l=5.58
X84 top_segment_2_0.DEC1[0].t1 top_segment_2_0.DEC1[3].t2 a_41787_18542.t1 VDDH.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X85 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t5 VDD.t223 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X86 top_segment_3_0.rseg_3_v3_0.v4.t0 top_segment_3_0.rseg_3_v3_0.v5.t0 GND.t23 sky130_fd_pr__res_xhigh_po_1p41 l=3.53
X87 top_segment_1_0.rseg_1_v3_1.v50.t1 top_segment_2_0.DEC2[3].t3 a_26443_5238.t4 GND.t609 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X88 GND.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 a_42609_20641.t1 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X89 top_segment_4_1.b3.t1 top_segment_4_1.bb3.t4 VDDH.t101 VDDH.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X90 VDDH.t168 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t7 a_42271_11884.t0 VDDH.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X91 a_42802_2702.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t4 GND.t478 GND.t477 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X92 GND.t597 GND.t598 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X93 top_segment_1_0.rseg_1_v3_1.v2.t2 top_segment_2_0.DEC2[0].t4 a_26443_5238.t3 GND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X94 top_segment_2_0.rseg_2_v3_0.v44.t0 top_segment_2_0.rseg_2_v3_0.v43.t1 GND.t181 sky130_fd_pr__res_xhigh_po_1p41 l=5.58
X95 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t2 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X96 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t1 VDDH.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X97 a_27429_5238.t4 top_segment_2_0.DEC2[3].t4 top_segment_1_0.rseg_1_v3_1.v53.t2 GND.t610 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X98 a_42781_5984.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t0 GND.t592 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X99 top_segment_2_0.rseg_2_v3_0.v26.t1 top_segment_2_0.rseg_2_v3_0.v25.t1 GND.t122 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X100 a_14416_5238.t0 top_segment_4_1.b3.t3 a_19045_7938.t0 VDDH.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X101 GND.t364 GND.t365 GND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=3.94
X102 a_42609_19573.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 GND.t80 GND.t79 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X103 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t1 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X104 top_segment_1_0.rseg_1_v3_1.v34.t2 top_segment_2_0.DEC2[2].t4 a_26443_5238.t1 GND.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X105 top_segment_2_0.rseg_2_v3_0.v8.t0 top_segment_2_0.rseg_2_v3_0.v7.t0 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=6.65
X106 VDD.t22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t1 VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X107 a_42245_15684.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t2 a_42271_16280.t1 VDDH.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X108 a_43890_3610.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t7 a_43890_3526.t1 GND.t113 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X109 top_segment_1_0.rseg_1_v3_1.v31.t2 top_segment_1_0.rseg_1_v3_1.v32.t2 GND.t188 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X110 top_segment_3_0.rseg_3_v3_0.v12.t2 top_segment_3_0.rseg_3_v3_0.v13.t0 GND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=4.6
X111 a_14452_6674.t4 top_segment_4_1.bb3.t5 a_17823_7938.t2 VDDH.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X112 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t1 GND.t192 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X113 top_segment_2_0.rseg_2_v3_0.v2.t1 top_segment_2_0.rseg_2_v3_0.v1.t0 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=10.24
X114 a_42609_20997.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 GND.t422 GND.t421 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X115 a_18099_7938.t1 top_segment_4_1.b3.t4 a_13154_5238.t0 VDDH.t71 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X116 top_segment_1_0.rseg_1_v3_1.v18.t0 top_segment_2_0.DEC2[1].t5 a_26443_5238.t0 GND.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X117 a_41938_2314.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t5 a_41938_2230.t0 GND.t78 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X118 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t0 DIN7.t1 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X119 VDD.t7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t1 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X120 top_segment_1_0.rseg_1_v3_1.v42.t2 top_segment_2_0.DEC2[2].t5 a_28879_6674.t2 GND.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X121 GND.t611 top_segment_2_0.DEC2[3].t5 top_segment_4_1.DEC3.t0 GND.t339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X122 a_18493_7938.t2 top_segment_4_1.bb3.t6 a_15438_6674.t4 VDDH.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X123 VDDH.t266 VDDH.t264 VDDH.t265 VDDH.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X124 a_27429_5238.t0 top_segment_2_0.DEC2[1].t6 top_segment_1_0.rseg_1_v3_1.v21.t0 GND.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X125 top_segment_2_0.rseg_2_v3_0.v22.t0 top_segment_2_0.rseg_2_v3_0.v23.t0 GND.t8 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X126 a_41787_17802.t0 top_segment_2_0.DEC2[1].t7 a_41529_17802.t0 VDDH.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X127 VDD.t72 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t0 VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X128 top_segment_2_0.rseg_2_v3_0.v40.t0 top_segment_2_0.rseg_2_v3_0.v41.t1 GND.t324 sky130_fd_pr__res_xhigh_po_1p41 l=5.22
X129 top_segment_2_0.rseg_2_v3_0.v36.t1 top_segment_2_0.rseg_2_v3_0.v35.t1 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X130 top_segment_1_0.rseg_1_v3_1.v8.t1 top_segment_2_0.DEC2[0].t5 a_28327_6674.t3 GND.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X131 VDD.t120 DIN6.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t1 VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X132 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t5 a_43890_2518.t1 GND.t392 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X133 a_41787_20308.t1 top_segment_2_0.DEC0[2].t3 a_41529_20308.t1 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X134 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t2 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X135 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t3 DIN4.t0 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X136 top_segment_1_0.rseg_1_v3_1.v7.t2 top_segment_1_0.rseg_1_v3_1.v8.t2 GND.t86 sky130_fd_pr__res_xhigh_po_1p41 l=2.5
X137 top_segment_1_0.rseg_1_v3_1.v19.t1 top_segment_1_0.rseg_1_v3_1.v20.t1 GND.t49 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X138 top_segment_1_0.rseg_1_v3_1.v47.t2 top_segment_1_0.rseg_1_v3_1.v48.t1 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X139 top_segment_2_0.DEC2[1].t1 top_segment_2_0.DEC2[3].t6 a_41787_17460.t1 VDDH.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X140 a_32851_7938.t0 top_segment_4_1.b3.t5 a_29589_6674.t1 GND.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X141 top_segment_2_0.rseg_2_v3_0.v34.t1 top_segment_2_0.rseg_2_v3_0.v33.t1 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X142 top_segment_2_0.rseg_2_v3_0.v30.t0 top_segment_2_0.DEC0[1].t2 a_19646_19162.t0 GND.t468 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X143 a_41271_19226.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t6 VDDH.t42 VDDH.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X144 top_segment_2_0.rseg_2_v3_0.v42.t0 top_segment_2_0.DEC0[2].t4 a_19094_19162.t0 GND.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X145 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t4 a_43890_3610.t0 GND.t158 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X146 top_segment_3_0.b[6].t1 top_segment_3_0.bb[6].t3 VDDH.t212 VDDH.t211 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X147 a_18217_7938.t2 top_segment_4_1.bb3.t7 a_15162_6674.t4 VDDH.t104 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X148 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t5 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X149 a_43890_3526.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t5 GND.t139 GND.t138 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X150 a_13645_18854.t2 top_segment_3_0.b[6].t2 top_segment_4_1.V0.t3 VDDH.t306 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X151 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t0 GND.t48 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X152 a_22176_17121.t3 top_segment_2_0.DEC2[0].t6 VH2.t2 GND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X153 a_19479_9019.t0 top_segment_4_1.b2.t4 a_17271_7938.t0 VDDH.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X154 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t6 a_42802_2150.t1 GND.t140 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X155 GND.t211 GND.t212 GND.t122 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X156 top_segment_2_0.V0.t0 top_segment_2_0.DEC0[0].t4 a_22406_19162.t2 GND.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X157 a_34000_9019.t0 top_segment_4_1.b2.t5 a_33403_7938.t0 GND.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X158 top_segment_3_0.rseg_3_v3_0.v10.t1 top_segment_3_0.rseg_3_v3_0.v9.t1 GND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=4.09
X159 GND.t472 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t4 a_42781_10934.t1 GND.t471 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X160 top_segment_1_0.rseg_1_v3_1.v26.t0 top_segment_2_0.DEC2[1].t8 a_28879_6674.t0 GND.t570 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X161 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t5 VDD.t150 VDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X162 a_18899_9019.t2 top_segment_4_1.bb2.t5 a_18769_7938.t0 VDDH.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X163 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t2 a_35435_18774.t1 GND.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X164 a_42245_8754.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t9 a_42781_9310.t0 GND.t593 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X165 VDD.t152 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t0 VDD.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X166 GND.t182 GND.t183 GND.t49 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X167 a_18899_9019.t1 top_segment_4_1.bb1.t2 a_18319_9019.t1 VDDH.t188 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X168 a_33724_9019.t1 top_segment_4_1.b1.t3 a_33116_9019.t2 GND.t404 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X169 a_41529_17802.t1 top_segment_2_0.DEC2[0].t7 a_41271_17802.t1 VDDH.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X170 top_segment_1_0.rseg_1_v3_1.v59.t2 top_segment_1_0.rseg_1_v3_1.v60.t2 GND.t201 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X171 top_segment_2_0.rseg_2_v3_0.v9.t1 top_segment_2_0.DEC0[0].t5 a_21026_19162.t1 GND.t538 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X172 GND.t10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t3 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X173 a_43890_2518.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t7 GND.t418 GND.t417 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X174 a_29865_6674.t0 top_segment_2_0.DEC2[1].t9 top_segment_1_0.rseg_1_v3_1.v29.t0 GND.t571 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X175 top_segment_2_0.rseg_2_v3_0.v29.t0 top_segment_2_0.DEC0[1].t3 a_20474_19162.t0 GND.t469 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X176 a_41529_20308.t0 top_segment_2_0.DEC0[0].t6 a_41271_20308.t0 VDDH.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X177 VDD.t145 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t0 VDD.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X178 GND.t414 DIN1.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t3 GND.t413 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X179 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t1 GND.t187 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X180 a_14140_5238.t3 top_segment_4_1.DEC1.t4 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t1 VDDH.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X181 a_41787_19568.t1 top_segment_2_0.DEC1[1].t2 a_41529_19568.t0 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X182 a_42271_8360.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t8 VDDH.t170 VDDH.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X183 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t5 VDD.t181 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X184 VDDH.t172 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t9 a_42271_15844.t1 VDDH.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X185 VDD.t91 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t1 VDD.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X186 GND.t205 DIN4.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t0 GND.t204 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X187 top_segment_1_0.rseg_1_v3_1.v17.t2 top_segment_1_0.rseg_1_v3_1.v18.t2 GND.t49 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X188 GND.t164 GND.t165 GND.t21 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X189 a_13495_17684.t2 top_segment_3_0.b[6].t3 top_segment_3_0.rseg_3_v3_0.v13.t2 VDDH.t307 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X190 a_15438_6674.t3 top_segment_4_1.DEC0.t3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t1 VDDH.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X191 GND.t362 GND.t363 GND.t192 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X192 VDD.t214 DIN0.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t1 VDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X193 SH[2].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t2 VDDH.t302 VDDH.t301 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X194 top_segment_2_0.rseg_2_v3_0.v26.t0 top_segment_2_0.DEC0[1].t4 a_19094_19162.t3 GND.t470 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X195 VDD.t196 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t0 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X196 top_segment_1_0.rseg_1_v3_1.v49.t0 top_segment_1_0.rseg_1_v3_1.v48.t0 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X197 a_42609_17081.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t6 top_segment_2_0.DEC2[0].t1 GND.t432 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X198 a_42781_9944.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t0 GND.t594 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X199 a_42271_7924.t1 a_42245_7764.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t1 VDDH.t197 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X200 a_13864_5238.t2 top_segment_4_1.DEC2.t3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t1 VDDH.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X201 a_21854_19162.t3 top_segment_2_0.DEC1[1].t3 a_20740_17121.t2 GND.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X202 a_27153_5238.t2 top_segment_4_1.bb3.t8 a_32851_7938.t2 GND.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X203 a_18015_9019.t1 top_segment_4_1.bb0.t2 VS4.t1 VDDH.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X204 top_segment_1_0.rseg_1_v3_1.v1.t0 GND.t87 GND.t86 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X205 GND.t134 GND.t135 GND.t48 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X206 VDD.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X207 GND.t342 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t2 a_42781_7964.t1 GND.t341 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X208 a_41271_18144.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t7 VDDH.t290 VDDH.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X209 top_segment_2_0.rseg_2_v3_0.v4.t1 top_segment_2_0.DEC0[0].t7 a_21854_19162.t1 GND.t539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X210 a_27981_5238.t2 top_segment_4_1.bb3.t9 a_33679_7938.t2 GND.t535 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X211 a_15714_6674.t2 top_segment_4_1.DEC2.t4 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t0 VDDH.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X212 VDD.t172 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t0 VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X213 top_segment_1_0.rseg_1_v3_1.v33.t0 top_segment_1_0.rseg_1_v3_1.v32.t0 GND.t72 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X214 GND.t315 GND.t316 GND.t23 sky130_fd_pr__res_xhigh_po_1p41 l=3.83
X215 a_43570_18700.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t6 GND.t406 GND.t405 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X216 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t5 GND.t198 GND.t197 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X217 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t0 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X218 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t6 VDD.t212 VDD.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X219 top_segment_1_0.rseg_1_v3_1.v25.t1 top_segment_1_0.rseg_1_v3_1.v24.t2 GND.t188 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X220 top_segment_1_0.rseg_1_v3_1.v1.t2 top_segment_2_0.DEC2[0].t8 a_26167_5238.t3 GND.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X221 top_segment_2_0.rseg_2_v3_0.v10.t0 top_segment_2_0.rseg_2_v3_0.v11.t1 GND.t21 sky130_fd_pr__res_xhigh_po_1p41 l=5.94
X222 top_segment_1_0.rseg_1_v3_1.v53.t1 top_segment_1_0.rseg_1_v3_1.v52.t0 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X223 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t1 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X224 a_42781_10300.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t4 GND.t261 GND.t260 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X225 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t1 GND.t149 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X226 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t4 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X227 VDD.t99 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t1 VDD.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X228 a_41938_2230.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t7 a_41938_2146.t0 GND.t407 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X229 a_27153_5238.t3 top_segment_2_0.DEC2[0].t9 top_segment_1_0.rseg_1_v3_1.v4.t1 GND.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X230 top_segment_2_0.rseg_2_v3_0.v46.t2 top_segment_2_0.DEC0[2].t5 a_19646_19162.t3 GND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X231 a_41529_19568.t1 top_segment_2_0.DEC1[0].t2 a_41271_19568.t1 VDDH.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X232 a_13645_18854.t1 top_segment_3_0.bb[5].t3 a_14165_17684.t1 VDDH.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X233 a_22682_19162.t2 top_segment_2_0.DEC1[1].t4 a_22176_17121.t1 GND.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X234 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t6 VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X235 SH[4].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t2 GND.t117 GND.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X236 a_15990_6674.t3 top_segment_4_1.DEC0.t4 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t1 VDDH.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X237 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t7 GND.t142 GND.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X238 top_segment_2_0.rseg_2_v3_0.v24.t1 top_segment_2_0.rseg_2_v3_0.v25.t0 GND.t122 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X239 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t0 DIN0.t1 VDD.t216 VDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X240 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t8 VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X241 top_segment_1_0.rseg_1_v3_1.v45.t0 top_segment_1_0.rseg_1_v3_1.v46.t1 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X242 GND.t266 GND.t267 GND.t149 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X243 top_segment_1_0.rseg_1_v3_1.v17.t0 top_segment_2_0.DEC2[1].t10 a_26167_5238.t0 GND.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X244 top_segment_2_0.rseg_2_v3_0.v8.t2 top_segment_2_0.rseg_2_v3_0.v9.t2 GND.t21 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X245 a_35435_18538.t2 a_35435_18774.t6 GND.t467 GND.t465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X246 a_16831_17684.t2 top_segment_3_0.bb[4].t2 a_14165_17684.t2 VDDH.t277 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X247 top_segment_4_1.bb1.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t2 GND.t596 GND.t595 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X248 GND.t396 DIN9.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t0 GND.t395 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X249 VDD.t11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X250 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t1 DIN3.t0 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X251 top_segment_1_0.rseg_1_v3_1.v48.t2 top_segment_2_0.DEC2[3].t7 a_25891_5238.t4 GND.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X252 top_segment_2_0.rseg_2_v3_0.v18.t1 top_segment_2_0.rseg_2_v3_0.v19.t2 GND.t8 sky130_fd_pr__res_xhigh_po_1p41 l=4.96
X253 top_segment_2_0.rseg_2_v3_0.v16.t3 top_segment_2_0.DEC0[1].t5 a_22406_19162.t0 GND.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X254 a_17823_7938.t1 top_segment_4_1.b3.t6 a_12878_5238.t0 VDDH.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X255 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t7 VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X256 a_43570_18976.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t9 GND.t582 GND.t270 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X257 a_42271_12320.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t10 VDDH.t174 VDDH.t173 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X258 top_segment_1_0.rseg_1_v3_1.v57.t0 top_segment_1_0.rseg_1_v3_1.v58.t1 GND.t201 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X259 top_segment_3_0.rseg_3_v3_0.v14.t1 top_segment_3_0.rseg_3_v3_0.v13.t1 GND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X260 a_15714_6674.t1 top_segment_4_1.DEC1.t5 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t0 VDDH.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X261 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t0 GND.t149 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X262 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t2 top_segment_4_1.DEC3.t3 a_13154_5238.t1 VDDH.t192 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X263 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t5 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t5 VDDH.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X264 top_segment_1_0.rseg_1_v3_1.v5.t1 top_segment_1_0.rseg_1_v3_1.v4.t2 GND.t86 sky130_fd_pr__res_xhigh_po_1p41 l=3.12
X265 a_14416_5238.t4 top_segment_4_1.DEC0.t5 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t1 VDDH.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X266 top_segment_3_0.rseg_3_v3_0.v12.t1 top_segment_3_0.rseg_3_v3_0.v11.t1 GND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=4.45
X267 a_42245_8754.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t3 a_42271_9350.t1 VDDH.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X268 a_13864_5238.t0 top_segment_4_1.b3.t7 a_18493_7938.t0 VDDH.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X269 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t2 VDDH.t26 VDDH.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X270 top_segment_1_0.rseg_1_v3_1.v32.t1 top_segment_2_0.DEC2[2].t6 a_25891_5238.t1 GND.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X271 top_segment_2_0.rseg_2_v3_0.v25.t2 top_segment_2_0.DEC0[1].t6 a_21026_19162.t0 GND.t648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X272 a_42781_7330.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t2 GND.t19 GND.t18 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X273 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t7 a_43570_18976.t0 GND.t505 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X274 a_41938_3162.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t5 GND.t263 GND.t262 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X275 VDD.t102 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t2 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X276 a_14140_5238.t1 top_segment_4_1.DEC3.t4 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t2 VDDH.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X277 GND.t232 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t6 a_42781_14894.t1 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X278 top_segment_4_1.b2.t0 top_segment_4_1.bb2.t6 GND.t228 GND.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X279 a_13900_6674.t4 top_segment_4_1.bb3.t10 a_17271_7938.t2 VDDH.t283 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X280 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t4 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X281 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t8 a_41714_2426.t0 GND.t506 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X282 a_14867_17684.t2 top_segment_3_0.b[6].t4 top_segment_3_0.rseg_3_v3_0.v11.t2 VDDH.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X283 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t6 a_43570_20400.t1 GND.t523 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X284 a_16279_17684.t0 top_segment_3_0.b[4].t3 a_13061_17684.t1 VDDH.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X285 a_41938_2146.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t7 GND.t613 GND.t612 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X286 top_segment_2_0.DEC0[2].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t2 a_41787_20650.t1 VDDH.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X287 a_29155_6674.t1 top_segment_4_1.b3.t8 a_32733_7938.t0 GND.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X288 a_42245_10734.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t11 a_42781_11290.t0 GND.t356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X289 GND.t54 GND.t55 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X290 top_segment_2_0.rseg_2_v3_0.v21.t1 top_segment_2_0.DEC0[1].t7 a_23234_19162.t0 GND.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X291 GND.t380 GND.t381 GND.t86 sky130_fd_pr__res_xhigh_po_1p41 l=2.5
X292 a_43570_20124.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t3 GND.t169 GND.t168 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X293 a_13771_17684.t1 top_segment_3_0.bb[5].t4 a_13613_17684.t2 VDDH.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X294 a_22958_19162.t2 top_segment_2_0.DEC1[1].t5 a_21016_17121.t3 GND.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X295 top_segment_2_0.rseg_2_v3_0.v47.t2 top_segment_2_0.DEC0[2].t6 a_20198_19162.t3 GND.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X296 a_33403_7938.t1 top_segment_4_1.b3.t9 a_30141_6674.t1 GND.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X297 a_41787_19966.t0 top_segment_2_0.DEC0[2].t7 a_41529_19966.t1 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X298 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t4 GND.t331 GND.t330 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X299 GND.t584 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t3 GND.t583 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X300 top_segment_1_0.rseg_1_v3_1.v35.t1 top_segment_1_0.rseg_1_v3_1.v34.t1 GND.t72 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X301 GND.t296 DIN3.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t3 GND.t295 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X302 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t7 GND.t234 GND.t233 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X303 a_34304_9019.t2 top_segment_4_1.bb2.t7 a_32181_7938.t0 GND.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X304 top_segment_1_0.rseg_1_v3_1.v25.t0 top_segment_2_0.DEC2[1].t11 a_28603_6674.t0 GND.t476 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X305 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t0 DIN1.t1 GND.t240 GND.t239 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X306 top_segment_1_0.rseg_1_v3_1.v55.t1 top_segment_1_0.rseg_1_v3_1.v54.t1 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X307 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t8 VDDH.t19 VDDH.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X308 top_segment_2_0.rseg_2_v3_0.v20.t1 top_segment_2_0.DEC0[1].t8 a_21854_19162.t0 GND.t649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X309 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t2 top_segment_4_1.DEC1.t6 a_12878_5238.t3 VDDH.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X310 a_42271_12874.t1 a_42245_12714.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t1 VDDH.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X311 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t8 a_43570_19252.t1 GND.t614 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X312 a_42781_11924.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t0 GND.t357 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X313 VDDH.t82 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t11 a_42271_7924.t0 VDDH.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X314 a_41714_3622.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t8 GND.t185 GND.t184 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X315 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t0 GND.t11 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X316 top_segment_3_0.rseg_3_v3_0.v6.t1 top_segment_3_0.rseg_3_v3_0.v7.t1 GND.t23 sky130_fd_pr__res_xhigh_po_1p41 l=3.68
X317 top_segment_4_1.b0.t1 top_segment_4_1.bb0.t3 VDDH.t50 VDDH.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X318 a_15695_17684.t0 top_segment_3_0.b[6].t5 top_segment_3_0.rseg_3_v3_0.v8.t3 VDDH.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X319 a_13613_17684.t0 top_segment_3_0.b[5].t3 a_15143_17684.t2 VDDH.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X320 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t3 VDD.t75 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X321 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t8 VDD.t135 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X322 a_41271_18542.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t8 VDDH.t291 VDDH.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X323 a_20474_19162.t2 top_segment_2_0.DEC1[0].t3 a_22176_17121.t4 GND.t510 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X324 a_18623_9019.t0 top_segment_4_1.bb1.t3 a_18015_9019.t0 VDDH.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X325 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t3 VDD.t131 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X326 top_segment_1_0.rseg_1_v3_1.v3.t1 top_segment_1_0.rseg_1_v3_1.v2.t1 GND.t86 sky130_fd_pr__res_xhigh_po_1p41 l=3.73
X327 top_segment_3_0.rseg_3_v3_0.v8.t1 top_segment_3_0.rseg_3_v3_0.v9.t0 GND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=3.94
X328 top_segment_3_0.V0.t3 top_segment_2_0.DEC0[2].t8 a_19922_19162.t0 GND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X329 a_41714_2426.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t9 GND.t485 GND.t484 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X330 a_23510_19162.t0 top_segment_2_0.DEC1[2].t2 a_21016_17121.t0 GND.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X331 top_segment_2_0.rseg_2_v3_0.v41.t0 top_segment_2_0.DEC0[2].t9 a_21026_19162.t2 GND.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X332 a_42781_14260.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t6 GND.t90 GND.t89 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X333 top_segment_1_0.rseg_1_v3_1.v45.t2 top_segment_1_0.rseg_1_v3_1.v44.t1 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X334 a_42609_18861.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t7 top_segment_2_0.DEC1[1].t0 GND.t270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X335 a_42245_12714.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t2 a_42271_13310.t1 VDDH.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X336 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t0 top_segment_4_1.DEC2.t5 a_14452_6674.t1 VDDH.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X337 top_segment_1_0.rseg_1_v3_1.v24.t0 top_segment_2_0.DEC2[1].t12 a_28327_6674.t0 GND.t378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X338 top_segment_1_0.rseg_1_v3_1.v17.t1 top_segment_1_0.rseg_1_v3_1.v16.t1 GND.t49 sky130_fd_pr__res_xhigh_po_1p41 l=1.58
X339 VDD.t199 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t2 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X340 top_segment_2_0.rseg_2_v3_0.v5.t2 top_segment_2_0.DEC0[0].t8 a_23234_19162.t1 GND.t540 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X341 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t5 GND.t160 GND.t159 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X342 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t2 top_segment_4_1.DEC1.t7 a_12602_5238.t3 VDDH.t199 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X343 top_segment_2_0.rseg_2_v3_0.v17.t0 top_segment_2_0.DEC0[1].t9 a_22682_19162.t0 GND.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X344 a_15438_6674.t1 top_segment_4_1.DEC2.t6 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t1 VDDH.t138 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X345 top_segment_1_0.rseg_1_v3_1.v51.t1 top_segment_1_0.rseg_1_v3_1.v52.t1 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X346 a_41529_19966.t0 top_segment_2_0.DEC0[1].t10 a_41271_19966.t0 VDDH.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X347 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t2 top_segment_4_1.DEC0.t6 a_13900_6674.t2 VDDH.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X348 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t7 a_43026_2242.t0 GND.t578 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X349 a_14140_5238.t2 top_segment_4_1.DEC2.t7 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t2 VDDH.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X350 top_segment_3_0.bb[5].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t2 GND.t39 GND.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X351 a_13588_5238.t4 top_segment_4_1.DEC1.t8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t2 VDDH.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X352 GND.t619 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 a_42609_17793.t0 GND.t618 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X353 a_42609_17437.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 GND.t265 GND.t264 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X354 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t1 GND.t192 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X355 top_segment_2_0.DEC2[0].t0 top_segment_2_0.DEC2[3].t8 a_41787_17118.t0 VDDH.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X356 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t7 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t1 VDDH.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X357 a_41787_18884.t0 top_segment_2_0.DEC1[2].t3 a_41529_18884.t0 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X358 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t2 top_segment_4_1.DEC0.t7 a_14728_6674.t3 VDDH.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X359 GND.t616 GND.t617 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X360 a_42271_16280.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t12 VDDH.t84 VDDH.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X361 VDD.t173 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t2 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X362 top_segment_2_0.rseg_2_v3_0.v10.t1 top_segment_2_0.rseg_2_v3_0.v9.t0 GND.t21 sky130_fd_pr__res_xhigh_po_1p41 l=6.14
X363 top_segment_2_0.rseg_2_v3_0.v12.t1 top_segment_2_0.DEC0[0].t9 a_19370_19162.t1 GND.t541 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X364 top_segment_2_0.rseg_2_v3_0.v32.t1 top_segment_2_0.rseg_2_v3_0.v33.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X365 a_42271_15844.t0 a_42245_15684.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t1 VDDH.t164 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X366 GND.t508 GND.t509 GND.t188 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X367 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t0 GND.t44 sky130_fd_pr__res_xhigh_po_1p41 l=1.94
X368 a_15419_17684.t0 top_segment_3_0.bb[6].t4 top_segment_3_0.rseg_3_v3_0.v1.t0 VDDH.t213 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X369 VL3.t1 top_segment_4_1.bb3.t11 a_16555_17684.t2 VDDH.t284 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X370 a_42781_14894.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t0 GND.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X371 top_segment_2_0.rseg_2_v3_0.v43.t2 top_segment_2_0.DEC0[2].t10 a_20750_19162.t2 GND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X372 a_41271_17460.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t9 VDDH.t292 VDDH.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X373 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t8 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t5 VDDH.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X374 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t9 VDD.t137 VDD.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X375 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t8 VDD.t204 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X376 a_17547_7938.t1 top_segment_4_1.b3.t10 a_12602_5238.t0 VDDH.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X377 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t9 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X378 top_segment_1_0.rseg_1_v3_1.v16.t0 top_segment_2_0.DEC2[1].t13 a_25891_5238.t0 GND.t379 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X379 a_13771_17684.t0 top_segment_3_0.bb[6].t5 top_segment_3_0.rseg_3_v3_0.v6.t0 VDDH.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X380 a_42245_14694.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t14 a_42781_15250.t0 GND.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X381 top_segment_4_1.bb3.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t3 VDDH.t11 VDDH.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X382 top_segment_1_0.rseg_1_v3_1.v40.t2 top_segment_2_0.DEC2[2].t7 a_28327_6674.t2 GND.t310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X383 GND.t580 top_segment_2_0.DEC2[1].t14 top_segment_4_1.DEC1.t0 GND.t339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X384 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t2 top_segment_4_1.DEC3.t5 a_12878_5238.t1 VDDH.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X385 top_segment_2_0.rseg_2_v3_0.v38.t0 top_segment_2_0.rseg_2_v3_0.v39.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=5.01
X386 a_13588_5238.t0 top_segment_4_1.b3.t11 a_18217_7938.t0 VDDH.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X387 VDDH.t263 VDDH.t261 VDDH.t262 VDDH.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X388 top_segment_2_0.rseg_2_v3_0.v35.t2 top_segment_2_0.DEC0[2].t11 a_22958_19162.t3 GND.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X389 top_segment_1_0.rseg_1_v3_1.v59.t0 top_segment_1_0.rseg_1_v3_1.v58.t0 GND.t201 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X390 a_42245_5784.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t15 a_42781_6340.t0 GND.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X391 top_segment_2_0.rseg_2_v3_0.v2.t0 top_segment_2_0.rseg_2_v3_0.v3.t0 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=9.22
X392 a_37219_19465.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t8 GND.t272 GND.t271 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1769 pd=1.8 as=0.1769 ps=1.8 w=0.61 l=9.7
X393 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t2 GND.t149 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X394 a_13864_5238.t1 top_segment_4_1.DEC3.t6 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t1 VDDH.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X395 a_42609_20285.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t9 top_segment_2_0.DEC0[1].t1 GND.t202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X396 a_41529_18884.t1 top_segment_2_0.DEC1[0].t4 a_41271_18884.t1 VDDH.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X397 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t1 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=1.63
X398 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t10 VDD.t138 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X399 a_28879_6674.t1 top_segment_4_1.b3.t12 a_32457_7938.t0 GND.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X400 top_segment_2_0.rseg_2_v3_0.v38.t2 top_segment_2_0.DEC0[2].t12 a_21578_19162.t3 GND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X401 a_23234_19162.t2 top_segment_2_0.DEC1[2].t4 a_22176_17121.t2 GND.t410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X402 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t2 top_segment_4_1.DEC0.t8 a_12878_5238.t4 VDDH.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X403 top_segment_3_0.b[4].t1 top_segment_3_0.bb[4].t3 VDDH.t279 VDDH.t278 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X404 VDDH.t86 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t13 a_42271_12874.t0 VDDH.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X405 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t2 GND.t44 sky130_fd_pr__res_xhigh_po_1p41 l=2.4
X406 a_43026_3242.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t4 a_43026_3158.t1 GND.t50 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X407 a_42802_3602.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t3 a_42802_3518.t0 GND.t507 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X408 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t0 GND.t11 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X409 top_segment_3_0.rseg_3_v3_0.v2.t2 top_segment_3_0.rseg_3_v3_0.v3.t2 GND.t23 sky130_fd_pr__res_xhigh_po_1p41 l=3.32
X410 a_37853_19465.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t5 GND.t256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X411 a_33127_7938.t1 top_segment_4_1.b3.t13 a_29865_6674.t1 GND.t209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X412 a_13864_5238.t4 top_segment_4_1.DEC0.t9 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t2 VDDH.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X413 a_42781_6974.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t0 GND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X414 top_segment_2_0.rseg_2_v3_0.v42.t1 top_segment_2_0.rseg_2_v3_0.v43.t0 GND.t181 sky130_fd_pr__res_xhigh_po_1p41 l=5.47
X415 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t2 GND.t44 sky130_fd_pr__res_xhigh_po_1p41 l=1.78
X416 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t0 GND.t192 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X417 VDD.t154 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t0 VDD.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X418 a_13588_5238.t3 top_segment_4_1.DEC3.t7 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t0 VDDH.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X419 top_segment_3_0.rseg_3_v3_0.v8.t2 top_segment_3_0.rseg_3_v3_0.v7.t2 GND.t23 sky130_fd_pr__res_xhigh_po_1p41 l=3.83
X420 a_35435_18774.t0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t1 GND.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X421 top_segment_1_0.rseg_1_v3_1.v53.t0 top_segment_1_0.rseg_1_v3_1.v54.t0 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X422 VDD.t104 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 VDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X423 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t8 a_43570_17276.t1 GND.t235 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X424 top_segment_2_0.rseg_2_v3_0.v32.t3 top_segment_2_0.DEC0[2].t13 a_22406_19162.t3 GND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X425 a_21026_19162.t3 top_segment_2_0.DEC1[3].t3 a_22176_17121.t5 GND.t645 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X426 a_41394_3894.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t1 VDD.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X427 a_35957_18086.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t5 GND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X428 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t2 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X429 top_segment_3_0.bb[6].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t3 VDDH.t47 VDDH.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X430 top_segment_1_0.rseg_1_v3_1.v11.t0 top_segment_1_0.rseg_1_v3_1.v12.t0 GND.t40 sky130_fd_pr__res_xhigh_po_1p41 l=1.99
X431 a_42609_17793.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t10 top_segment_2_0.DEC2[2].t1 GND.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X432 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t0 top_segment_4_1.DEC2.t8 a_12326_5238.t2 VDDH.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X433 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t4 a_43026_3242.t0 GND.t292 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X434 a_41394_2698.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t0 VDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X435 a_43026_2242.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t11 GND.t214 GND.t213 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X436 top_segment_1_0.rseg_1_v3_1.v55.t0 top_segment_1_0.rseg_1_v3_1.v56.t0 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X437 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t4 GND.t504 GND.t503 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X438 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t3 a_42802_3602.t1 GND.t479 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X439 top_segment_3_0.rseg_3_v3_0.v6.t2 top_segment_3_0.rseg_3_v3_0.v5.t2 GND.t23 sky130_fd_pr__res_xhigh_po_1p41 l=3.58
X440 a_43026_3158.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t4 GND.t92 GND.t91 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X441 SH[1].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t2 GND.t200 GND.t199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X442 a_42802_3518.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t3 a_42802_3434.t0 GND.t520 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X443 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t1 top_segment_4_1.DEC1.t9 a_12326_5238.t3 VDDH.t201 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X444 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t10 VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X445 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t1 top_segment_4_1.DEC2.t9 a_13154_5238.t2 VDDH.t127 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X446 a_43570_18104.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t5 GND.t153 GND.t152 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X447 a_33116_9019.t0 top_segment_4_1.b0.t2 VS1.t1 GND.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X448 VDD.t124 DIN9.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t1 VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X449 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t9 VDD.t206 VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X450 a_30417_6674.t3 top_segment_2_0.DEC2[0].t10 top_segment_1_0.rseg_1_v3_1.v15.t2 GND.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X451 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t2 GND.t149 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X452 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t2 top_segment_4_1.DEC1.t10 a_13154_5238.t3 VDDH.t202 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X453 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t1 GND.t186 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X454 top_segment_2_0.rseg_2_v3_0.v37.t2 top_segment_2_0.DEC0[2].t14 a_23234_19162.t3 GND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X455 a_42609_18505.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t11 top_segment_2_0.DEC1[0].t0 GND.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X456 a_15990_6674.t1 top_segment_4_1.DEC2.t10 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t0 VDDH.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X457 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t7 a_43570_17552.t0 GND.t128 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X458 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t4 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X459 top_segment_2_0.DEC2[2].t0 top_segment_2_0.DEC2[3].t9 a_41787_17802.t1 VDDH.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X460 top_segment_1_0.rseg_1_v3_1.v37.t1 top_segment_1_0.rseg_1_v3_1.v38.t1 GND.t72 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X461 a_35435_18774.t5 a_35435_18774.t4 GND.t466 GND.t465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X462 a_42245_5784.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t3 a_42271_6380.t0 VDDH.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X463 top_segment_2_0.rseg_2_v3_0.v26.t2 top_segment_2_0.rseg_2_v3_0.v27.t2 GND.t122 sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X464 a_43570_17276.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t8 GND.t346 GND.t345 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X465 top_segment_2_0.DEC0[1].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t3 a_41787_20308.t0 VDDH.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X466 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t1 top_segment_4_1.DEC0.t10 a_14452_6674.t3 VDDH.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X467 VDD.t48 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t3 VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X468 GND.t333 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t5 a_42781_11924.t0 GND.t332 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X469 a_20750_19162.t3 top_segment_2_0.DEC1[3].t4 a_21016_17121.t5 GND.t646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X470 top_segment_2_0.rseg_2_v3_0.v13.t1 top_segment_2_0.DEC0[0].t10 a_20474_19162.t1 GND.t542 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X471 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t0 GND.t44 sky130_fd_pr__res_xhigh_po_1p41 l=2.04
X472 a_41271_20650.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t10 VDDH.t293 VDDH.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X473 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t8 a_41938_2314.t0 GND.t579 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X474 SH[3].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t2 VDDH.t273 VDDH.t272 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X475 top_segment_1_0.rseg_1_v3_1.v29.t2 top_segment_1_0.rseg_1_v3_1.v30.t2 GND.t188 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X476 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t9 VDD.t198 VDD.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X477 a_30141_6674.t4 top_segment_2_0.DEC2[3].t10 top_segment_1_0.rseg_1_v3_1.v62.t2 GND.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X478 VDD.t193 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t2 VDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X479 a_42271_8914.t1 a_42245_8754.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t1 VDDH.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X480 a_42802_3150.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t12 a_42802_3066.t1 GND.t446 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X481 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t0 VDDH.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X482 top_segment_2_0.rseg_2_v3_0.v15.t1 top_segment_2_0.DEC0[0].t11 a_20198_19162.t1 GND.t566 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X483 VDD.t50 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t0 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X484 a_21302_19162.t4 top_segment_2_0.DEC1[3].t5 a_22756_17121.t4 GND.t647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X485 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t6 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X486 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t9 VDDH.t20 VDDH.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X487 a_20198_19162.t2 top_segment_2_0.DEC1[0].t5 a_21016_17121.t4 GND.t511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X488 GND.t402 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t2 a_42781_8954.t0 GND.t401 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X489 a_15990_6674.t2 top_segment_4_1.DEC1.t11 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t0 VDDH.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X490 GND.t433 GND.t434 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X491 top_segment_2_0.rseg_2_v3_0.v8.t1 top_segment_2_0.DEC0[0].t12 a_21302_19162.t2 GND.t567 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X492 VDD.t183 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 VDD.t182 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X493 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t0 DIN6.t1 VDD.t122 VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X494 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t10 VDD.t164 VDD.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X495 top_segment_2_0.rseg_2_v3_0.v14.t0 top_segment_2_0.rseg_2_v3_0.v13.t0 GND.t21 sky130_fd_pr__res_xhigh_po_1p41 l=5.47
X496 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t2 GND.t192 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X497 top_segment_2_0.DEC1[3].t0 top_segment_2_0.DEC1[2].t5 a_41787_19568.t0 VDDH.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X498 a_14176_6674.t4 top_segment_4_1.bb3.t12 a_17547_7938.t2 VDDH.t285 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X499 a_41938_2866.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t10 a_41938_2782.t1 GND.t438 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X500 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t1 top_segment_4_1.DEC3.t8 a_12326_5238.t1 VDDH.t222 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X501 GND.t241 GND.t242 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=1.63
X502 a_13588_5238.t1 top_segment_4_1.DEC0.t11 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t2 VDDH.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X503 VDDH.t260 VDDH.t258 VDDH.t259 VDDH.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X504 a_42781_11290.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t4 GND.t627 GND.t626 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X505 top_segment_2_0.rseg_2_v3_0.v28.t0 top_segment_2_0.DEC0[1].t11 a_19370_19162.t0 GND.t437 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X506 a_41787_20992.t0 top_segment_2_0.DEC0[1].t12 a_41529_20992.t0 VDDH.t204 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X507 a_42245_9744.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t2 a_42271_10340.t1 VDDH.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X508 a_15990_6674.t0 top_segment_4_1.DEC3.t9 VDDH.t224 VDDH.t223 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X509 a_43890_2966.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t3 a_43890_2882.t0 GND.t127 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X510 VDDH.t257 VDDH.t255 VDDH.t256 VDDH.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X511 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t2 top_segment_4_1.DEC1.t12 a_14728_6674.t2 VDDH.t295 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X512 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t0 GND.t44 sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X513 a_16279_17684.t2 top_segment_3_0.bb[4].t4 a_13613_17684.t3 VDDH.t280 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X514 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t12 a_42802_3150.t0 GND.t599 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X515 a_42802_2150.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t10 GND.t108 GND.t107 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X516 top_segment_2_0.rseg_2_v3_0.v28.t1 top_segment_2_0.rseg_2_v3_0.v29.t2 GND.t122 sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X517 a_19370_19162.t2 top_segment_2_0.DEC1[0].t6 a_22756_17121.t3 GND.t512 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X518 top_segment_4_1.bb2.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t4 GND.t15 GND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X519 a_28327_6674.t1 top_segment_4_1.b3.t14 a_31905_7938.t0 GND.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X520 a_42802_3066.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t12 GND.t216 GND.t215 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X521 top_segment_2_0.rseg_2_v3_0.v40.t1 top_segment_2_0.rseg_2_v3_0.v39.t1 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X522 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t13 VDD.t203 VDD.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X523 GND.t348 GND.t349 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=4.76
X524 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t5 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t7 a_35435_18538.t0 GND.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X525 VL3.t0 top_segment_4_1.b3.t15 a_16279_17684.t1 VDDH.t237 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X526 a_42802_3434.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t4 GND.t409 GND.t408 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X527 a_42271_13310.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t14 VDDH.t88 VDDH.t87 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X528 top_segment_2_0.rseg_2_v3_0.v11.t2 top_segment_2_0.DEC0[0].t13 a_20750_19162.t1 GND.t568 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X529 a_41271_17118.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t11 VDDH.t77 VDDH.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X530 GND.t563 DIN6.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t3 GND.t562 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X531 VDD.t218 DIN2.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t1 VDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X532 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t1 DIN4.t2 GND.t207 GND.t206 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X533 a_42781_8320.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t5 GND.t223 GND.t222 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X534 VDD.t141 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t1 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X535 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t1 top_segment_4_1.DEC2.t11 a_12878_5238.t2 VDDH.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X536 GND.t600 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t14 a_42781_15884.t1 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X537 top_segment_4_1.b3.t0 top_segment_4_1.bb3.t13 GND.t537 GND.t536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X538 top_segment_4_1.bb0.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t3 GND.t294 GND.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X539 VDD.t140 DIN5.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t3 VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X540 VDD.t165 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t1 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X541 top_segment_2_0.rseg_2_v3_0.v16.t2 top_segment_2_0.rseg_2_v3_0.v17.t1 GND.t8 sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X542 a_13645_18854.t0 top_segment_3_0.bb[6].t6 top_segment_3_0.rseg_3_v3_0.v8.t0 VDDH.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X543 GND.t151 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 a_42609_18505.t0 GND.t150 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X544 a_42609_17437.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t12 top_segment_2_0.DEC2[1].t0 GND.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X545 GND.t280 GND.t281 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X546 a_41529_20992.t1 top_segment_2_0.DEC0[0].t14 a_41271_20992.t0 VDDH.t294 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X547 a_42245_11724.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t17 a_42781_12280.t0 GND.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X548 a_34304_9019.t1 top_segment_4_1.b2.t6 a_33127_7938.t0 GND.t289 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X549 top_segment_1_0.rseg_1_v3_1.v29.t1 top_segment_1_0.rseg_1_v3_1.v28.t2 GND.t188 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X550 a_19203_9019.t2 top_segment_4_1.bb2.t8 a_18493_7938.t1 VDDH.t267 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X551 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t7 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X552 GND.t419 GND.t420 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X553 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t1 top_segment_4_1.DEC0.t12 a_14176_6674.t3 VDDH.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X554 GND.t635 GND.t636 GND.t8 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X555 top_segment_2_0.rseg_2_v3_0.v24.t0 top_segment_2_0.DEC0[1].t13 a_21302_19162.t0 GND.t488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X556 GND.t435 GND.t436 GND.t40 sky130_fd_pr__res_xhigh_po_1p41 l=1.68
X557 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t7 GND.t451 GND.t450 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X558 top_segment_1_0.rseg_1_v3_1.v5.t2 top_segment_1_0.rseg_1_v3_1.v6.t2 GND.t86 sky130_fd_pr__res_xhigh_po_1p41 l=2.86
X559 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t0 top_segment_4_1.DEC2.t12 a_12602_5238.t2 VDDH.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X560 VDDH.t157 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t15 a_42271_5944.t0 VDDH.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X561 top_segment_2_0.rseg_2_v3_0.v18.t2 top_segment_2_0.rseg_2_v3_0.v17.t2 GND.t8 sky130_fd_pr__res_xhigh_po_1p41 l=5.06
X562 a_42271_13864.t0 a_42245_13704.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t0 VDDH.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X563 a_31905_7938.t2 top_segment_4_1.bb3.t14 a_25891_5238.t2 GND.t531 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X564 a_15143_17684.t0 top_segment_3_0.b[6].t6 top_segment_3_0.rseg_3_v3_0.v10.t2 VDDH.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X565 a_42781_12914.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t0 GND.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X566 VDD.t89 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t1 VDD.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X567 VDDH.t159 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t16 a_42271_8914.t0 VDDH.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X568 a_15162_6674.t3 top_segment_4_1.DEC0.t13 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t2 VDDH.t121 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X569 top_segment_4_1.b1.t0 top_segment_4_1.bb1.t4 VDDH.t39 VDDH.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X570 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t5 VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X571 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t1 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X572 top_segment_2_0.rseg_2_v3_0.v32.t0 top_segment_2_0.DEC0[1].t14 a_19922_19162.t3 GND.t489 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X573 GND.t629 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t2 GND.t628 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X574 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t2 DIN2.t1 VDD.t220 VDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X575 GND.t302 DIN8.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t1 GND.t301 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X576 GND.t130 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t2 GND.t129 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X577 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t11 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X578 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t5 VDD.t195 VDD.t194 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X579 a_32733_7938.t2 top_segment_4_1.bb3.t15 a_26719_5238.t4 GND.t532 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X580 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t10 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t3 VDDH.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X581 a_21016_17121.t2 top_segment_2_0.DEC2[3].t11 VL2.t3 GND.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X582 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t0 DIN5.t1 VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X583 a_42609_19573.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t13 top_segment_2_0.DEC1[3].t1 GND.t632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X584 GND.t102 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t3 GND.t101 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X585 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t12 VDD.t16 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X586 a_13921_18854.t2 top_segment_3_0.b[6].t7 top_segment_3_0.rseg_3_v3_0.v15.t2 VDDH.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X587 top_segment_2_0.DEC0[0].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t4 a_41787_19966.t1 VDDH.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X588 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t9 VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X589 GND.t283 DIN0.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t3 GND.t282 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X590 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t2 DIN9.t2 GND.t398 GND.t397 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X591 a_29865_6674.t4 top_segment_2_0.DEC2[3].t12 top_segment_1_0.rseg_1_v3_1.v61.t2 GND.t604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X592 a_27705_5238.t2 top_segment_4_1.bb3.t16 a_33403_7938.t2 GND.t533 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X593 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t1 GND.t44 sky130_fd_pr__res_xhigh_po_1p41 l=2.14
X594 a_42781_15250.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t6 GND.t155 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X595 top_segment_2_0.rseg_2_v3_0.v1.t1 top_segment_2_0.DEC0[0].t15 a_22682_19162.t1 GND.t569 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X596 a_42609_20997.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t0 GND.t633 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X597 a_42245_13704.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t3 a_42271_14300.t1 VDDH.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X598 top_segment_2_0.rseg_2_v3_0.v18.t0 top_segment_2_0.DEC0[1].t15 a_22130_19162.t0 GND.t490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X599 top_segment_3_0.b[6].t0 top_segment_3_0.bb[6].t7 GND.t453 GND.t452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X600 a_14165_17684.t0 top_segment_3_0.b[5].t4 a_13219_17684.t1 VDDH.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X601 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t0 GND.t149 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X602 a_30417_6674.t4 top_segment_2_0.DEC2[3].t13 top_segment_1_0.rseg_1_v3_1.v63.t2 GND.t605 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X603 top_segment_3_0.bb[6].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t4 GND.t82 GND.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X604 top_segment_2_0.rseg_2_v3_0.v27.t0 top_segment_2_0.DEC0[1].t16 a_20750_19162.t0 GND.t624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X605 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t7 a_43570_20676.t0 GND.t361 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X606 GND.t291 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 a_42609_19929.t1 GND.t290 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X607 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t1 GND.t149 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X608 VDDH.t25 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t1 VDDH.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X609 a_43570_20400.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t3 GND.t203 GND.t202 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X610 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t9 GND.t132 GND.t131 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X611 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t2 top_segment_4_1.DEC1.t13 a_14452_6674.t2 VDDH.t296 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X612 GND.t360 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t3 GND.t359 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X613 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t2 top_segment_4_1.DEC0.t14 a_13154_5238.t4 VDDH.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X614 top_segment_2_0.rseg_2_v3_0.v7.t1 top_segment_2_0.DEC0[0].t16 a_23510_19162.t1 GND.t325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X615 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t10 GND.t104 GND.t103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X616 VDD.t189 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t1 VDD.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X617 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t0 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X618 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t2 DIN0.t3 GND.t285 GND.t284 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X619 a_15438_6674.t2 top_segment_4_1.DEC1.t14 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t0 VDDH.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X620 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t1 GND.t186 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X621 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t2 GND.t186 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X622 a_13337_17684.t0 top_segment_3_0.b[5].t5 a_15419_17684.t1 VDDH.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X623 a_42781_15884.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t0 GND.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X624 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t13 GND.t448 GND.t447 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X625 a_14140_5238.t4 top_segment_4_1.DEC0.t15 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t1 VDDH.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X626 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t2 DIN3.t2 GND.t298 GND.t297 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X627 top_segment_2_0.rseg_2_v3_0.v2.t2 top_segment_2_0.DEC0[0].t17 a_22130_19162.t1 GND.t326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X628 GND.t253 GND.t254 GND.t44 sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X629 top_segment_2_0.DEC1[1].t1 top_segment_2_0.DEC1[3].t6 a_41787_18884.t1 VDDH.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X630 a_43570_19252.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t15 GND.t384 GND.t383 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X631 top_segment_3_0.bb[4].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t4 VDDH.t115 VDDH.t114 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X632 GND.t424 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t0 GND.t423 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X633 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t4 a_37219_19465.t2 GND.t429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X634 a_15438_6674.t0 top_segment_4_1.DEC3.t10 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 VDDH.t225 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X635 top_segment_2_0.rseg_2_v3_0.v4.t2 top_segment_2_0.rseg_2_v3_0.v3.t2 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=8.5
X636 a_41271_17802.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t12 VDDH.t78 VDDH.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X637 a_14867_17684.t0 top_segment_3_0.bb[6].t8 top_segment_3_0.rseg_3_v3_0.v3.t0 VDDH.t216 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X638 a_43570_20676.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t5 GND.t137 GND.t136 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X639 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t0 GND.t11 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X640 a_42245_6774.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t20 a_42781_7330.t0 GND.t334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X641 a_27981_5238.t4 top_segment_2_0.DEC2[3].t14 top_segment_1_0.rseg_1_v3_1.v55.t2 GND.t606 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X642 a_41271_20308.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t13 VDDH.t79 VDDH.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X643 a_22406_19162.t1 top_segment_2_0.DEC1[1].t6 a_22756_17121.t2 GND.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X644 a_42609_18149.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 GND.t148 GND.t147 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X645 VDDH.t254 VDDH.t252 VDDH.t253 VDDH.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X646 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t12 a_43026_2518.t1 GND.t439 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X647 a_42271_6380.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t17 VDDH.t161 VDDH.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X648 top_segment_3_0.V0.t2 top_segment_3_0.rseg_3_v3_0.v1.t2 GND.t23 sky130_fd_pr__res_xhigh_po_1p41 l=3.17
X649 VDDH.t163 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t18 a_42271_13864.t1 VDDH.t162 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X650 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t12 a_43026_2886.t1 GND.t603 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X651 a_27981_5238.t1 top_segment_2_0.DEC2[2].t8 top_segment_1_0.rseg_1_v3_1.v39.t2 GND.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X652 top_segment_2_0.rseg_2_v3_0.v14.t1 top_segment_2_0.DEC0[0].t18 a_19646_19162.t1 GND.t327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X653 a_42781_7964.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t0 GND.t335 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X654 top_segment_1_0.rseg_1_v3_1.v57.t2 top_segment_1_0.rseg_1_v3_1.v56.t2 GND.t201 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X655 a_42271_5944.t1 a_42245_5784.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t1 VDDH.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X656 VDDH.t89 top_segment_2_0.DEC2[0].t11 top_segment_4_1.DEC0.t1 VDDH.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X657 a_34304_9019.t0 top_segment_4_1.bb1.t5 a_33116_9019.t1 GND.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X658 GND.t556 GND.t557 GND.t11 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X659 a_19479_9019.t1 top_segment_4_1.b1.t4 a_18319_9019.t2 VDDH.t189 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X660 a_19045_7938.t2 top_segment_4_1.bb3.t17 a_15990_6674.t4 VDDH.t282 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X661 a_15695_17684.t2 top_segment_3_0.bb[6].t9 top_segment_3_0.V0.t0 VDDH.t217 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X662 VDD.t158 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 VDD.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X663 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t2 DIN8.t1 GND.t304 GND.t303 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X664 a_41787_19226.t0 top_segment_2_0.DEC1[1].t7 a_41529_19226.t0 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X665 GND.t179 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t3 a_42781_5984.t0 GND.t178 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X666 GND.t431 a_35435_18774.t2 a_35435_18774.t3 GND.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X667 top_segment_1_0.rseg_1_v3_1.v10.t1 top_segment_2_0.DEC2[0].t12 a_28879_6674.t3 GND.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X668 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t0 GND.t186 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X669 top_segment_2_0.rseg_2_v3_0.v28.t2 top_segment_2_0.rseg_2_v3_0.v27.t1 GND.t122 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X670 top_segment_1_0.rseg_1_v3_1.v43.t0 top_segment_1_0.rseg_1_v3_1.v42.t1 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X671 a_21854_19162.t2 top_segment_2_0.DEC1[2].t6 a_22756_17121.t0 GND.t411 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X672 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t1 GND.t11 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X673 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t1 top_segment_4_1.DEC2.t13 a_14176_6674.t1 VDDH.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X674 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t1 GND.t192 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X675 a_16555_17684.t0 top_segment_3_0.b[4].t4 a_13337_17684.t1 VDDH.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X676 a_21596_17121.t0 top_segment_2_0.DEC2[1].t15 VH2.t0 GND.t581 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X677 a_32457_7938.t2 top_segment_4_1.bb3.t18 a_26443_5238.t2 GND.t534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X678 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t8 a_43570_20952.t0 GND.t524 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X679 a_29865_6674.t3 top_segment_2_0.DEC2[0].t13 top_segment_1_0.rseg_1_v3_1.v13.t2 GND.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X680 top_segment_2_0.rseg_2_v3_0.v23.t2 top_segment_2_0.DEC0[1].t17 a_23510_19162.t3 GND.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X681 VDD.t143 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 VDD.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X682 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t15 a_41714_3346.t1 GND.t449 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X683 VDD.t18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t0 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X684 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t0 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=1.27
X685 a_41271_19568.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t14 VDDH.t80 VDDH.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X686 a_27429_5238.t2 top_segment_4_1.bb3.t19 a_33127_7938.t2 GND.t191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X687 a_15162_6674.t1 top_segment_4_1.DEC2.t14 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t1 VDDH.t132 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X688 VDD.t74 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t2 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X689 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t0 GND.t149 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X690 top_segment_2_0.rseg_2_v3_0.v45.t2 top_segment_2_0.DEC0[2].t15 a_20474_19162.t3 GND.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X691 a_43026_2518.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t14 GND.t318 GND.t317 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X692 top_segment_1_0.rseg_1_v3_1.v15.t1 top_segment_1_0.rseg_1_v3_1.v16.t2 GND.t40 sky130_fd_pr__res_xhigh_po_1p41 l=1.68
X693 top_segment_2_0.rseg_2_v3_0.v30.t2 top_segment_2_0.rseg_2_v3_0.v29.t1 GND.t122 sky130_fd_pr__res_xhigh_po_1p41 l=4.65
X694 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t11 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t2 VDDH.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X695 SH[2].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t3 GND.t367 GND.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X696 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t10 VDDH.t22 VDDH.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X697 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t13 a_41714_2150.t1 GND.t217 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X698 a_29589_6674.t4 top_segment_2_0.DEC2[3].t15 top_segment_1_0.rseg_1_v3_1.v60.t1 GND.t607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X699 a_43026_2886.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t15 GND.t320 GND.t319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X700 VDD.t68 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t4 a_41394_3894.t0 VDD.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X701 top_segment_3_0.rseg_3_v3_0.v4.t2 top_segment_3_0.rseg_3_v3_0.v3.t1 GND.t23 sky130_fd_pr__res_xhigh_po_1p41 l=3.37
X702 a_42609_19217.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t15 top_segment_2_0.DEC1[2].t0 GND.t634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X703 GND.t399 GND.t400 GND.t186 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X704 a_42271_9350.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t19 VDDH.t230 VDDH.t229 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X705 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t2 GND.t11 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X706 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t13 VDD.t208 VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X707 VDD.t160 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t0 VDD.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X708 a_42271_10340.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t20 VDDH.t232 VDDH.t231 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X709 a_41529_19226.t1 top_segment_2_0.DEC1[0].t7 a_41271_19226.t1 VDDH.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X710 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t0 VDDH.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X711 top_segment_3_0.rseg_3_v3_0.v2.t1 top_segment_3_0.rseg_3_v3_0.v1.t1 GND.t23 sky130_fd_pr__res_xhigh_po_1p41 l=3.27
X712 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t15 VDD.t162 VDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X713 a_42245_6774.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t4 a_42271_7370.t0 VDDH.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X714 a_30417_6674.t0 top_segment_2_0.DEC2[1].t16 top_segment_1_0.rseg_1_v3_1.v31.t0 GND.t351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X715 GND.t601 GND.t602 GND.t201 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X716 VDDH.t13 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t11 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t0 VDDH.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X717 a_21578_19162.t1 top_segment_2_0.DEC1[2].t7 a_21596_17121.t4 GND.t412 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X718 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t0 top_segment_4_1.DEC1.t15 a_14176_6674.t2 VDDH.t298 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X719 GND.t442 GND.t443 GND.t8 sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X720 top_segment_2_0.rseg_2_v3_0.v40.t2 top_segment_2_0.DEC0[2].t16 a_21302_19162.t3 GND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X721 a_41787_18144.t0 top_segment_2_0.DEC2[1].t17 a_41529_18144.t0 VDDH.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X722 a_17271_7938.t1 top_segment_4_1.b3.t16 a_12326_5238.t0 VDDH.t238 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X723 GND.t114 GND.t115 GND.t48 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X724 GND.t561 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t6 a_42781_12914.t1 GND.t560 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X725 top_segment_4_1.b0.t0 top_segment_4_1.bb0.t4 GND.t84 GND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X726 a_38483_21071.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t1 VDDH.t154 sky130_fd_pr__pfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=1
X727 VDDH.t304 top_segment_2_0.DEC2[3].t16 top_segment_4_1.DEC3.t1 VDDH.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X728 a_15162_6674.t2 top_segment_4_1.DEC1.t16 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t1 VDDH.t299 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X729 a_41714_3346.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t16 GND.t386 GND.t385 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X730 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t2 top_segment_4_1.DEC3.t11 a_12602_5238.t1 VDDH.t226 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X731 GND.t393 GND.t394 GND.t149 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X732 top_segment_2_0.rseg_2_v3_0.v38.t1 top_segment_2_0.rseg_2_v3_0.v37.t1 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=5.01
X733 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t4 GND.t244 GND.t243 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X734 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t12 VDD.t191 VDD.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X735 top_segment_2_0.rseg_2_v3_0.v24.t2 top_segment_2_0.rseg_2_v3_0.v23.t1 GND.t8 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X736 a_21016_17121.t1 top_segment_2_0.DEC2[2].t9 VH2.t1 GND.t312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X737 SH[4].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t4 VDDH.t1 VDDH.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X738 a_15162_6674.t0 top_segment_4_1.DEC3.t12 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t2 VDDH.t227 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X739 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t10 a_42802_2426.t0 GND.t133 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X740 VDD.t97 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 VDD.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X741 top_segment_4_1.bb0.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t4 VDDH.t68 VDDH.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X742 a_42271_9904.t1 a_42245_9744.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t1 VDDH.t209 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X743 a_28603_6674.t2 top_segment_4_1.b3.t17 a_32181_7938.t1 GND.t463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X744 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t14 VDD.t210 VDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X745 top_segment_1_0.rseg_1_v3_1.v27.t1 top_segment_1_0.rseg_1_v3_1.v28.t1 GND.t188 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X746 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t1 top_segment_4_1.DEC0.t16 a_12602_5238.t4 VDDH.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X747 a_19094_19162.t1 top_segment_2_0.DEC1[3].t7 a_21596_17121.t1 GND.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X748 a_42271_10894.t1 a_42245_10734.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t1 VDDH.t310 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X749 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t0 GND.t186 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X750 top_segment_1_0.rseg_1_v3_1.v63.t0 top_segment_1_0.rseg_1_v3_1.v62.t1 GND.t201 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X751 a_27705_5238.t4 top_segment_2_0.DEC2[3].t17 top_segment_1_0.rseg_1_v3_1.v54.t2 GND.t543 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X752 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t2 GND.t149 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X753 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t0 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X754 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t2 GND.t48 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X755 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t2 GND.t186 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X756 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t6 VDD.t146 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X757 a_27705_5238.t3 top_segment_2_0.DEC2[0].t14 top_segment_1_0.rseg_1_v3_1.v6.t1 GND.t177 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X758 a_41529_18144.t1 top_segment_2_0.DEC2[0].t15 a_41271_18144.t1 VDDH.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X759 VDD.t83 DIN8.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t3 VDD.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X760 VDD.t26 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t0 VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X761 GND.t370 GND.t371 GND.t44 sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X762 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t2 GND.t192 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X763 a_27705_5238.t1 top_segment_2_0.DEC2[2].t10 top_segment_1_0.rseg_1_v3_1.v38.t2 GND.t313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X764 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t3 DIN9.t3 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X765 top_segment_4_1.V0.t0 top_segment_3_0.rseg_3_v3_0.v15.t0 GND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=5.42
X766 top_segment_2_0.rseg_2_v3_0.v46.t0 top_segment_2_0.rseg_2_v3_0.v47.t0 GND.t181 sky130_fd_pr__res_xhigh_po_1p41 l=6.09
X767 a_42781_12280.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t4 GND.t300 GND.t299 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X768 top_segment_1_0.rseg_1_v3_1.v43.t1 top_segment_2_0.DEC2[2].t11 a_29155_6674.t2 GND.t314 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X769 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t8 VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X770 VDDH.t181 top_segment_2_0.DEC2[2].t12 top_segment_4_1.DEC2.t1 VDDH.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X771 a_42245_10734.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t3 a_42271_11330.t1 VDDH.t207 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X772 top_segment_1_0.rseg_1_v3_1.v43.t2 top_segment_1_0.rseg_1_v3_1.v44.t2 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X773 a_41271_19966.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t15 VDDH.t182 VDDH.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X774 a_27705_5238.t0 top_segment_2_0.DEC2[1].t18 top_segment_1_0.rseg_1_v3_1.v22.t0 GND.t376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X775 a_43570_17552.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t10 GND.t382 GND.t69 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X776 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t16 a_42802_2702.t0 GND.t389 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X777 top_segment_1_0.rseg_1_v3_1.v21.t2 top_segment_1_0.rseg_1_v3_1.v20.t2 GND.t49 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X778 VDDH.t208 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t1 GND.t44 sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X779 a_30141_6674.t2 top_segment_2_0.DEC2[2].t13 top_segment_1_0.rseg_1_v3_1.v46.t2 GND.t337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X780 top_segment_2_0.rseg_2_v3_0.v31.t0 top_segment_2_0.DEC0[1].t18 a_20198_19162.t0 GND.t625 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X781 a_19203_9019.t1 top_segment_4_1.b1.t5 a_18015_9019.t2 VDDH.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X782 a_42802_2426.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t15 GND.t640 GND.t639 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X783 top_segment_4_1.bb3.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t4 GND.t17 GND.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X784 top_segment_1_0.rseg_1_v3_1.v9.t0 top_segment_1_0.rseg_1_v3_1.v8.t0 GND.t40 sky130_fd_pr__res_xhigh_po_1p41 l=2.35
X785 top_segment_2_0.rseg_2_v3_0.v6.t2 top_segment_2_0.rseg_2_v3_0.v7.t2 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=7.01
X786 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t2 top_segment_4_1.DEC2.t15 a_13900_6674.t0 VDDH.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X787 GND.t585 GND.t586 GND.t201 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X788 a_13771_17684.t2 top_segment_3_0.b[6].t8 top_segment_3_0.rseg_3_v3_0.v14.t2 VDDH.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X789 top_segment_2_0.rseg_2_v3_0.v36.t2 top_segment_2_0.DEC0[2].t17 a_21854_19162.t4 GND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X790 a_29589_6674.t3 top_segment_2_0.DEC2[0].t16 top_segment_1_0.rseg_1_v3_1.v12.t2 GND.t551 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X791 a_19370_19162.t4 top_segment_2_0.DEC1[3].t8 a_20740_17121.t4 GND.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X792 top_segment_3_0.rseg_3_v3_0.v10.t0 top_segment_3_0.rseg_3_v3_0.v11.t0 GND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=4.19
X793 a_42271_14300.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t21 VDDH.t234 VDDH.t233 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X794 a_18319_9019.t0 top_segment_4_1.b0.t3 VS4.t0 VDDH.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X795 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t2 top_segment_4_1.V0.t2 GND.t11 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X796 a_27429_5238.t1 top_segment_2_0.DEC2[2].t14 top_segment_1_0.rseg_1_v3_1.v37.t2 GND.t338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X797 a_13219_17684.t2 top_segment_3_0.bb[5].t5 a_13061_17684.t2 VDDH.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X798 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t0 top_segment_4_1.DEC2.t16 a_14728_6674.t1 VDDH.t308 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X799 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t1 top_segment_2_0.DEC0[2].t18 a_41787_20992.t1 VDDH.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X800 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t12 VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X801 a_30141_6674.t3 top_segment_2_0.DEC2[0].t17 top_segment_1_0.rseg_1_v3_1.v14.t2 GND.t552 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X802 GND.t630 GND.t631 GND.t192 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X803 top_segment_1_0.rseg_1_v3_1.v59.t1 top_segment_2_0.DEC2[3].t18 a_29155_6674.t4 GND.t544 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X804 GND.t481 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 a_42609_19217.t1 GND.t480 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X805 a_42609_18149.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t16 top_segment_2_0.DEC2[3].t0 GND.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X806 top_segment_2_0.V0.t1 top_segment_2_0.rseg_2_v3_0.v1.t2 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=11.57
X807 a_19203_9019.t0 top_segment_4_1.b2.t7 a_17547_7938.t0 VDDH.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X808 a_41787_18542.t0 top_segment_2_0.DEC1[2].t8 a_41529_18542.t0 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X809 top_segment_3_0.b[4].t0 top_segment_3_0.bb[4].t5 GND.t517 GND.t516 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X810 a_34580_9019.t0 top_segment_4_1.bb1.t6 a_33420_9019.t0 GND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X811 VDD.t114 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t1 VDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X812 top_segment_2_0.rseg_2_v3_0.v30.t1 top_segment_2_0.rseg_2_v3_0.v31.t1 GND.t122 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X813 VDD.t38 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X814 VDD.t64 DIN1.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t1 VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X815 a_33724_9019.t2 top_segment_4_1.bb2.t9 a_32733_7938.t1 GND.t497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X816 a_42245_12714.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t22 a_42781_13270.t0 GND.t336 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X817 top_segment_4_1.bb1.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t4 VDDH.t206 VDDH.t205 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X818 VDD.t57 DIN4.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t2 VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X819 a_18623_9019.t1 top_segment_4_1.b2.t8 a_18099_7938.t0 VDDH.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X820 top_segment_2_0.rseg_2_v3_0.v33.t2 top_segment_2_0.DEC0[2].t19 a_22682_19162.t3 GND.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X821 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t14 a_43890_2242.t0 GND.t415 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X822 top_segment_2_0.rseg_2_v3_0.v20.t2 top_segment_2_0.rseg_2_v3_0.v19.t1 GND.t8 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X823 a_19922_19162.t1 top_segment_2_0.DEC1[0].t8 a_20740_17121.t3 GND.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X824 a_30141_6674.t0 top_segment_2_0.DEC2[1].t19 top_segment_1_0.rseg_1_v3_1.v30.t0 GND.t377 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X825 top_segment_2_0.rseg_2_v3_0.v44.t2 top_segment_2_0.DEC0[2].t20 a_19370_19162.t3 GND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X826 top_segment_1_0.rseg_1_v3_1.v23.t2 top_segment_1_0.rseg_1_v3_1.v22.t1 GND.t49 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X827 a_41271_18884.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t16 VDDH.t183 VDDH.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X828 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t4 VDD.t175 VDD.t174 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X829 top_segment_2_0.rseg_2_v3_0.v14.t2 top_segment_2_0.rseg_2_v3_0.v15.t2 GND.t21 sky130_fd_pr__res_xhigh_po_1p41 l=5.32
X830 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t16 a_41938_2866.t1 GND.t170 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X831 a_22756_17121.t1 top_segment_2_0.DEC2[0].t18 VL2.t2 GND.t553 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X832 top_segment_1_0.rseg_1_v3_1.v58.t2 top_segment_2_0.DEC2[3].t19 a_28879_6674.t4 GND.t545 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X833 top_segment_2_0.rseg_2_v3_0.v34.t0 top_segment_2_0.rseg_2_v3_0.v35.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=4.81
X834 VDDH.t15 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t12 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t0 VDDH.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X835 a_41938_2782.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t15 a_41938_2698.t1 GND.t416 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X836 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t2 GND.t186 sky130_fd_pr__res_xhigh_po_1p41 l=1.22
X837 GND.t258 GND.t259 GND.t23 sky130_fd_pr__res_xhigh_po_1p41 l=3.17
X838 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t0 GND.t11 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X839 a_42781_13904.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t1 GND.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X840 VDDH.t236 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t22 a_42271_9904.t0 VDDH.t235 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X841 a_43890_2882.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t4 GND.t157 GND.t156 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X842 top_segment_1_0.rseg_1_v3_1.v41.t1 top_segment_1_0.rseg_1_v3_1.v42.t0 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X843 top_segment_4_1.b2.t1 top_segment_4_1.bb2.t10 VDDH.t269 VDDH.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X844 VDDH.t147 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t23 a_42271_10894.t0 VDDH.t146 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X845 top_segment_1_0.rseg_1_v3_1.v13.t1 top_segment_1_0.rseg_1_v3_1.v14.t0 GND.t40 sky130_fd_pr__res_xhigh_po_1p41 l=1.84
X846 top_segment_3_0.V0.t1 top_segment_2_0.rseg_2_v3_0.v47.t1 GND.t279 sky130_fd_pr__res_xhigh_po_1p41 l=6.35
X847 a_37219_19465.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t3 GND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X848 top_segment_1_0.rseg_1_v3_1.v7.t0 top_segment_1_0.rseg_1_v3_1.v6.t0 GND.t86 sky130_fd_pr__res_xhigh_po_1p41 l=2.66
X849 top_segment_1_0.rseg_1_v3_1.v63.t1 top_segment_2_0.V0.t2 GND.t201 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X850 a_41529_18542.t1 top_segment_2_0.DEC1[1].t8 a_41271_18542.t1 VDDH.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X851 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t2 GND.t48 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X852 VDDH.t251 VDDH.t248 VDDH.t250 VDDH.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X853 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t11 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X854 top_segment_1_0.rseg_1_v3_1.v15.t0 top_segment_1_0.rseg_1_v3_1.v14.t1 GND.t40 sky130_fd_pr__res_xhigh_po_1p41 l=1.73
X855 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t2 GND.t186 sky130_fd_pr__res_xhigh_po_1p41 l=1.12
X856 a_42781_16240.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t17 GND.t390 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X857 top_segment_4_1.V0.t1 top_segment_4_1.DEC0.t17 a_12326_5238.t4 VDDH.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X858 a_42245_14694.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t3 a_42271_15290.t0 VDDH.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X859 GND.t548 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t0 GND.t547 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X860 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t0 DIN8.t3 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X861 top_segment_3_0.rseg_3_v3_0.v14.t0 top_segment_3_0.rseg_3_v3_0.v15.t1 GND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=5.12
X862 a_13219_17684.t3 top_segment_3_0.b[6].t9 top_segment_3_0.rseg_3_v3_0.v12.t0 VDDH.t178 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X863 a_41787_17460.t0 top_segment_2_0.DEC2[2].t15 a_41529_17460.t0 VDDH.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X864 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t2 top_segment_4_1.DEC3.t13 a_14728_6674.t0 VDDH.t228 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X865 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t2 GND.t4 sky130_fd_pr__res_xhigh_po_1p41 l=1.48
X866 GND.t575 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t1 GND.t574 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X867 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t5 VDD.t170 VDD.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X868 VDD.t156 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t1 VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X869 a_42609_18861.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 GND.t274 GND.t273 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X870 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t18 a_43570_19528.t0 GND.t391 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X871 VDD.t148 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t3 VDD.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X872 a_27429_5238.t3 top_segment_2_0.DEC2[0].t19 top_segment_1_0.rseg_1_v3_1.v5.t0 GND.t554 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X873 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t2 DIN6.t3 GND.t565 GND.t564 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X874 a_15714_6674.t3 top_segment_4_1.DEC3.t14 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t0 VDDH.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X875 a_13495_17684.t1 top_segment_3_0.bb[5].t6 a_13337_17684.t2 VDDH.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X876 a_42245_15684.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t24 a_42781_16240.t1 GND.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X877 a_42541_21510.t1 ROUT.t2 ROUT.t3 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X878 a_41938_2698.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t16 GND.t321 GND.t230 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X879 GND.t615 a_35435_18774.t7 a_35435_18538.t3 GND.t430 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X880 top_segment_1_0.rseg_1_v3_1.v1.t1 top_segment_1_0.rseg_1_v3_1.v2.t0 GND.t86 sky130_fd_pr__res_xhigh_po_1p41 l=4.24
X881 GND.t354 GND.t355 GND.t186 sky130_fd_pr__res_xhigh_po_1p41 l=1.02
X882 top_segment_1_0.rseg_1_v3_1.v49.t1 top_segment_2_0.DEC2[3].t20 a_26167_5238.t4 GND.t546 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X883 top_segment_2_0.rseg_2_v3_0.v22.t1 top_segment_2_0.DEC0[1].t19 a_21578_19162.t0 GND.t268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X884 a_42541_21510.t3 ROUT.t4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t0 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X885 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t17 a_43570_18700.t1 GND.t171 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X886 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t5 a_43890_2966.t1 GND.t255 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X887 GND.t340 top_segment_2_0.DEC2[2].t16 top_segment_4_1.DEC2.t0 GND.t339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X888 a_27153_5238.t4 top_segment_2_0.DEC2[3].t21 top_segment_1_0.rseg_1_v3_1.v52.t2 GND.t513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X889 a_15419_17684.t2 top_segment_3_0.b[6].t10 top_segment_3_0.rseg_3_v3_0.v9.t2 VDDH.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X890 a_22176_17121.t0 top_segment_2_0.DEC2[1].t20 VL2.t0 GND.t623 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X891 a_14140_5238.t0 top_segment_4_1.b3.t18 a_18769_7938.t1 VDDH.t239 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X892 top_segment_1_0.rseg_1_v3_1.v33.t2 top_segment_2_0.DEC2[2].t17 a_26167_5238.t1 GND.t305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X893 a_19646_19162.t2 top_segment_2_0.DEC1[0].t9 a_21596_17121.t2 GND.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X894 top_segment_3_0.b[5].t0 top_segment_3_0.bb[5].t7 VDDH.t63 VDDH.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X895 top_segment_1_0.rseg_1_v3_1.v11.t1 top_segment_1_0.rseg_1_v3_1.v10.t0 GND.t40 sky130_fd_pr__res_xhigh_po_1p41 l=2.09
X896 a_29865_6674.t2 top_segment_2_0.DEC2[2].t18 top_segment_1_0.rseg_1_v3_1.v45.t1 GND.t306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X897 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t4 VDDH.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X898 top_segment_2_0.rseg_2_v3_0.v6.t1 top_segment_2_0.DEC0[0].t19 a_21578_19162.t2 GND.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X899 VDD.t30 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X900 GND.t491 GND.t492 GND.t44 sky130_fd_pr__res_xhigh_po_1p41 l=2.55
X901 a_14416_5238.t1 top_segment_4_1.DEC3.t15 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t1 VDDH.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X902 a_41529_17460.t1 top_segment_2_0.DEC2[0].t20 a_41271_17460.t1 VDDH.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X903 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t18 GND.t577 GND.t576 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X904 top_segment_3_0.bb[5].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t4 VDDH.t31 VDDH.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X905 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t7 VDD.t167 VDD.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X906 GND.t559 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t3 GND.t558 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X907 a_27153_5238.t1 top_segment_2_0.DEC2[2].t19 top_segment_1_0.rseg_1_v3_1.v36.t2 GND.t307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X908 a_27981_5238.t3 top_segment_2_0.DEC2[0].t21 top_segment_1_0.rseg_1_v3_1.v7.t1 GND.t555 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X909 a_43570_19528.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t16 GND.t642 GND.t641 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X910 VDD.t42 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t0 VDD.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X911 VDD.t81 DIN3.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t0 VDD.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X912 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t12 VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X913 top_segment_1_0.rseg_1_v3_1.v11.t2 top_segment_2_0.DEC2[0].t22 a_29155_6674.t3 GND.t218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X914 a_13495_17684.t0 top_segment_3_0.bb[6].t10 top_segment_3_0.rseg_3_v3_0.v5.t1 VDDH.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X915 GND.t494 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t7 a_42781_9944.t1 GND.t493 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X916 GND.t71 DIN7.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t1 GND.t70 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X917 GND.t109 GND.t110 GND.t40 sky130_fd_pr__res_xhigh_po_1p41 l=2.35
X918 top_segment_1_0.rseg_1_v3_1.v39.t0 top_segment_1_0.rseg_1_v3_1.v40.t1 GND.t72 sky130_fd_pr__res_xhigh_po_1p41 l=0.86
X919 top_segment_2_0.rseg_2_v3_0.v46.t1 top_segment_2_0.rseg_2_v3_0.v45.t1 GND.t181 sky130_fd_pr__res_xhigh_po_1p41 l=5.88
X920 a_42541_21510.t2 ROUT.t5 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t1 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X921 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t2 DIN1.t3 VDD.t66 VDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X922 a_42245_7764.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t25 a_42781_8320.t0 GND.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X923 a_42609_19929.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t17 top_segment_2_0.DEC0[0].t0 GND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X924 a_20740_17121.t1 top_segment_2_0.DEC2[3].t22 VH2.t3 GND.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X925 GND.t638 DIN2.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t3 GND.t637 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X926 a_33679_7938.t1 top_segment_4_1.b3.t19 a_30417_6674.t1 GND.t464 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X927 VDD.t187 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t3 VDD.t186 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X928 a_43890_2242.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t17 GND.t644 GND.t643 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X929 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t1 GND.t48 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X930 GND.t373 DIN5.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t1 GND.t372 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X931 a_16555_17684.t3 top_segment_3_0.bb[4].t6 a_13889_17684.t2 VDDH.t281 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X932 a_42609_20285.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 GND.t94 GND.t93 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X933 a_34000_9019.t2 top_segment_4_1.bb2.t11 a_32457_7938.t1 GND.t498 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X934 VDDH.t149 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t24 a_38483_21071.t2 VDDH.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9.2
X935 a_42271_7370.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t25 VDDH.t151 VDDH.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X936 VDDH.t153 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t26 a_42271_14854.t0 VDDH.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X937 a_18899_9019.t0 top_segment_4_1.b2.t9 a_17823_7938.t0 VDDH.t276 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X938 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t6 a_41938_3162.t1 GND.t249 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X939 top_segment_1_0.rseg_1_v3_1.v27.t2 top_segment_1_0.rseg_1_v3_1.v26.t1 GND.t188 sky130_fd_pr__res_xhigh_po_1p41 l=1.17
X940 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t1 GND.t192 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X941 SH[1].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t4 VDDH.t66 VDDH.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X942 a_42781_8954.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t26 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t0 GND.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X943 top_segment_1_0.rseg_1_v3_1.v61.t0 top_segment_1_0.rseg_1_v3_1.v62.t0 GND.t201 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X944 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t1 GND.t11 sky130_fd_pr__res_xhigh_po_1p41 l=0.55
X945 a_42271_6934.t1 a_42245_6774.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t1 VDDH.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X946 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t2 a_38483_21071.t0 VDDH.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=1
X947 top_segment_1_0.rseg_1_v3_1.v13.t0 top_segment_1_0.rseg_1_v3_1.v12.t1 GND.t40 sky130_fd_pr__res_xhigh_po_1p41 l=1.89
X948 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t1 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X949 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t13 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t0 VDDH.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X950 a_33420_9019.t1 top_segment_4_1.bb0.t5 VS1.t0 GND.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X951 top_segment_1_0.rseg_1_v3_1.v57.t1 top_segment_2_0.DEC2[3].t23 a_28603_6674.t1 GND.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X952 top_segment_2_0.rseg_2_v3_0.v20.t0 top_segment_2_0.rseg_2_v3_0.v21.t0 GND.t8 sky130_fd_pr__res_xhigh_po_1p41 l=4.86
X953 a_13921_18854.t1 top_segment_3_0.bb[5].t8 a_13889_17684.t1 VDDH.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X954 a_22130_19162.t2 top_segment_2_0.DEC1[1].t9 a_21596_17121.t3 GND.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X955 VDDH.t17 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t13 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t2 VDDH.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=1
X956 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t5 a_43570_20124.t0 GND.t347 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X957 GND.t622 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t2 GND.t416 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X958 GND.t457 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t7 a_42781_6974.t1 GND.t456 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X959 GND.t487 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t2 GND.t486 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X960 GND.t343 GND.t344 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=6.65
X961 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t2 DIN7.t3 GND.t112 GND.t111 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X962 a_13921_18854.t0 top_segment_3_0.bb[6].t11 top_segment_3_0.rseg_3_v3_0.v7.t0 VDDH.t219 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X963 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t8 GND.t496 GND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X964 GND.t166 GND.t167 GND.t33 sky130_fd_pr__res_xhigh_po_1p41 l=5.42
X965 VDDH.t6 top_segment_2_0.DEC2[1].t21 top_segment_4_1.DEC1.t1 VDDH.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X966 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t19 VDD.t176 VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X967 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t17 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X968 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t0 DIN2.t3 GND.t455 GND.t454 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X969 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t8 GND.t550 GND.t549 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X970 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t5 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X971 top_segment_1_0.rseg_1_v3_1.v3.t0 top_segment_1_0.rseg_1_v3_1.v4.t0 GND.t86 sky130_fd_pr__res_xhigh_po_1p41 l=3.37
X972 a_37853_19465.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t3 GND.t256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
X973 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t16 VDD.t133 VDD.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X974 top_segment_1_0.rseg_1_v3_1.v23.t1 top_segment_1_0.rseg_1_v3_1.v24.t1 GND.t49 sky130_fd_pr__res_xhigh_po_1p41 l=1.32
X975 a_42541_21510.t0 ROUT.t0 ROUT.t1 VDDH.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=20
X976 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t2 DIN5.t3 GND.t375 GND.t374 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X977 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t1 GND.t48 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X978 a_14416_5238.t2 top_segment_4_1.DEC2.t17 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t2 VDDH.t309 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X979 a_29589_6674.t0 top_segment_2_0.DEC2[1].t22 top_segment_1_0.rseg_1_v3_1.v28.t0 GND.t473 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X980 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t13 a_41714_3622.t0 GND.t123 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X981 top_segment_2_0.rseg_2_v3_0.v12.t0 top_segment_2_0.rseg_2_v3_0.v11.t0 GND.t21 sky130_fd_pr__res_xhigh_po_1p41 l=5.73
X982 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t5 VDD.t130 VDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X983 top_segment_1_0.rseg_1_v3_1.v21.t1 top_segment_1_0.rseg_1_v3_1.v22.t2 GND.t49 sky130_fd_pr__res_xhigh_po_1p41 l=1.37
X984 GND.t12 GND.t13 GND.t11 sky130_fd_pr__res_xhigh_po_1p41 l=0.61
X985 a_13864_5238.t3 top_segment_4_1.DEC1.t17 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t1 VDDH.t300 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X986 SH[3].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t3 GND.t500 GND.t499 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X987 GND.t482 GND.t483 GND.t324 sky130_fd_pr__res_xhigh_po_1p41 l=5.22
X988 top_segment_2_0.DEC1[2].t1 top_segment_2_0.DEC1[3].t9 a_41787_19226.t1 VDDH.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X989 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t1 top_segment_4_1.DEC3.t16 a_14452_6674.t0 VDDH.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X990 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t4 GND.t428 GND.t427 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X991 top_segment_1_0.rseg_1_v3_1.v51.t0 top_segment_1_0.rseg_1_v3_1.v50.t0 GND.t3 sky130_fd_pr__res_xhigh_po_1p41 l=0.71
X992 a_37853_19465.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t27 GND.t514 GND.t513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=5.3
X993 a_43570_20952.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t9 GND.t238 GND.t237 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X994 a_41787_20650.t0 top_segment_2_0.DEC0[1].t20 a_41529_20650.t0 VDDH.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X995 a_13219_17684.t0 top_segment_3_0.bb[6].t12 top_segment_3_0.rseg_3_v3_0.v4.t1 VDDH.t220 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X996 top_segment_2_0.rseg_2_v3_0.v19.t0 top_segment_2_0.DEC0[1].t21 a_22958_19162.t0 GND.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X997 a_42271_11330.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t27 VDDH.t287 VDDH.t286 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
X998 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t4 GND.t231 GND.t230 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X999 top_segment_1_0.rseg_1_v3_1.v37.t0 top_segment_1_0.rseg_1_v3_1.v36.t0 GND.t72 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X1000 GND.t444 GND.t445 GND.t45 sky130_fd_pr__res_xhigh_po_1p41 l=11.57
X1001 a_42245_7764.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t4 a_42271_8360.t1 VDDH.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.8
X1002 top_segment_1_0.rseg_1_v3_1.v41.t0 top_segment_1_0.rseg_1_v3_1.v40.t0 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=0.91
X1003 top_segment_2_0.rseg_2_v3_0.v44.t1 top_segment_2_0.rseg_2_v3_0.v45.t0 GND.t181 sky130_fd_pr__res_xhigh_po_1p41 l=5.73
X1004 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t2 GND.t48 sky130_fd_pr__res_xhigh_po_1p41 l=0.81
X1005 a_42781_6340.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t2 GND.t388 GND.t387 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1006 GND.t220 top_segment_2_0.DEC2[0].t23 a_25891_5238.t3 GND.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1007 top_segment_2_0.rseg_2_v3_0.v32.t2 top_segment_2_0.rseg_2_v3_0.v31.t2 GND.t122 sky130_fd_pr__res_xhigh_po_1p41 l=4.71
X1008 GND.t106 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t12 a_42781_13904.t1 GND.t105 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1009 top_segment_4_1.b1.t1 top_segment_4_1.bb1.t7 GND.t573 GND.t572 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
X1010 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t1 top_segment_4_1.DEC3.t17 a_14176_6674.t0 VDDH.t145 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1011 top_segment_1_0.rseg_1_v3_1.v41.t2 top_segment_2_0.DEC2[2].t20 a_28603_6674.t3 GND.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1012 top_segment_2_0.rseg_2_v3_0.v3.t1 top_segment_2_0.DEC0[0].t20 a_22958_19162.t1 GND.t329 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1013 a_41271_20992.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t17 VDDH.t185 VDDH.t184 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.2436 ps=2.26 w=0.84 l=1
X1014 GND.t322 GND.t323 GND.t188 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X1015 a_27153_5238.t0 top_segment_2_0.DEC2[1].t23 top_segment_1_0.rseg_1_v3_1.v20.t0 GND.t474 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1016 top_segment_2_0.rseg_2_v3_0.v34.t2 top_segment_2_0.DEC0[2].t21 a_22130_19162.t3 GND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1017 top_segment_1_0.rseg_1_v3_1.v3.t2 top_segment_2_0.DEC2[0].t24 a_26719_5238.t2 GND.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1018 a_13889_17684.t0 top_segment_3_0.b[5].t6 a_14867_17684.t1 VDDH.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1019 top_segment_1_0.rseg_1_v3_1.v51.t2 top_segment_2_0.DEC2[3].t24 a_26719_5238.t1 GND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1020 a_29589_6674.t2 top_segment_2_0.DEC2[2].t21 top_segment_1_0.rseg_1_v3_1.v44.t0 GND.t309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1021 a_42245_9744.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t28 a_42781_10300.t0 GND.t515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1022 a_35957_18086.t3 a_35957_18086.t2 GND.t121 GND.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1856 pd=1.86 as=0.1856 ps=1.86 w=0.64 l=12
X1023 top_segment_1_0.rseg_1_v3_1.v61.t1 top_segment_1_0.rseg_1_v3_1.v60.t0 GND.t201 sky130_fd_pr__res_xhigh_po_1p41 l=0.66
X1024 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t9 GND.t526 GND.t525 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1025 VDD.t134 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t0 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1026 a_27981_5238.t0 top_segment_2_0.DEC2[1].t24 top_segment_1_0.rseg_1_v3_1.v23.t0 GND.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1027 a_42609_20641.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t18 top_segment_2_0.DEC0[2].t0 GND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1028 VH3.t1 top_segment_4_1.bb3.t20 a_16831_17684.t1 VDDH.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1029 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t8 a_43570_17828.t0 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1030 VDD.t108 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t4 a_41394_2698.t1 VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1031 top_segment_2_0.rseg_2_v3_0.v22.t2 top_segment_2_0.rseg_2_v3_0.v21.t2 GND.t8 sky130_fd_pr__res_xhigh_po_1p41 l=4.81
X1032 top_segment_2_0.rseg_2_v3_0.v36.t0 top_segment_2_0.rseg_2_v3_0.v37.t0 GND.t0 sky130_fd_pr__res_xhigh_po_1p41 l=4.91
X1033 VDDH.t247 VDDH.t245 VDDH.t246 VDDH.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1034 a_21302_19162.t1 top_segment_2_0.DEC1[2].t9 a_20740_17121.t0 GND.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1035 top_segment_1_0.rseg_1_v3_1.v31.t1 top_segment_1_0.rseg_1_v3_1.v30.t1 GND.t188 sky130_fd_pr__res_xhigh_po_1p41 l=1.07
X1036 a_30417_6674.t2 top_segment_2_0.DEC2[2].t22 top_segment_1_0.rseg_1_v3_1.v47.t1 GND.t521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1037 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t0 GND.t192 sky130_fd_pr__res_xhigh_po_1p41 l=0.96
X1038 VDDH.t244 VDDH.t241 VDDH.t243 VDDH.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.522 pd=4.18 as=0 ps=0 w=1.8 l=1
X1039 a_41529_20650.t1 top_segment_2_0.DEC0[0].t21 a_41271_20650.t0 VDDH.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.13 as=0.1218 ps=1.13 w=0.84 l=1
X1040 top_segment_1_0.rseg_1_v3_1.v35.t2 top_segment_2_0.DEC2[2].t23 a_26719_5238.t3 GND.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1041 top_segment_2_0.rseg_2_v3_0.v16.t0 top_segment_2_0.rseg_2_v3_0.v15.t0 GND.t21 sky130_fd_pr__res_xhigh_po_1p41 l=5.17
X1042 top_segment_2_0.DEC2[3].t1 top_segment_2_0.DEC2[2].t24 a_41787_18144.t1 VDDH.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2436 pd=2.26 as=0.1218 ps=1.13 w=0.84 l=1
X1043 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t0 GND.t53 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X1044 a_42271_11884.t1 a_42245_11724.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t1 VDDH.t305 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.8
X1045 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t20 VDD.t178 VDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1046 a_14728_6674.t4 top_segment_4_1.bb3.t21 a_18099_7938.t2 VDDH.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.5
X1047 GND.t57 GND.t58 GND.t56 sky130_fd_pr__res_xhigh_po_1p41 l=0.76
X1048 VDDH.t289 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t28 a_42271_6934.t0 VDDH.t288 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.8
R0 GND.n126 GND.n123 93338.2
R1 GND.n1080 GND.n124 75097.7
R2 GND.n418 GND.n162 74752.4
R3 GND.n1370 GND.n13 52236.1
R4 GND.n1136 GND.n124 49116.3
R5 GND.n1079 GND.n161 40814.8
R6 GND.n983 GND.n980 39303.2
R7 GND.n1135 GND.n126 35921.1
R8 GND.n1113 GND.n146 32324.4
R9 GND.n1112 GND.n147 32324.4
R10 GND.n147 GND.n146 32321.1
R11 GND.n1113 GND.n1112 32321.1
R12 GND.n1077 GND.n162 31697.7
R13 GND.n1080 GND.n159 30691.4
R14 GND.n947 GND.n98 28676.6
R15 GND.n947 GND.n99 28676.6
R16 GND.n1168 GND.n98 28673.3
R17 GND.n1168 GND.n99 28673.3
R18 GND.n1165 GND.n100 27409.3
R19 GND.n1165 GND.n101 27409.3
R20 GND.n1141 GND.n100 27406
R21 GND.n1141 GND.n101 27406
R22 GND.n1270 GND.t199 19674.4
R23 GND.n975 GND.n971 19032.4
R24 GND.t499 GND.t116 15956
R25 GND.t366 GND.t499 15956
R26 GND.t199 GND.t366 15956
R27 GND.t243 GND.t172 15812.5
R28 GND.n363 GND.t452 15691
R29 GND.n900 GND.n60 15303.1
R30 GND.n1270 GND.t243 15099.2
R31 GND.n970 GND.n161 14517.6
R32 GND.n1079 GND.n160 14097.4
R33 GND.t116 GND.t293 13619
R34 GND.n382 GND.n367 13432.1
R35 GND.n382 GND.n368 13432.1
R36 GND.n379 GND.n367 13432.1
R37 GND.n379 GND.n368 13432.1
R38 GND.n1236 GND.n1201 12669.3
R39 GND.t81 GND.t275 11314.3
R40 GND.t38 GND.t516 11314.3
R41 GND.t458 GND.t536 11314.3
R42 GND.t16 GND.t227 11314.3
R43 GND.t14 GND.t572 11314.3
R44 GND.n983 GND.n981 11217.1
R45 GND.n1139 GND.n121 10583.4
R46 GND.n1078 GND.n1077 10105.7
R47 GND.n1080 GND.n1079 10065.1
R48 GND.n1128 GND.n132 10050.6
R49 GND.n1126 GND.n132 10050.6
R50 GND.n1370 GND.n1369 9941.15
R51 GND.n975 GND.n122 9936.26
R52 GND.t230 GND.t579 9900
R53 GND.n980 GND.n979 9777.78
R54 GND.n1128 GND.n133 9474.26
R55 GND.n1126 GND.n134 9474.26
R56 GND.n978 GND.n977 9451.85
R57 GND.n976 GND.n121 9253.97
R58 GND.n979 GND.n978 9201.59
R59 GND.n977 GND.n976 8875.66
R60 GND.n1077 GND.n167 8850.66
R61 GND.n1089 GND.n158 8548.9
R62 GND.n1088 GND.n158 8548.9
R63 GND.n1119 GND.n140 8548.9
R64 GND.n1120 GND.n140 8548.9
R65 GND.n1185 GND.n1184 8242.76
R66 GND.n1270 GND.n28 8095.54
R67 GND.n1089 GND.n151 7972.6
R68 GND.n1110 GND.n151 7972.6
R69 GND.n1110 GND.n141 7972.6
R70 GND.n1119 GND.n141 7972.6
R71 GND.n1088 GND.n1083 7972.6
R72 GND.n1083 GND.n150 7972.6
R73 GND.n150 GND.n139 7972.6
R74 GND.n1120 GND.n139 7972.6
R75 GND.t172 GND.t249 7871.88
R76 GND.n1371 GND.t612 7700
R77 GND.n1073 GND.n169 7416.07
R78 GND.n1073 GND.n170 7416.07
R79 GND.n169 GND.n168 7416.07
R80 GND.n170 GND.n168 7416.07
R81 GND.n1248 GND.n55 7376.47
R82 GND.n1224 GND.n1222 7376.47
R83 GND.n1269 GND.t595 7333.33
R84 GND.n238 GND.n237 7323.68
R85 GND.n1135 GND.n125 7195.46
R86 GND.n165 GND.n164 6513.16
R87 GND.n380 GND.n123 6249.61
R88 GND.n1236 GND.n1235 6156.3
R89 GND.t432 GND.n363 6141.67
R90 GND.n1250 GND.n44 6036.13
R91 GND.n525 GND.n524 5949.49
R92 GND.n1140 GND.n1139 5698.84
R93 GND.t7 GND.t633 5438.89
R94 GND.t202 GND.t7 5438.89
R95 GND.t202 GND.t6 5438.89
R96 GND.t632 GND.t6 5438.89
R97 GND.t632 GND.t634 5438.89
R98 GND.t68 GND.t270 5438.89
R99 GND.t5 GND.t68 5438.89
R100 GND.t5 GND.t67 5438.89
R101 GND.t67 GND.t69 5438.89
R102 GND.t69 GND.t432 5438.89
R103 GND.n971 GND.n970 5191.76
R104 GND.n525 GND.n162 5155.69
R105 GND.n1040 GND.n194 5016.93
R106 GND.n973 GND.n121 5009.74
R107 GND.n983 GND.n79 4999.47
R108 GND.n935 GND.n211 4924.62
R109 GND.n1020 GND.n211 4924.62
R110 GND.n976 GND.n975 4726.5
R111 GND.n885 GND.n884 4714.29
R112 GND.n866 GND.n743 4714.29
R113 GND.n857 GND.n856 4714.29
R114 GND.n838 GND.n775 4714.29
R115 GND.n829 GND.n828 4714.29
R116 GND.t452 GND.t81 4641.76
R117 GND.t275 GND.t38 4641.76
R118 GND.t516 GND.t458 4641.76
R119 GND.t536 GND.t16 4641.76
R120 GND.t227 GND.t14 4641.76
R121 GND.t572 GND.t595 4641.76
R122 GND.t293 GND.t83 4641.76
R123 GND.n1133 GND.n127 4597.17
R124 GND.n1133 GND.n128 4597.17
R125 GND.n1138 GND.n122 4537.46
R126 GND.n485 GND.n420 4533.07
R127 GND.n485 GND.n421 4533.07
R128 GND.n1053 GND.n177 4458.86
R129 GND.n184 GND.n177 4458.86
R130 GND.n184 GND.n176 4458.86
R131 GND.n1053 GND.n176 4458.86
R132 GND.n1000 GND.n220 4458.86
R133 GND.n1000 GND.n221 4458.86
R134 GND.n904 GND.n221 4458.86
R135 GND.n904 GND.n220 4458.86
R136 GND.n1201 GND.n61 4458.86
R137 GND.n907 GND.n61 4458.86
R138 GND.n907 GND.n62 4458.86
R139 GND.n1201 GND.n62 4458.86
R140 GND.n1183 GND.n80 4458.86
R141 GND.n88 GND.n80 4458.86
R142 GND.n88 GND.n81 4458.86
R143 GND.n1183 GND.n81 4458.86
R144 GND.n1187 GND.n76 4458.86
R145 GND.n1187 GND.n77 4458.86
R146 GND.n78 GND.n77 4458.86
R147 GND.n78 GND.n76 4458.86
R148 GND.n1067 GND.n1061 4458.86
R149 GND.n1065 GND.n1061 4458.86
R150 GND.n1065 GND.n1060 4458.86
R151 GND.n1067 GND.n1060 4458.86
R152 GND.n1175 GND.n94 4458.86
R153 GND.n1173 GND.n94 4458.86
R154 GND.n1173 GND.n93 4458.86
R155 GND.n1175 GND.n93 4458.86
R156 GND.n986 GND.n236 4458.86
R157 GND.n968 GND.n236 4458.86
R158 GND.n968 GND.n235 4458.86
R159 GND.n986 GND.n235 4458.86
R160 GND.n993 GND.n228 4458.86
R161 GND.n995 GND.n228 4458.86
R162 GND.n995 GND.n227 4458.86
R163 GND.n993 GND.n227 4458.86
R164 GND.n1193 GND.n69 4458.86
R165 GND.n1193 GND.n70 4458.86
R166 GND.n1195 GND.n69 4458.86
R167 GND.n1195 GND.n70 4458.86
R168 GND.n977 GND.n974 4451.25
R169 GND.n978 GND.n971 4206.29
R170 GND.n133 GND.n128 4020.88
R171 GND.n134 GND.n127 4020.88
R172 GND.n933 GND.n193 3998.27
R173 GND.t83 GND.n1269 3980.95
R174 GND.n1043 GND.n193 3956.88
R175 GND.n1007 GND.n1006 3883.67
R176 GND.n1006 GND.n1004 3842.28
R177 GND.n1079 GND.n1078 3789.17
R178 GND.n979 GND.n969 3752.03
R179 GND.n923 GND.n909 3641.73
R180 GND.n1136 GND.n122 3460.47
R181 GND.n980 GND.n161 3386.33
R182 GND.t579 GND.t78 3300
R183 GND.n1269 GND.n36 3253.78
R184 GND.n517 GND.n308 3250.5
R185 GND.n709 GND.n308 3250.5
R186 GND.n709 GND.n309 3250.5
R187 GND.n705 GND.n309 3250.5
R188 GND.n705 GND.n313 3250.5
R189 GND.n701 GND.n313 3250.5
R190 GND.n701 GND.n325 3250.5
R191 GND.n696 GND.n325 3250.5
R192 GND.n696 GND.n633 3250.5
R193 GND.t634 GND.n486 3193.06
R194 GND.n715 GND.n303 3151.5
R195 GND.n310 GND.n303 3151.5
R196 GND.n311 GND.n310 3151.5
R197 GND.n312 GND.n311 3151.5
R198 GND.n328 GND.n312 3151.5
R199 GND.n329 GND.n328 3151.5
R200 GND.n631 GND.n329 3151.5
R201 GND.n632 GND.n631 3151.5
R202 GND.n638 GND.n632 3151.5
R203 GND.n1004 GND.n203 3036.9
R204 GND.t78 GND.t407 2887.5
R205 GND.t407 GND.t612 2887.5
R206 GND.n916 GND.n202 2801.33
R207 GND.n1137 GND.n123 2780.4
R208 GND.n526 GND.n525 2710.35
R209 GND.n1012 GND.n210 2463.9
R210 GND.n1050 GND.n185 2381.13
R211 GND.n1373 GND.n1372 2374.87
R212 GND.n1040 GND.n195 2266.53
R213 GND.t226 GND.t52 2200
R214 GND.t51 GND.t403 2200
R215 GND.t404 GND.t85 2200
R216 GND.t85 GND.t66 2200
R217 GND.n1136 GND.n1135 2119.27
R218 GND.n1050 GND.n186 2101
R219 GND.n1023 GND.n209 2040.52
R220 GND.t52 GND.t51 1997.37
R221 GND.t403 GND.t404 1997.37
R222 GND.t533 GND.t535 1997.37
R223 GND.t191 GND.t533 1997.37
R224 GND.t225 GND.t191 1997.37
R225 GND.t532 GND.t534 1997.37
R226 GND.t534 GND.t224 1997.37
R227 GND.t224 GND.t531 1997.37
R228 GND.t338 GND.t313 1997.37
R229 GND.t307 GND.t338 1997.37
R230 GND.t97 GND.t522 1997.37
R231 GND.t305 GND.t97 1997.37
R232 GND.t99 GND.t305 1997.37
R233 GND.t376 GND.t180 1997.37
R234 GND.t100 GND.t376 1997.37
R235 GND.t474 GND.t100 1997.37
R236 GND.t46 GND.t350 1997.37
R237 GND.t350 GND.t475 1997.37
R238 GND.t475 GND.t379 1997.37
R239 GND.t555 GND.t177 1997.37
R240 GND.t177 GND.t554 1997.37
R241 GND.t554 GND.t77 1997.37
R242 GND.t221 GND.t73 1997.37
R243 GND.t73 GND.t76 1997.37
R244 GND.t76 GND.t219 1997.37
R245 GND.t351 GND.t377 1997.37
R246 GND.t377 GND.t571 1997.37
R247 GND.t571 GND.t473 1997.37
R248 GND.t47 GND.t570 1997.37
R249 GND.t570 GND.t476 1997.37
R250 GND.t476 GND.t378 1997.37
R251 GND.t552 GND.t174 1997.37
R252 GND.t176 GND.t552 1997.37
R253 GND.t551 GND.t176 1997.37
R254 GND.t175 GND.t218 1997.37
R255 GND.t352 GND.t175 1997.37
R256 GND.t74 GND.t352 1997.37
R257 GND.n1043 GND.n186 1951.38
R258 GND.n984 GND.n983 1773.03
R259 GND.t219 GND.n94 1687.7
R260 GND.n88 GND.t74 1687.7
R261 GND.n1007 GND.n209 1664.88
R262 GND.t423 GND.n28 1608.12
R263 GND.n1138 GND.n1137 1581.82
R264 GND.n1323 GND.t159 1576.25
R265 GND.t40 GND.t86 1548.86
R266 GND.t66 GND.n159 1541.45
R267 GND.t535 GND.n167 1541.45
R268 GND.t531 GND.n160 1541.45
R269 GND.n237 GND.t99 1541.45
R270 GND.t180 GND.n238 1541.45
R271 GND.t379 GND.n984 1541.45
R272 GND.n981 GND.t555 1541.45
R273 GND.t310 GND.n165 1541.45
R274 GND.n164 GND.t351 1541.45
R275 GND.t378 GND.n1185 1541.45
R276 GND.n210 GND.n195 1464.33
R277 GND.n1269 GND.n1268 1460.5
R278 GND.n933 GND.n185 1438.87
R279 GND.t4 GND.t44 1346.78
R280 GND.t174 GND.n79 1346.05
R281 GND.n1372 GND.n1371 1339.85
R282 GND.t229 GND.n1074 1302.63
R283 GND.t49 GND.t188 1261.42
R284 GND.n34 GND.n21 1255.62
R285 GND.n970 GND.n124 1240.24
R286 GND.n1237 GND.n1236 1220.17
R287 GND.n893 GND.n892 1219.11
R288 GND.n35 GND.n24 1198.25
R289 GND.n1337 GND.n25 1198.25
R290 GND.n30 GND.n17 1198.25
R291 GND.n1324 GND.n1323 1198.25
R292 GND.n1322 GND.n1321 1198.25
R293 GND.n1311 GND.n1310 1198.25
R294 GND.n1309 GND.n1308 1198.25
R295 GND.n668 GND.n654 1198.25
R296 GND.n11 GND.n10 1198.25
R297 GND.n529 GND.n526 1198.25
R298 GND.n540 GND.n359 1198.25
R299 GND.n551 GND.n355 1198.25
R300 GND.n562 GND.n351 1198.25
R301 GND.n573 GND.n347 1198.25
R302 GND.n584 GND.n343 1198.25
R303 GND.n595 GND.n339 1198.25
R304 GND.n606 GND.n335 1198.25
R305 GND.n629 GND.n628 1198.25
R306 GND.n630 GND.n2 1198.25
R307 GND.n1374 GND.n1373 1198.25
R308 GND.n1297 GND.n1294 1198.01
R309 GND.t186 GND.t4 1185.54
R310 GND.n418 GND 1178.42
R311 GND GND.n487 1177.5
R312 GND.n416 GND 1177.5
R313 GND GND.n430 1177.5
R314 GND.n429 GND 1177.5
R315 GND.n515 GND 1177.5
R316 GND.n1129 GND.n131 1153.51
R317 GND.n1137 GND.n1136 1146.44
R318 GND.n983 GND.t49 1142.5
R319 GND.t192 GND.n969 1134.47
R320 GND.n974 GND.t53 1108.21
R321 GND GND.t479 1104.21
R322 GND.t187 GND.t149 1102.37
R323 GND.n973 GND.t11 1095.81
R324 GND.n1130 GND.n1129 1083.11
R325 GND.n1125 GND.n135 1083.11
R326 GND.n523 GND.t154 1034.5
R327 GND.n1078 GND.n79 1020.1
R328 GND.n982 GND.t72 1011.91
R329 GND.n1066 GND.t225 998.684
R330 GND.n1066 GND.t532 998.684
R331 GND.n994 GND.t307 998.684
R332 GND.n994 GND.t522 998.684
R333 GND.n985 GND.t474 998.684
R334 GND.n985 GND.t46 998.684
R335 GND.n1174 GND.t77 998.684
R336 GND.n1174 GND.t221 998.684
R337 GND.n1186 GND.t473 998.684
R338 GND.n1186 GND.t47 998.684
R339 GND.n87 GND.t551 998.684
R340 GND.t218 GND.n87 998.684
R341 GND.n1057 GND.n1056 982.966
R342 GND.n1087 GND.n1084 981.836
R343 GND.n1167 GND.t86 938.22
R344 GND.t506 GND.t484 938.072
R345 GND.t154 GND.n516 935.114
R346 GND.n1087 GND.n1086 911.436
R347 GND.n1086 GND.n1085 911.436
R348 GND.n1085 GND.n136 911.436
R349 GND.n1012 GND.n209 904.067
R350 GND.n1023 GND.n203 900.884
R351 GND.t78 GND.t217 893.402
R352 GND.t407 GND.t529 893.402
R353 GND.n894 GND.n893 890.795
R354 GND.n892 GND.n722 887.395
R355 GND.n886 GND.n722 887.395
R356 GND.n886 GND.n885 887.395
R357 GND.n884 GND.n732 887.395
R358 GND.n878 GND.n732 887.395
R359 GND.n878 GND.n877 887.395
R360 GND.n877 GND.n876 887.395
R361 GND.n876 GND.n743 887.395
R362 GND.n866 GND.n865 887.395
R363 GND.n865 GND.n864 887.395
R364 GND.n864 GND.n754 887.395
R365 GND.n858 GND.n754 887.395
R366 GND.n858 GND.n857 887.395
R367 GND.n856 GND.n764 887.395
R368 GND.n850 GND.n764 887.395
R369 GND.n850 GND.n849 887.395
R370 GND.n849 GND.n848 887.395
R371 GND.n848 GND.n775 887.395
R372 GND.n838 GND.n837 887.395
R373 GND.n837 GND.n836 887.395
R374 GND.n836 GND.n786 887.395
R375 GND.n830 GND.n786 887.395
R376 GND.n830 GND.n829 887.395
R377 GND.n828 GND.n796 887.395
R378 GND.n822 GND.n796 887.395
R379 GND.n822 GND.n821 887.395
R380 GND.n821 GND.n820 887.395
R381 GND.n820 GND.n36 887.395
R382 GND.n1268 GND.n37 887.395
R383 GND.n1262 GND.n37 887.395
R384 GND.n1262 GND.n1261 887.395
R385 GND.n1261 GND.n1260 887.395
R386 GND.n1260 GND.n44 887.395
R387 GND.n1250 GND.n1249 887.395
R388 GND.n1249 GND.n1248 887.395
R389 GND.n1238 GND.n55 887.395
R390 GND.n1238 GND.n1237 887.395
R391 GND.n1235 GND.n1202 887.395
R392 GND.n1222 GND.n1202 887.395
R393 GND.n1224 GND.n1223 887.395
R394 GND.n1223 GND.n13 887.395
R395 GND.t172 GND 859.899
R396 GND.n1072 GND.n1071 852.33
R397 GND.n1072 GND.n171 852.33
R398 GND GND.n30 848.731
R399 GND.t159 GND 842.913
R400 GND.n923 GND.n916 840.4
R401 GND GND.n35 837.563
R402 GND.t33 GND.n380 835.664
R403 GND.n487 GND.n416 827.04
R404 GND.n430 GND.n429 827.04
R405 GND.n1369 GND 826.396
R406 GND.n1077 GND.t229 817.764
R407 GND.n381 GND.t23 790.207
R408 GND.t48 GND.n972 786.471
R409 GND.n174 GND.n172 781.929
R410 GND.n1070 GND.n172 781.929
R411 GND GND.t184 781.726
R412 GND.t385 GND 781.726
R413 GND.t599 GND.t292 775.48
R414 GND.n276 GND.n259 769.572
R415 GND.n285 GND.n261 769.572
R416 GND.n294 GND.n263 769.572
R417 GND.n267 GND.n264 769.572
R418 GND.n516 GND.n515 765.375
R419 GND.n1166 GND.t44 758.747
R420 GND.n1125 GND.n1124 739.765
R421 GND.t427 GND 714.721
R422 GND.t230 GND 714.721
R423 GND GND.t612 714.721
R424 GND.n1323 GND.n1271 708.047
R425 GND.t91 GND.t50 708.047
R426 GND.t317 GND.t439 708.047
R427 GND.t213 GND.t578 708.047
R428 GND.n1372 GND.n12 708.047
R429 GND.t438 GND.t416 708.047
R430 GND.t416 GND.t230 708.047
R431 GND.t23 GND.n369 701.784
R432 GND.n363 GND.t246 700.206
R433 GND.n1074 GND.t226 694.737
R434 GND.t449 GND 681.218
R435 GND.n143 GND.n138 675.013
R436 GND.n966 GND.n95 669.365
R437 GND.n381 GND.t33 656.327
R438 GND.n33 GND.n32 649.043
R439 GND.n1178 GND.n90 646.4
R440 GND.n524 GND.n523 634.702
R441 GND.n1140 GND.t11 623.778
R442 GND GND.n12 623.755
R443 GND.t579 GND 603.047
R444 GND.n1086 GND.n135 601.977
R445 GND.n1124 GND.n136 601.977
R446 GND.n1123 GND.n1122 601.977
R447 GND.n1369 GND.n1368 599.125
R448 GND.n1293 GND.n12 599.125
R449 GND.n1328 GND.n28 599.125
R450 GND.n1039 GND.n196 592.888
R451 GND.n1270 GND.t592 590.955
R452 GND.t262 GND.n33 590.039
R453 GND.t319 GND 590.038
R454 GND GND.t477 590.038
R455 GND GND.t639 590.038
R456 GND.n293 GND.n292 585
R457 GND.n291 GND.n262 585
R458 GND.n945 GND.n262 585
R459 GND.n284 GND.n283 585
R460 GND.n282 GND.n260 585
R461 GND.n945 GND.n260 585
R462 GND.n275 GND.n274 585
R463 GND.n273 GND.n258 585
R464 GND.n945 GND.n258 585
R465 GND.n944 GND.n943 585
R466 GND.n945 GND.n944 585
R467 GND.n266 GND.n265 585
R468 GND.n1220 GND.n1219 585
R469 GND.n1220 GND.n13 585
R470 GND.n1221 GND.n1214 585
R471 GND.n1223 GND.n1221 585
R472 GND.n1226 GND.n1225 585
R473 GND.n1225 GND.n1224 585
R474 GND.n1231 GND.n1211 585
R475 GND.n1222 GND.n1211 585
R476 GND.n1232 GND.n1203 585
R477 GND.n1203 GND.n1202 585
R478 GND.n1234 GND.n1233 585
R479 GND.n1235 GND.n1234 585
R480 GND.n1204 GND.n59 585
R481 GND.n1237 GND.n59 585
R482 GND.n1239 GND.n58 585
R483 GND.n1239 GND.n1238 585
R484 GND.n1241 GND.n1240 585
R485 GND.n1240 GND.n55 585
R486 GND.n1247 GND.n1246 585
R487 GND.n1248 GND.n1247 585
R488 GND.n54 GND.n53 585
R489 GND.n1249 GND.n54 585
R490 GND.n1252 GND.n1251 585
R491 GND.n1251 GND.n1250 585
R492 GND.n1257 GND.n45 585
R493 GND.n45 GND.n44 585
R494 GND.n1259 GND.n1258 585
R495 GND.n1260 GND.n1259 585
R496 GND.n43 GND.n42 585
R497 GND.n1261 GND.n43 585
R498 GND.n1264 GND.n1263 585
R499 GND.n1263 GND.n1262 585
R500 GND.n1265 GND.n38 585
R501 GND.n38 GND.n37 585
R502 GND.n1267 GND.n1266 585
R503 GND.n1268 GND.n1267 585
R504 GND.n817 GND.n807 585
R505 GND.n807 GND.n36 585
R506 GND.n819 GND.n818 585
R507 GND.n820 GND.n819 585
R508 GND.n806 GND.n805 585
R509 GND.n821 GND.n806 585
R510 GND.n824 GND.n823 585
R511 GND.n823 GND.n822 585
R512 GND.n825 GND.n797 585
R513 GND.n797 GND.n796 585
R514 GND.n827 GND.n826 585
R515 GND.n828 GND.n827 585
R516 GND.n795 GND.n794 585
R517 GND.n829 GND.n795 585
R518 GND.n832 GND.n831 585
R519 GND.n831 GND.n830 585
R520 GND.n833 GND.n787 585
R521 GND.n787 GND.n786 585
R522 GND.n835 GND.n834 585
R523 GND.n836 GND.n835 585
R524 GND.n785 GND.n784 585
R525 GND.n837 GND.n785 585
R526 GND.n840 GND.n839 585
R527 GND.n839 GND.n838 585
R528 GND.n845 GND.n776 585
R529 GND.n776 GND.n775 585
R530 GND.n847 GND.n846 585
R531 GND.n848 GND.n847 585
R532 GND.n774 GND.n773 585
R533 GND.n849 GND.n774 585
R534 GND.n852 GND.n851 585
R535 GND.n851 GND.n850 585
R536 GND.n853 GND.n765 585
R537 GND.n765 GND.n764 585
R538 GND.n855 GND.n854 585
R539 GND.n856 GND.n855 585
R540 GND.n763 GND.n762 585
R541 GND.n857 GND.n763 585
R542 GND.n860 GND.n859 585
R543 GND.n859 GND.n858 585
R544 GND.n861 GND.n755 585
R545 GND.n755 GND.n754 585
R546 GND.n863 GND.n862 585
R547 GND.n864 GND.n863 585
R548 GND.n753 GND.n752 585
R549 GND.n865 GND.n753 585
R550 GND.n868 GND.n867 585
R551 GND.n867 GND.n866 585
R552 GND.n873 GND.n744 585
R553 GND.n744 GND.n743 585
R554 GND.n875 GND.n874 585
R555 GND.n876 GND.n875 585
R556 GND.n742 GND.n741 585
R557 GND.n877 GND.n742 585
R558 GND.n880 GND.n879 585
R559 GND.n879 GND.n878 585
R560 GND.n881 GND.n733 585
R561 GND.n733 GND.n732 585
R562 GND.n883 GND.n882 585
R563 GND.n884 GND.n883 585
R564 GND.n731 GND.n730 585
R565 GND.n885 GND.n731 585
R566 GND.n888 GND.n887 585
R567 GND.n887 GND.n886 585
R568 GND.n889 GND.n723 585
R569 GND.n723 GND.n722 585
R570 GND.n891 GND.n890 585
R571 GND.n892 GND.n891 585
R572 GND.n721 GND.n720 585
R573 GND.n182 GND 583.907
R574 GND.n1018 GND.n213 582.4
R575 GND.n1102 GND.n134 576.293
R576 GND.n1102 GND.n133 576.293
R577 GND.n1082 GND.n151 576.293
R578 GND.n1083 GND.n1082 576.293
R579 GND.n1105 GND.n141 576.293
R580 GND.n1105 GND.n139 576.293
R581 GND.n1122 GND.n1121 568.095
R582 GND.n389 GND.n388 566.203
R583 GND.t246 GND.n302 562.423
R584 GND.n1117 GND.n143 542.871
R585 GND GND.t408 539.465
R586 GND GND.t215 539.465
R587 GND.n891 GND.n721 539.294
R588 GND.n891 GND.n723 539.294
R589 GND.n887 GND.n723 539.294
R590 GND.n887 GND.n731 539.294
R591 GND.n883 GND.n733 539.294
R592 GND.n879 GND.n733 539.294
R593 GND.n879 GND.n742 539.294
R594 GND.n875 GND.n742 539.294
R595 GND.n875 GND.n744 539.294
R596 GND.n867 GND.n753 539.294
R597 GND.n863 GND.n753 539.294
R598 GND.n863 GND.n755 539.294
R599 GND.n859 GND.n755 539.294
R600 GND.n859 GND.n763 539.294
R601 GND.n855 GND.n765 539.294
R602 GND.n851 GND.n765 539.294
R603 GND.n851 GND.n774 539.294
R604 GND.n847 GND.n774 539.294
R605 GND.n847 GND.n776 539.294
R606 GND.n839 GND.n785 539.294
R607 GND.n835 GND.n785 539.294
R608 GND.n835 GND.n787 539.294
R609 GND.n831 GND.n787 539.294
R610 GND.n831 GND.n795 539.294
R611 GND.n827 GND.n797 539.294
R612 GND.n823 GND.n797 539.294
R613 GND.n823 GND.n806 539.294
R614 GND.n819 GND.n806 539.294
R615 GND.n819 GND.n807 539.294
R616 GND.n1267 GND.n38 539.294
R617 GND.n1263 GND.n38 539.294
R618 GND.n1263 GND.n43 539.294
R619 GND.n1259 GND.n43 539.294
R620 GND.n1259 GND.n45 539.294
R621 GND.n1251 GND.n54 539.294
R622 GND.n1247 GND.n54 539.294
R623 GND.n1240 GND.n1239 539.294
R624 GND.n1239 GND.n59 539.294
R625 GND.n1234 GND.n1203 539.294
R626 GND.n1211 GND.n1203 539.294
R627 GND.n1225 GND.n1221 539.294
R628 GND.n1221 GND.n1220 539.294
R629 GND.n274 GND.n258 539.294
R630 GND.n283 GND.n260 539.294
R631 GND.n292 GND.n262 539.294
R632 GND.n944 GND.n265 539.294
R633 GND.n35 GND.t123 536.042
R634 GND.n30 GND.t506 536.042
R635 GND.n1132 GND.n1131 530.072
R636 GND.n423 GND.n422 525.178
R637 GND.n484 GND.n483 525.178
R638 GND GND.t133 522.606
R639 GND GND.t140 522.606
R640 GND.n1236 GND.n60 517.648
R641 GND.n939 GND.n213 516.841
R642 GND.n1109 GND.n1093 514.26
R643 GND.n1068 GND.n1058 514.26
R644 GND.n1054 GND.n175 514.26
R645 GND.n1176 GND.n92 514.26
R646 GND.n903 GND.n223 514.26
R647 GND.n1200 GND.n63 514.26
R648 GND.n89 GND.n86 514.26
R649 GND.n1200 GND.n1199 514.26
R650 GND.n1169 GND.n97 511.591
R651 GND.n1032 GND.n202 502.967
R652 GND.n929 GND.n909 502.967
R653 GND.t172 GND.t449 502.538
R654 GND.n1032 GND.n195 499.784
R655 GND.n929 GND.n194 499.784
R656 GND.n906 GND.n185 499.784
R657 GND.n920 GND.n186 499.784
R658 GND.n909 GND.n906 496.601
R659 GND.n920 GND.n916 496.601
R660 GND.n1118 GND.n142 496.188
R661 GND.n1090 GND.n157 494.683
R662 GND.n375 GND.n374 492.817
R663 GND.t123 GND.n25 491.372
R664 GND.n1084 GND.n157 487.154
R665 GND.n1114 GND.n145 483.003
R666 GND.t197 GND.t507 480.461
R667 GND.t243 GND.t423 480.204
R668 GND.n1108 GND.n1107 475.86
R669 GND.n1164 GND.n1163 475.536
R670 GND.n1077 GND.t72 473.488
R671 GND.n931 GND.n192 472.848
R672 GND.n1044 GND.n192 472.848
R673 GND.n1092 GND.n1091 472.471
R674 GND GND.t446 472.031
R675 GND.n935 GND.n194 471.134
R676 GND.n1020 GND.n210 471.134
R677 GND.t358 GND.t591 470.267
R678 GND.t245 GND.t336 470.267
R679 GND.t196 GND.t195 470.267
R680 GND.t357 GND.t356 470.267
R681 GND.t515 GND.t257 470.267
R682 GND.t594 GND.t593 470.267
R683 GND.t248 GND.t247 470.267
R684 GND GND.t78 469.036
R685 GND.n376 GND.n375 461.243
R686 GND.n388 GND.n387 461.243
R687 GND.n1115 GND.n1114 461.243
R688 GND.n1142 GND.n120 461.243
R689 GND.n949 GND.n948 461.243
R690 GND.n1143 GND.n1142 459.964
R691 GND.n1131 GND.n1130 459.671
R692 GND.n1123 GND.n137 459.671
R693 GND.n1009 GND.n217 459.295
R694 GND.n218 GND.n217 459.295
R695 GND.n948 GND.n257 459.111
R696 GND.n1164 GND.n103 458.043
R697 GND.t243 GND.t427 457.868
R698 GND.n371 GND.n370 449.296
R699 GND.n32 GND.t170 446.745
R700 GND.t170 GND.n31 446.745
R701 GND.t184 GND.n25 446.702
R702 GND.n183 GND.n181 443.86
R703 GND.n183 GND.n182 443.86
R704 GND.n1064 GND.n74 443.86
R705 GND.n1064 GND.n1063 443.86
R706 GND.n1172 GND.n95 443.86
R707 GND.n998 GND.n223 443.86
R708 GND.n997 GND.n996 443.86
R709 GND.n996 GND.n225 443.86
R710 GND.n967 GND.n239 443.86
R711 GND.n1177 GND.n1176 443.86
R712 GND.n1192 GND.n1191 443.86
R713 GND.n1188 GND.n75 443.86
R714 GND.n86 GND.n82 443.86
R715 GND.n1199 GND.n1198 443.86
R716 GND.n1197 GND.n1196 443.86
R717 GND.n1196 GND.n68 443.86
R718 GND.n232 GND.n231 443.86
R719 GND.n231 GND.n85 443.86
R720 GND.n1181 GND.n1180 443.86
R721 GND.n1180 GND.n1179 443.86
R722 GND.t361 GND 442.539
R723 GND GND.t614 442.539
R724 GND GND.t20 442.539
R725 GND.n1091 GND.n1090 438.966
R726 GND.n1118 GND.n1117 438.966
R727 GND.n1294 GND.t107 438.315
R728 GND.n1271 GND.n1270 436.238
R729 GND.n1109 GND.n1108 435.577
R730 GND.n1069 GND.n1057 431.812
R731 GND.n924 GND.n910 430.252
R732 GND.n1181 GND.n85 428.8
R733 GND.n967 GND.n966 427.671
R734 GND.n137 GND.n129 415.248
R735 GND.n1107 GND.n142 415.248
R736 GND.n1189 GND.n1188 414.872
R737 GND.t507 GND 413.027
R738 GND.n1062 GND.n82 399.812
R739 GND GND.n74 399.06
R740 GND.n1093 GND.n1092 397.176
R741 GND.n387 GND.n386 390.416
R742 GND.n239 GND.n225 380.988
R743 GND.n990 GND.n989 380.988
R744 GND.n1076 GND.n1075 380.676
R745 GND.n1139 GND.n1138 375.947
R746 GND.t249 GND.n34 370.882
R747 GND.n1322 GND.t408 370.882
R748 GND.n1310 GND.t603 370.882
R749 GND.t389 GND.n1309 370.882
R750 GND.n218 GND.n204 364.048
R751 GND GND.n371 362.88
R752 GND.n31 GND.t438 362.454
R753 GND.n1170 GND.n1169 361.601
R754 GND.n1198 GND.n64 350.872
R755 GND.n1197 GND.n66 350.872
R756 GND.n230 GND.n68 350.872
R757 GND.n991 GND.n232 350.872
R758 GND.n988 GND.n85 350.872
R759 GND.n1181 GND.n83 350.872
R760 GND.n1179 GND.n1178 350.872
R761 GND.n1030 GND.n203 350.168
R762 GND.n1030 GND.n202 346.983
R763 GND.n903 GND.n64 345.976
R764 GND.n1124 GND.n1123 343.341
R765 GND.n1122 GND.n136 343.341
R766 GND.n972 GND.t192 342.896
R767 GND.n1191 GND.n1190 338.825
R768 GND.n232 GND.n68 338.825
R769 GND.n34 GND.t262 337.166
R770 GND.t520 GND.n1322 337.166
R771 GND.n1310 GND.t319 337.166
R772 GND.n1309 GND.t477 337.166
R773 GND GND.t249 335.026
R774 GND.n181 GND.n180 332.8
R775 GND.n182 GND.n71 332.8
R776 GND.n1189 GND.n74 332.8
R777 GND.n1063 GND.n1062 332.8
R778 GND.n915 GND.n201 330.865
R779 GND.t591 GND.t89 328.938
R780 GND.t105 GND.t245 328.938
R781 GND.t336 GND.t589 328.938
R782 GND.t560 GND.t196 328.938
R783 GND.t195 GND.t299 328.938
R784 GND.t332 GND.t357 328.938
R785 GND.t356 GND.t626 328.938
R786 GND.t257 GND.t471 328.938
R787 GND.t260 GND.t515 328.938
R788 GND.t493 GND.t594 328.938
R789 GND.t593 GND.t501 328.938
R790 GND.t401 GND.t248 328.938
R791 GND.t479 GND.t197 328.736
R792 GND.n998 GND.n997 317.365
R793 GND.n229 GND.n222 317.365
R794 GND.n180 GND.n179 313.601
R795 GND.n390 GND.n389 312.353
R796 GND.n222 GND.n66 310.589
R797 GND.n1121 GND.n138 306.825
R798 GND.t523 GND.t202 304.7
R799 GND.t128 GND.t69 304.7
R800 GND GND.n129 303.06
R801 GND.n179 GND.n178 301.553
R802 GND.n1198 GND.n1197 301.553
R803 GND.n392 GND.n391 299.553
R804 GND.n138 GND 298.918
R805 GND.t158 GND 296.161
R806 GND.n1172 GND.n1171 295.906
R807 GND GND.t520 295.019
R808 GND.n1055 GND.n1054 294.776
R809 GND.n1014 GND.n212 291.205
R810 GND.t7 GND.t136 290.19
R811 GND.t634 GND.t383 290.19
R812 GND.t67 GND.t527 290.19
R813 GND.n991 GND.n990 289.13
R814 GND.n1049 GND.n187 281.601
R815 GND.t524 GND.t633 275.68
R816 GND.t632 GND.t391 275.68
R817 GND.t5 GND.t88 275.68
R818 GND.n1287 GND.t216 274.812
R819 GND.n1315 GND.t92 274.812
R820 GND.n680 GND.t139 274.812
R821 GND.n669 GND.t157 274.812
R822 GND.n178 GND.n71 272.565
R823 GND.t292 GND 269.733
R824 GND.t603 GND 269.733
R825 GND.n377 GND.n376 259.873
R826 GND.n230 GND.n229 259.765
R827 GND GND.t385 256.853
R828 GND.n1038 GND.n197 256.753
R829 GND.t136 GND 253.917
R830 GND.t202 GND 253.917
R831 GND.t168 GND 253.917
R832 GND.t383 GND 253.917
R833 GND GND.t270 253.917
R834 GND GND.t405 253.917
R835 GND.t527 GND 253.917
R836 GND.t69 GND 253.917
R837 GND.t345 GND 253.917
R838 GND.n391 GND.n390 253.26
R839 GND GND.t389 252.875
R840 GND.t439 GND 252.875
R841 GND.t578 GND 252.875
R842 GND.n395 GND.n145 251.339
R843 GND.n397 GND.n396 249.207
R844 GND.t270 GND.n417 246.237
R845 GND.n1151 GND.t220 242.202
R846 GND.n1024 GND.n208 241.319
R847 GND.n90 GND.n83 241.319
R848 GND.n1055 GND.n174 240.565
R849 GND.n1070 GND.n1069 240.565
R850 GND.n1048 GND.n188 237.177
R851 GND.t215 GND 236.016
R852 GND.n962 GND.n96 235.98
R853 GND.n1044 GND.n188 235.672
R854 GND GND.t93 232.153
R855 GND.t6 GND.n416 232.153
R856 GND.n487 GND.t632 232.153
R857 GND.t273 GND 232.153
R858 GND.n430 GND.t68 232.153
R859 GND.n429 GND.t5 232.153
R860 GND GND.t264 232.153
R861 GND.n515 GND.t432 232.153
R862 GND.t633 GND.n418 230.849
R863 GND.n399 GND.n398 229.579
R864 GND.n419 GND.t523 228.524
R865 GND.n428 GND.t128 228.524
R866 GND.t335 GND.t334 228.131
R867 GND.t193 GND.t194 228.131
R868 GND.n394 GND.n393 226.544
R869 GND.n988 GND.n987 226.26
R870 GND.t1 GND.t237 224.898
R871 GND.t641 GND.t480 224.898
R872 GND.t152 GND.t618 224.898
R873 GND.n914 GND.t514 222.188
R874 GND.n214 GND.t466 222.023
R875 GND.n214 GND.t615 221.905
R876 GND.n206 GND.t431 221.851
R877 GND.n206 GND.t467 221.851
R878 GND.n1036 GND.t272 221.738
R879 GND.n989 GND.n988 217.601
R880 GND.n419 GND 214.016
R881 GND GND.n486 214.016
R882 GND GND.n428 214.016
R883 GND.t421 GND.t524 210.387
R884 GND.t93 GND.t347 210.387
R885 GND.t391 GND.t79 210.387
R886 GND.t171 GND.t273 210.387
R887 GND.t88 GND.t147 210.387
R888 GND.t264 GND.t235 210.387
R889 GND.n242 GND.n241 207.393
R890 GND.n524 GND.t358 205.118
R891 GND.n987 GND.n83 202.542
R892 GND.n1008 GND.n208 201.788
R893 GND.n945 GND.n263 200.215
R894 GND.n945 GND.n261 200.215
R895 GND.n945 GND.n259 200.215
R896 GND.n945 GND.n264 200.215
R897 GND.n374 GND.n366 196.726
R898 GND.n644 GND.n638 196.256
R899 GND.t290 GND.t168 195.879
R900 GND.t405 GND.t150 195.879
R901 GND.t518 GND.t345 195.879
R902 GND.n1171 GND.n92 195.766
R903 GND.n1184 GND.n79 195.395
R904 GND.n370 GND.n365 192.034
R905 GND.n1167 GND.n1166 189.688
R906 GND.n396 GND.n395 188.194
R907 GND.t639 GND 185.441
R908 GND.t107 GND 185.441
R909 GND.n486 GND.n417 184.678
R910 GND.n292 GND.n263 184.572
R911 GND.n283 GND.n261 184.572
R912 GND.n274 GND.n259 184.572
R913 GND.n265 GND.n264 184.572
R914 GND.n386 GND.n157 184.471
R915 GND.n1091 GND.n156 184.471
R916 GND.n1093 GND.n152 184.471
R917 GND.n1108 GND.n1100 184.471
R918 GND.n1097 GND.n142 184.471
R919 GND.n1117 GND.n1116 184.471
R920 GND.n992 GND.n230 184.095
R921 GND.n526 GND.t359 183.065
R922 GND.n359 GND.t628 183.065
R923 GND.n355 GND.t486 183.065
R924 GND.n351 GND.t547 183.065
R925 GND.n347 GND.t101 183.065
R926 GND.n343 GND.t9 183.065
R927 GND.n339 GND.t574 183.065
R928 GND.n335 GND.t583 183.065
R929 GND.t558 GND.n629 183.065
R930 GND.t129 GND.n630 183.065
R931 GND.n1162 GND.n1161 180.087
R932 GND.n400 GND.n399 179.019
R933 GND.n1116 GND.n1115 179.004
R934 GND.t484 GND.t579 178.68
R935 GND.n932 GND.n187 175.06
R936 GND.n385 GND.n384 173.474
R937 GND.n212 GND.n197 172.746
R938 GND.n246 GND.n245 172.619
R939 GND.n252 GND.n251 171.554
R940 GND.n115 GND.n114 171.339
R941 GND.n1149 GND.n1148 171.339
R942 GND.n963 GND.n962 171.339
R943 GND.n256 GND.n255 171.339
R944 GND.n951 GND.n950 171.339
R945 GND.n955 GND.n954 171.339
R946 GND.n1192 GND.n71 171.294
R947 GND.n1158 GND.n1157 171.126
R948 GND.n1096 GND.n144 170.487
R949 GND.n1095 GND.n1094 170.274
R950 GND.n119 GND.n118 170.274
R951 GND.n110 GND.n109 170.274
R952 GND.n106 GND.n105 170.274
R953 GND.n960 GND.n959 170.274
R954 GND.n1145 GND.n1144 170.06
R955 GND.n219 GND.n64 168.282
R956 GND.n373 GND.n372 163.874
R957 GND.n530 GND.t360 162.471
R958 GND.n535 GND.t283 162.471
R959 GND.n541 GND.t629 162.471
R960 GND.n546 GND.t414 162.471
R961 GND.n552 GND.t487 162.471
R962 GND.n557 GND.t638 162.471
R963 GND.n563 GND.t548 162.471
R964 GND.n568 GND.t296 162.471
R965 GND.n574 GND.t102 162.471
R966 GND.n579 GND.t205 162.471
R967 GND.n585 GND.t10 162.471
R968 GND.n590 GND.t373 162.471
R969 GND.n596 GND.t575 162.471
R970 GND.n601 GND.t563 162.471
R971 GND.n607 GND.t584 162.471
R972 GND.n612 GND.t71 162.471
R973 GND.n331 GND.t559 162.471
R974 GND.n622 GND.t302 162.471
R975 GND.n1387 GND.t130 162.471
R976 GND.n1384 GND.t396 162.471
R977 GND.n369 GND.n125 161.903
R978 GND GND.t282 161.149
R979 GND GND.t413 161.149
R980 GND GND.t637 161.149
R981 GND GND.t295 161.149
R982 GND GND.t204 161.149
R983 GND GND.t372 161.149
R984 GND GND.t562 161.149
R985 GND GND.t70 161.149
R986 GND.t301 GND 161.149
R987 GND.t395 GND 161.149
R988 GND.n534 GND.t496 160.017
R989 GND.n358 GND.t285 160.017
R990 GND.n545 GND.t451 160.017
R991 GND.n354 GND.t240 160.017
R992 GND.n556 GND.t331 160.017
R993 GND.n350 GND.t455 160.017
R994 GND.n567 GND.t550 160.017
R995 GND.n346 GND.t298 160.017
R996 GND.n578 GND.t104 160.017
R997 GND.n342 GND.t207 160.017
R998 GND.n589 GND.t234 160.017
R999 GND.n338 GND.t375 160.017
R1000 GND.n600 GND.t577 160.017
R1001 GND.n334 GND.t565 160.017
R1002 GND.n611 GND.t448 160.017
R1003 GND.n330 GND.t112 160.017
R1004 GND.n623 GND.t142 160.017
R1005 GND.n618 GND.t304 160.017
R1006 GND.n1385 GND.t132 160.017
R1007 GND.n5 GND.t398 160.017
R1008 GND.t341 GND.t335 159.571
R1009 GND.t334 GND.t18 159.571
R1010 GND.t194 GND.t456 159.571
R1011 GND.t387 GND.t193 159.571
R1012 GND.t178 GND.t592 159.571
R1013 GND.n1275 GND.t160 158.361
R1014 GND.n1282 GND.t198 158.361
R1015 GND.n20 GND.t504 158.361
R1016 GND.n22 GND.t173 158.361
R1017 GND.n650 GND.t526 158.361
R1018 GND.n1354 GND.t231 155.63
R1019 GND.n992 GND.n991 154.73
R1020 GND.n1352 GND.t622 154.131
R1021 GND.n1329 GND.t424 154.131
R1022 GND.n272 GND.t611 153.707
R1023 GND.n1331 GND.t244 153.631
R1024 GND.n718 GND.n717 153.276
R1025 GND.n1332 GND.t428 152.381
R1026 GND.n1099 GND.n1098 152.139
R1027 GND.n152 GND.n148 151.779
R1028 GND.n1294 GND 151.725
R1029 GND.n250 GND.n249 151.714
R1030 GND.n155 GND.n154 151.5
R1031 GND.n117 GND.n116 151.5
R1032 GND.n108 GND.n107 151.5
R1033 GND.n1147 GND.n1146 151.5
R1034 GND.n953 GND.n952 151.5
R1035 GND.n957 GND.n956 151.5
R1036 GND.n643 GND.n642 151.256
R1037 GND.n644 GND.n643 151.256
R1038 GND.n641 GND.n640 151.256
R1039 GND.n642 GND.n641 151.256
R1040 GND.n639 GND.n323 151.256
R1041 GND.n640 GND.n639 151.256
R1042 GND.n326 GND.n321 151.256
R1043 GND.n326 GND.n323 151.256
R1044 GND.n320 GND.n319 151.256
R1045 GND.n321 GND.n320 151.256
R1046 GND.n318 GND.n317 151.256
R1047 GND.n319 GND.n318 151.256
R1048 GND.n711 GND.n304 151.256
R1049 GND.n317 GND.n304 151.256
R1050 GND.n714 GND.n301 151.256
R1051 GND.n714 GND.n713 151.256
R1052 GND.n713 GND.n712 151.256
R1053 GND.n712 GND.n711 151.256
R1054 GND.n717 GND.n301 151.256
R1055 GND.n1298 GND.t214 150.922
R1056 GND.n1302 GND.t640 150.922
R1057 GND.n1303 GND.t318 150.922
R1058 GND.n1289 GND.t478 150.922
R1059 GND.n1288 GND.t320 150.922
R1060 GND.n1359 GND.t485 150.922
R1061 GND.n1347 GND.t263 150.922
R1062 GND.n1343 GND.t386 150.922
R1063 GND.n1338 GND.t185 150.922
R1064 GND.n1297 GND.t108 150.922
R1065 GND.n663 GND.t418 150.922
R1066 GND.n658 GND.t644 150.922
R1067 GND.n442 GND.t642 150.922
R1068 GND.n505 GND.t238 150.922
R1069 GND.n492 GND.t169 150.922
R1070 GND.n498 GND.t203 150.922
R1071 GND.n410 GND.t137 150.922
R1072 GND.n450 GND.t582 150.922
R1073 GND.n456 GND.t406 150.922
R1074 GND.n364 GND.t346 150.922
R1075 GND.n479 GND.t382 150.922
R1076 GND.n469 GND.t528 150.922
R1077 GND.n425 GND.t153 150.922
R1078 GND.n444 GND.t384 150.922
R1079 GND.n254 GND.n253 150.434
R1080 GND.n1354 GND.t321 149.493
R1081 GND.n1272 GND.t409 149.493
R1082 GND.n965 GND.n961 149.367
R1083 GND.n1056 GND.n1055 149.083
R1084 GND.n279 GND.t340 149.067
R1085 GND.n288 GND.t580 149.067
R1086 GND.n297 GND.t353 149.067
R1087 GND.n726 GND.t453 149.067
R1088 GND.n736 GND.t82 149.067
R1089 GND.n746 GND.t276 149.067
R1090 GND.n870 GND.t39 149.067
R1091 GND.n758 GND.t517 149.067
R1092 GND.n768 GND.t459 149.067
R1093 GND.n778 GND.t537 149.067
R1094 GND.n842 GND.t17 149.067
R1095 GND.n790 GND.t228 149.067
R1096 GND.n800 GND.t15 149.067
R1097 GND.n809 GND.t573 149.067
R1098 GND.n814 GND.t596 149.067
R1099 GND.n47 GND.t84 149.067
R1100 GND.n1254 GND.t294 149.067
R1101 GND.n1243 GND.t117 149.067
R1102 GND.n1207 GND.t500 149.067
R1103 GND.n1228 GND.t367 149.067
R1104 GND.n1216 GND.t200 149.067
R1105 GND.n1160 GND.n1159 148.087
R1106 GND.n1361 GND.t530 147.411
R1107 GND.n143 GND.n140 146.25
R1108 GND.n140 GND.n126 146.25
R1109 GND.n132 GND.n131 146.25
R1110 GND.n1081 GND.n132 146.25
R1111 GND.n1102 GND.n130 146.25
R1112 GND.n1103 GND.n1102 146.25
R1113 GND.n1133 GND.n1132 146.25
R1114 GND.n1134 GND.n1133 146.25
R1115 GND.n1084 GND.n158 146.25
R1116 GND.n1075 GND.n158 146.25
R1117 GND.n1082 GND.n153 146.25
R1118 GND.n1082 GND.n1081 146.25
R1119 GND.n1106 GND.n1105 146.25
R1120 GND.n1105 GND.n1104 146.25
R1121 GND.n1071 GND.n170 146.25
R1122 GND.n170 GND.n159 146.25
R1123 GND.n1060 GND.n1059 146.25
R1124 GND.n1060 GND.n167 146.25
R1125 GND.n1061 GND.n1058 146.25
R1126 GND.n1061 GND.n160 146.25
R1127 GND.n233 GND.n228 146.25
R1128 GND.n237 GND.n228 146.25
R1129 GND.n235 GND.n234 146.25
R1130 GND.n238 GND.n235 146.25
R1131 GND.n240 GND.n236 146.25
R1132 GND.n984 GND.n236 146.25
R1133 GND.n93 GND.n91 146.25
R1134 GND.n981 GND.n93 146.25
R1135 GND.n94 GND.n92 146.25
R1136 GND.n76 GND.n73 146.25
R1137 GND.n164 GND.n76 146.25
R1138 GND.n84 GND.n77 146.25
R1139 GND.n1185 GND.n77 146.25
R1140 GND.n1183 GND.n1182 146.25
R1141 GND.n1184 GND.n1183 146.25
R1142 GND.n72 GND.n70 146.25
R1143 GND.n165 GND.n70 146.25
R1144 GND.n89 GND.n88 146.25
R1145 GND.n1201 GND.n1200 146.25
R1146 GND.n904 GND.n903 146.25
R1147 GND.n905 GND.n904 146.25
R1148 GND.n1000 GND.n999 146.25
R1149 GND.n1001 GND.n1000 146.25
R1150 GND.n227 GND.n224 146.25
R1151 GND.n227 GND.n226 146.25
R1152 GND.n907 GND.n65 146.25
R1153 GND.n908 GND.n907 146.25
R1154 GND.n69 GND.n67 146.25
R1155 GND.n922 GND.n69 146.25
R1156 GND.n176 GND.n175 146.25
R1157 GND.n902 GND.n176 146.25
R1158 GND.n177 GND.n173 146.25
R1159 GND.n1002 GND.n177 146.25
R1160 GND.n171 GND.n169 146.25
R1161 GND.n918 GND.n169 146.25
R1162 GND.n1030 GND.n1029 146.25
R1163 GND.n1031 GND.n1030 146.25
R1164 GND.n1362 GND.t613 146.245
R1165 GND.t188 GND.n982 144.454
R1166 GND.n398 GND.n397 143.393
R1167 GND.n244 GND.n243 142.754
R1168 GND.n156 GND.n155 138.897
R1169 GND.n699 GND.t222 137.728
R1170 GND.n113 GND.n112 137.47
R1171 GND.n105 GND.n103 137.419
R1172 GND.n241 GND.n97 135.286
R1173 GND.n393 GND.n392 135.073
R1174 GND.n219 GND.n66 133.272
R1175 GND.n1100 GND.n1099 133.137
R1176 GND.n1154 GND.n1150 132.907
R1177 GND.n378 GND.n373 132.071
R1178 GND.n386 GND.n385 131.857
R1179 GND.n180 GND.n63 130.26
R1180 GND.n243 GND.n242 128.887
R1181 GND.n897 GND.t121 127.977
R1182 GND.n1097 GND.n1096 125.457
R1183 GND.t525 GND 125.046
R1184 GND.n893 GND.n721 121.496
R1185 GND.n1116 GND.n144 120.55
R1186 GND.n383 GND.n365 117.99
R1187 GND.n936 GND.n935 117.001
R1188 GND.n935 GND.n934 117.001
R1189 GND.n929 GND.n928 117.001
R1190 GND.n934 GND.n929 117.001
R1191 GND.n1020 GND.n1019 117.001
R1192 GND.n1021 GND.n1020 117.001
R1193 GND.n1033 GND.n1032 117.001
R1194 GND.n1032 GND.n1031 117.001
R1195 GND.n911 GND.n906 117.001
R1196 GND.n934 GND.n906 117.001
R1197 GND.n920 GND.n919 117.001
R1198 GND.n921 GND.n920 117.001
R1199 GND.n1132 GND.n129 114.825
R1200 GND.n1013 GND.n208 111.812
R1201 GND.n384 GND.n156 110.311
R1202 GND.t347 GND.t290 108.822
R1203 GND.t150 GND.t171 108.822
R1204 GND.t235 GND.t518 108.822
R1205 GND.t359 GND.t495 108.293
R1206 GND.t282 GND.t284 108.293
R1207 GND.t628 GND.t450 108.293
R1208 GND.t413 GND.t239 108.293
R1209 GND.t486 GND.t330 108.293
R1210 GND.t637 GND.t454 108.293
R1211 GND.t547 GND.t549 108.293
R1212 GND.t295 GND.t297 108.293
R1213 GND.t101 GND.t103 108.293
R1214 GND.t204 GND.t206 108.293
R1215 GND.t9 GND.t233 108.293
R1216 GND.t372 GND.t374 108.293
R1217 GND.t574 GND.t576 108.293
R1218 GND.t562 GND.t564 108.293
R1219 GND.t583 GND.t447 108.293
R1220 GND.t70 GND.t111 108.293
R1221 GND.t141 GND.t558 108.293
R1222 GND.t303 GND.t301 108.293
R1223 GND.t131 GND.t129 108.293
R1224 GND.t397 GND.t395 108.293
R1225 GND.n1098 GND.n1097 106.257
R1226 GND.n516 GND.n302 106.16
R1227 GND.n1163 GND.n1162 102.433
R1228 GND.n654 GND.t392 102.377
R1229 GND.n372 GND 100.496
R1230 GND.n964 GND.n963 100.299
R1231 GND.n1170 GND.n96 99.6436
R1232 GND.n924 GND.n915 99.3887
R1233 GND.n983 GND.t40 99.2212
R1234 GND.n1161 GND.n1160 98.1667
R1235 GND GND.n359 96.6896
R1236 GND GND.n355 96.6896
R1237 GND GND.n351 96.6896
R1238 GND GND.n347 96.6896
R1239 GND GND.n343 96.6896
R1240 GND GND.n339 96.6896
R1241 GND GND.n335 96.6896
R1242 GND.n629 GND 96.6896
R1243 GND.n630 GND 96.6896
R1244 GND.n1100 GND.n1095 96.4436
R1245 GND.n1371 GND.n1370 96.2411
R1246 GND.n961 GND.n960 96.0333
R1247 GND.n1025 GND.n204 95.2476
R1248 GND.t237 GND.t421 94.3121
R1249 GND.t79 GND.t641 94.3121
R1250 GND.t147 GND.t152 94.3121
R1251 GND.t255 GND 89.9457
R1252 GND.n522 GND.n521 89.504
R1253 GND GND.t415 89.2144
R1254 GND.n154 GND.n152 88.9769
R1255 GND.n717 GND.n716 88.7516
R1256 GND.t495 GND 86.3761
R1257 GND.t284 GND 86.3761
R1258 GND.t450 GND 86.3761
R1259 GND.t239 GND 86.3761
R1260 GND.t330 GND 86.3761
R1261 GND.t454 GND 86.3761
R1262 GND.t549 GND 86.3761
R1263 GND.t297 GND 86.3761
R1264 GND.t103 GND 86.3761
R1265 GND.t206 GND 86.3761
R1266 GND.t233 GND 86.3761
R1267 GND.t374 GND 86.3761
R1268 GND.t576 GND 86.3761
R1269 GND.t564 GND 86.3761
R1270 GND.t447 GND 86.3761
R1271 GND.t111 GND 86.3761
R1272 GND GND.t141 86.3761
R1273 GND GND.t303 86.3761
R1274 GND GND.t131 86.3761
R1275 GND GND.t397 86.3761
R1276 GND.n699 GND 86.3761
R1277 GND.n969 GND.t186 85.3595
R1278 GND.n245 GND.n244 84.94
R1279 GND.n107 GND.n106 82.8067
R1280 GND.n109 GND.n108 80.6733
R1281 GND.n1171 GND.n1170 80.0005
R1282 GND.n966 GND.n965 80.0005
R1283 GND GND.t525 77.5142
R1284 GND.n974 GND.t48 74.416
R1285 GND.n966 GND.n240 74.0272
R1286 GND.t325 GND.t540 72.1616
R1287 GND.t329 GND.t569 72.1616
R1288 GND.t569 GND.t252 72.1616
R1289 GND.t252 GND.t326 72.1616
R1290 GND.t326 GND.t539 72.1616
R1291 GND.t539 GND.t328 72.1616
R1292 GND.t567 GND.t328 72.1616
R1293 GND.t567 GND.t538 72.1616
R1294 GND.t568 GND.t538 72.1616
R1295 GND.t542 GND.t568 72.1616
R1296 GND.t566 GND.t542 72.1616
R1297 GND.t327 GND.t251 72.1616
R1298 GND.t541 GND.t327 72.1616
R1299 GND.t250 GND.t541 72.1616
R1300 GND.t163 GND.t161 72.1616
R1301 GND.t161 GND.t269 72.1616
R1302 GND.t269 GND.t162 72.1616
R1303 GND.t460 GND.t490 72.1616
R1304 GND.t36 GND.t28 72.1616
R1305 GND.t43 GND.t36 72.1616
R1306 GND.t35 GND.t43 72.1616
R1307 GND.n1159 GND.n1158 72.14
R1308 GND.n1157 GND.n1156 72.14
R1309 GND.n956 GND.n955 72.14
R1310 GND.n1182 GND.n82 70.4005
R1311 GND.n1182 GND.n1181 70.4005
R1312 GND.n84 GND.n75 70.4005
R1313 GND.n85 GND.n84 70.4005
R1314 GND.n1190 GND.n73 70.4005
R1315 GND.n232 GND.n73 70.4005
R1316 GND.n1092 GND.n153 70.4005
R1317 GND.n1086 GND.n153 70.4005
R1318 GND.n1107 GND.n1106 70.4005
R1319 GND.n1106 GND.n136 70.4005
R1320 GND.n135 GND.n131 70.4005
R1321 GND.n1123 GND.n130 70.4005
R1322 GND.n1130 GND.n130 70.4005
R1323 GND.n1071 GND.n1070 70.4005
R1324 GND.n174 GND.n171 70.4005
R1325 GND.n1056 GND.n173 70.4005
R1326 GND.n182 GND.n173 70.4005
R1327 GND.n1059 GND.n1057 70.4005
R1328 GND.n1059 GND.n74 70.4005
R1329 GND.n1063 GND.n1058 70.4005
R1330 GND.n181 GND.n175 70.4005
R1331 GND.n240 GND.n90 70.4005
R1332 GND.n1177 GND.n91 70.4005
R1333 GND.n95 GND.n91 70.4005
R1334 GND.n999 GND.n222 70.4005
R1335 GND.n999 GND.n998 70.4005
R1336 GND.n229 GND.n224 70.4005
R1337 GND.n997 GND.n224 70.4005
R1338 GND.n990 GND.n233 70.4005
R1339 GND.n233 GND.n225 70.4005
R1340 GND.n989 GND.n234 70.4005
R1341 GND.n239 GND.n234 70.4005
R1342 GND.n1191 GND.n72 70.4005
R1343 GND.n72 GND.n68 70.4005
R1344 GND.n178 GND.n67 70.4005
R1345 GND.n1197 GND.n67 70.4005
R1346 GND.n179 GND.n65 70.4005
R1347 GND.n1198 GND.n65 70.4005
R1348 GND.n1179 GND.n89 70.4005
R1349 GND.t113 GND.t158 70.2016
R1350 GND.t127 GND.t255 70.2016
R1351 GND.n383 GND.n366 69.7769
R1352 GND.n32 GND.t503 69.7227
R1353 GND.n1271 GND 69.4703
R1354 GND.t45 GND.t329 69.0242
R1355 GND.n253 GND.n252 67.4467
R1356 GND.t446 GND.t91 67.4335
R1357 GND.t133 GND.t317 67.4335
R1358 GND.t140 GND.t213 67.4335
R1359 GND.n1373 GND.n11 67.2766
R1360 GND.n247 GND.n246 66.9708
R1361 GND.n1077 GND.n1076 65.8868
R1362 GND.n959 GND.n958 65.3297
R1363 GND.n111 GND.n110 65.3133
R1364 GND.n251 GND.n250 65.3133
R1365 GND.n939 GND.n938 65.1299
R1366 GND.n31 GND 65.0093
R1367 GND.n1013 GND.n1012 65.0005
R1368 GND.n1012 GND.n163 65.0005
R1369 GND.t410 GND.t268 64.841
R1370 GND.t412 GND.t488 64.841
R1371 GND.t95 GND.t648 64.841
R1372 GND.n1033 GND.n201 64.377
R1373 GND.n911 GND.n187 64.0005
R1374 GND.n928 GND.n910 64.0005
R1375 GND.n928 GND.n196 64.0005
R1376 GND.n1033 GND.n197 64.0005
R1377 GND.n919 GND.n188 64.0005
R1378 GND.n911 GND.n910 63.624
R1379 GND.n919 GND.n915 63.624
R1380 GND.n114 GND.n113 63.18
R1381 GND.n952 GND.n951 63.18
R1382 GND.t138 GND.t113 61.4265
R1383 GND.t156 GND.t127 61.4265
R1384 GND.t392 GND.t417 61.4265
R1385 GND.t415 GND.t643 61.4265
R1386 GND.n1150 GND.n1149 61.0467
R1387 GND.n1148 GND.n1147 61.0467
R1388 GND.n954 GND.n953 61.0467
R1389 GND.n1019 GND.n212 60.6123
R1390 GND.t149 GND.n973 60.5543
R1391 GND.n936 GND.n196 60.2358
R1392 GND.t411 GND.n149 60.1348
R1393 GND.n116 GND.n115 58.9133
R1394 GND.n255 GND.n254 58.9133
R1395 GND.n257 GND.n256 58.9133
R1396 GND.t469 GND.t647 57.5203
R1397 GND.t625 GND.t645 57.5203
R1398 GND.t468 GND.t646 57.5203
R1399 GND.t437 GND.t144 57.5203
R1400 GND.t607 GND.t604 56.9878
R1401 GND.n118 GND.n117 56.78
R1402 GND.n1075 GND.t325 55.6901
R1403 GND.n1081 GND.t250 55.6901
R1404 GND.n654 GND 55.5764
R1405 GND.t89 GND.n362 55.0318
R1406 GND.n362 GND.t105 55.0318
R1407 GND.n708 GND.t589 55.0318
R1408 GND.n708 GND.t560 55.0318
R1409 GND.t299 GND.n707 55.0318
R1410 GND.n707 GND.t332 55.0318
R1411 GND.t626 GND.n706 55.0318
R1412 GND.n706 GND.t471 55.0318
R1413 GND.n327 GND.t260 55.0318
R1414 GND.n327 GND.t493 55.0318
R1415 GND.n700 GND.t501 55.0318
R1416 GND.n700 GND.t401 55.0318
R1417 GND.t34 GND.t511 54.9057
R1418 GND.t25 GND.t277 54.9057
R1419 GND.n33 GND 54.7689
R1420 GND.n1146 GND.n1145 54.6467
R1421 GND.n1144 GND.n1143 54.6467
R1422 GND.n950 GND.n949 54.6467
R1423 GND GND.n11 54.1138
R1424 GND.n120 GND.n119 52.0867
R1425 GND.t279 GND.t37 52.0297
R1426 GND.t417 GND 51.1888
R1427 GND.t643 GND 51.1888
R1428 GND.t470 GND.t512 50.1996
R1429 GND.t75 GND.t22 50.1996
R1430 GND GND.t138 46.8012
R1431 GND GND.t156 46.8012
R1432 GND.n1029 GND.n204 46.3064
R1433 GND.t162 GND.t8 46.0163
R1434 GND.n520 GND.n517 45.7159
R1435 GND.n308 GND.n306 45.7159
R1436 GND.n710 GND.n709 45.7159
R1437 GND.n316 GND.n309 45.7159
R1438 GND.n705 GND.n704 45.7159
R1439 GND.n703 GND.n313 45.7159
R1440 GND.n702 GND.n701 45.7159
R1441 GND.n636 GND.n325 45.7159
R1442 GND.n696 GND.n695 45.7159
R1443 GND.n694 GND.n633 45.7159
R1444 GND.n1029 GND.n201 45.5534
R1445 GND.n362 GND.n308 45.0005
R1446 GND.n709 GND.n708 45.0005
R1447 GND.n707 GND.n309 45.0005
R1448 GND.n706 GND.n705 45.0005
R1449 GND.n327 GND.n313 45.0005
R1450 GND.n701 GND.n700 45.0005
R1451 GND.n712 GND.n303 45.0005
R1452 GND.n362 GND.n303 45.0005
R1453 GND.n310 GND.n304 45.0005
R1454 GND.n708 GND.n310 45.0005
R1455 GND.n318 GND.n311 45.0005
R1456 GND.n707 GND.n311 45.0005
R1457 GND.n320 GND.n312 45.0005
R1458 GND.n706 GND.n312 45.0005
R1459 GND.n328 GND.n326 45.0005
R1460 GND.n328 GND.n327 45.0005
R1461 GND.n639 GND.n329 45.0005
R1462 GND.n700 GND.n329 45.0005
R1463 GND.n715 GND.n714 45.0005
R1464 GND.n1044 GND.n1043 45.0005
R1465 GND.n1043 GND.n1042 45.0005
R1466 GND.n698 GND.n325 45.0005
R1467 GND.n697 GND.n696 45.0005
R1468 GND.n637 GND.n633 45.0005
R1469 GND.n641 GND.n631 45.0005
R1470 GND.n698 GND.n631 45.0005
R1471 GND.n643 GND.n632 45.0005
R1472 GND.n697 GND.n632 45.0005
R1473 GND.n638 GND.n637 45.0005
R1474 GND.n104 GND.t492 44.7381
R1475 GND.n102 GND.t491 44.7381
R1476 GND.t37 GND.n1134 44.709
R1477 GND.t217 GND.t407 44.6706
R1478 GND.t529 GND.t612 44.6706
R1479 GND.n1001 GND.t309 44.5993
R1480 GND.t0 GND.t24 44.1861
R1481 GND.n691 GND.n690 43.9358
R1482 GND.t29 GND.t64 43.9247
R1483 GND.t30 GND.t59 43.9247
R1484 GND.n522 GND.n517 43.7886
R1485 GND.n716 GND.n715 43.7516
R1486 GND.n902 GND.t544 42.9475
R1487 GND.t623 GND.t41 42.8789
R1488 GND.n933 GND.n932 41.7862
R1489 GND.n934 GND.n933 41.7862
R1490 GND.n483 GND.n421 41.7076
R1491 GND.n499 GND.n411 39.8486
R1492 GND.n480 GND.n470 39.8486
R1493 GND.n449 GND.n434 39.8486
R1494 GND.n1080 GND.t163 39.7414
R1495 GND.n1127 GND.t236 39.7414
R1496 GND.t581 GND.n1101 39.7414
R1497 GND.n374 GND.t365 39.3159
R1498 GND.n366 GND.t364 39.3159
R1499 GND.n365 GND.t316 39.3159
R1500 GND.n370 GND.t315 39.3159
R1501 GND.n372 GND.t258 39.3159
R1502 GND.n373 GND.t259 39.3159
R1503 GND.n377 GND.t166 39.3159
R1504 GND.n376 GND.t167 39.3159
R1505 GND.n144 GND.t425 39.3159
R1506 GND.n1096 GND.t349 39.3159
R1507 GND.n145 GND.t483 39.3159
R1508 GND.n395 GND.t482 39.3159
R1509 GND.n396 GND.t617 39.3159
R1510 GND.n397 GND.t616 39.3159
R1511 GND.n398 GND.t369 39.3159
R1512 GND.n399 GND.t368 39.3159
R1513 GND.n400 GND.t636 39.3159
R1514 GND.n393 GND.t635 39.3159
R1515 GND.n392 GND.t462 39.3159
R1516 GND.n391 GND.t461 39.3159
R1517 GND.n390 GND.t344 39.3159
R1518 GND.n389 GND.t343 39.3159
R1519 GND.n387 GND.t444 39.3159
R1520 GND.n385 GND.t445 39.3159
R1521 GND.n384 GND.t164 39.3159
R1522 GND.n155 GND.t165 39.3159
R1523 GND.n154 GND.t442 39.3159
R1524 GND.n1094 GND.t443 39.3159
R1525 GND.n1095 GND.t211 39.3159
R1526 GND.n1099 GND.t212 39.3159
R1527 GND.n1098 GND.t348 39.3159
R1528 GND.n1115 GND.t426 39.3159
R1529 GND.n120 GND.t557 39.3159
R1530 GND.n119 GND.t556 39.3159
R1531 GND.n118 GND.t267 39.3159
R1532 GND.n117 GND.t266 39.3159
R1533 GND.n116 GND.t434 39.3159
R1534 GND.n115 GND.t433 39.3159
R1535 GND.n114 GND.t115 39.3159
R1536 GND.n113 GND.t114 39.3159
R1537 GND.n111 GND.t363 39.3159
R1538 GND.n110 GND.t362 39.3159
R1539 GND.n109 GND.t400 39.3159
R1540 GND.n108 GND.t399 39.3159
R1541 GND.n107 GND.t420 39.3159
R1542 GND.n106 GND.t419 39.3159
R1543 GND.n1163 GND.t253 39.3159
R1544 GND.n1162 GND.t254 39.3159
R1545 GND.n1161 GND.t241 39.3159
R1546 GND.n1160 GND.t242 39.3159
R1547 GND.n1159 GND.t354 39.3159
R1548 GND.n1158 GND.t355 39.3159
R1549 GND.n1157 GND.t630 39.3159
R1550 GND.n1156 GND.t631 39.3159
R1551 GND.n1150 GND.t134 39.3159
R1552 GND.n1149 GND.t135 39.3159
R1553 GND.n1148 GND.t54 39.3159
R1554 GND.n1147 GND.t55 39.3159
R1555 GND.n1146 GND.t393 39.3159
R1556 GND.n1145 GND.t394 39.3159
R1557 GND.n1144 GND.t12 39.3159
R1558 GND.n1143 GND.t13 39.3159
R1559 GND.n963 GND.t436 39.3159
R1560 GND.n962 GND.t145 39.3159
R1561 GND.n96 GND.t146 39.3159
R1562 GND.n97 GND.t381 39.3159
R1563 GND.n241 GND.t380 39.3159
R1564 GND.n242 GND.t110 39.3159
R1565 GND.n243 GND.t109 39.3159
R1566 GND.n244 GND.t441 39.3159
R1567 GND.n245 GND.t440 39.3159
R1568 GND.n246 GND.t509 39.3159
R1569 GND.n249 GND.t508 39.3159
R1570 GND.n250 GND.t588 39.3159
R1571 GND.n251 GND.t587 39.3159
R1572 GND.n252 GND.t598 39.3159
R1573 GND.n253 GND.t597 39.3159
R1574 GND.n254 GND.t281 39.3159
R1575 GND.n255 GND.t280 39.3159
R1576 GND.n256 GND.t586 39.3159
R1577 GND.n257 GND.t585 39.3159
R1578 GND.n949 GND.t601 39.3159
R1579 GND.n950 GND.t602 39.3159
R1580 GND.n951 GND.t189 39.3159
R1581 GND.n952 GND.t190 39.3159
R1582 GND.n953 GND.t57 39.3159
R1583 GND.n954 GND.t58 39.3159
R1584 GND.n955 GND.t620 39.3159
R1585 GND.n956 GND.t621 39.3159
R1586 GND.n957 GND.t322 39.3159
R1587 GND.n959 GND.t323 39.3159
R1588 GND.n960 GND.t182 39.3159
R1589 GND.n961 GND.t183 39.3159
R1590 GND.n964 GND.t435 39.3159
R1591 GND.n1004 GND.n218 39.0005
R1592 GND.n1004 GND.n1003 39.0005
R1593 GND.t251 GND.t21 38.4342
R1594 GND.n1104 GND.t278 38.4342
R1595 GND.t31 GND.n1103 38.4342
R1596 GND.n378 GND.n377 38.2036
R1597 GND.t339 GND.n945 37.5791
R1598 GND.t32 GND.t96 36.604
R1599 GND.t27 GND.t312 36.604
R1600 GND.n1008 GND.n1007 36.563
R1601 GND.n1007 GND.n163 36.563
R1602 GND GND.t6 36.2742
R1603 GND.t68 GND 36.2742
R1604 GND GND.t432 36.2742
R1605 GND.n275 GND.n273 36.1417
R1606 GND.n276 GND.n275 36.1417
R1607 GND.n284 GND.n282 36.1417
R1608 GND.n285 GND.n284 36.1417
R1609 GND.n293 GND.n291 36.1417
R1610 GND.n294 GND.n293 36.1417
R1611 GND.n267 GND.n266 36.1417
R1612 GND.n943 GND.n266 36.1417
R1613 GND.n894 GND.n720 36.1417
R1614 GND.n890 GND.n720 36.1417
R1615 GND.n890 GND.n889 36.1417
R1616 GND.n889 GND.n888 36.1417
R1617 GND.n888 GND.n730 36.1417
R1618 GND.n882 GND.n881 36.1417
R1619 GND.n881 GND.n880 36.1417
R1620 GND.n880 GND.n741 36.1417
R1621 GND.n874 GND.n741 36.1417
R1622 GND.n874 GND.n873 36.1417
R1623 GND.n868 GND.n752 36.1417
R1624 GND.n862 GND.n752 36.1417
R1625 GND.n862 GND.n861 36.1417
R1626 GND.n861 GND.n860 36.1417
R1627 GND.n860 GND.n762 36.1417
R1628 GND.n854 GND.n853 36.1417
R1629 GND.n853 GND.n852 36.1417
R1630 GND.n852 GND.n773 36.1417
R1631 GND.n846 GND.n773 36.1417
R1632 GND.n846 GND.n845 36.1417
R1633 GND.n840 GND.n784 36.1417
R1634 GND.n834 GND.n784 36.1417
R1635 GND.n834 GND.n833 36.1417
R1636 GND.n833 GND.n832 36.1417
R1637 GND.n832 GND.n794 36.1417
R1638 GND.n826 GND.n825 36.1417
R1639 GND.n825 GND.n824 36.1417
R1640 GND.n824 GND.n805 36.1417
R1641 GND.n818 GND.n805 36.1417
R1642 GND.n818 GND.n817 36.1417
R1643 GND.n1266 GND.n1265 36.1417
R1644 GND.n1265 GND.n1264 36.1417
R1645 GND.n1264 GND.n42 36.1417
R1646 GND.n1258 GND.n42 36.1417
R1647 GND.n1258 GND.n1257 36.1417
R1648 GND.n1252 GND.n53 36.1417
R1649 GND.n1246 GND.n53 36.1417
R1650 GND.n1241 GND.n58 36.1417
R1651 GND.n1204 GND.n58 36.1417
R1652 GND.n1233 GND.n1232 36.1417
R1653 GND.n1232 GND.n1231 36.1417
R1654 GND.n1226 GND.n1214 36.1417
R1655 GND.n1219 GND.n1214 36.1417
R1656 GND.n900 GND.t63 36.1338
R1657 GND.t610 GND.t124 36.1338
R1658 GND.t489 GND.t122 35.8196
R1659 GND.t27 GND.t96 35.5582
R1660 GND.t312 GND.t29 35.5582
R1661 GND.n104 GND.t371 35.1381
R1662 GND.n102 GND.t370 35.1381
R1663 GND.n1277 GND.n29 34.6358
R1664 GND.n1281 GND.n1280 34.6358
R1665 GND.n1283 GND.n1281 34.6358
R1666 GND.n1317 GND.n1316 34.6358
R1667 GND.n1363 GND.n1360 34.6358
R1668 GND.n690 GND.n646 34.6358
R1669 GND.n686 GND.n646 34.6358
R1670 GND.n686 GND.n685 34.6358
R1671 GND.n685 GND.n684 34.6358
R1672 GND.n684 GND.n648 34.6358
R1673 GND.n679 GND.n649 34.6358
R1674 GND.n675 GND.n674 34.6358
R1675 GND.n674 GND.n651 34.6358
R1676 GND.n670 GND.n651 34.6358
R1677 GND.n667 GND.n655 34.6358
R1678 GND.n662 GND.n656 34.6358
R1679 GND.n436 GND.n415 34.6358
R1680 GND.n507 GND.n506 34.6358
R1681 GND.n497 GND.n413 34.6358
R1682 GND.n504 GND.n409 34.6358
R1683 GND.n451 GND.n431 34.6358
R1684 GND.n478 GND.n472 34.6358
R1685 GND.n468 GND.n467 34.6358
R1686 GND.n462 GND.n461 34.6358
R1687 GND.n445 GND.n443 34.6358
R1688 GND.t271 GND.t61 33.8625
R1689 GND.t21 GND.t566 33.728
R1690 GND.n1104 GND.t510 33.728
R1691 GND.n1103 GND.t42 33.728
R1692 GND.t50 GND.t599 33.717
R1693 GND.n476 GND.n473 33.5688
R1694 GND.n440 GND.n437 33.5688
R1695 GND.n495 GND.n414 33.5688
R1696 GND.n407 GND.n406 33.5688
R1697 GND.n464 GND.n426 33.5688
R1698 GND.n453 GND.n432 33.5688
R1699 GND.n1363 GND.n1362 32.7534
R1700 GND.n1022 GND.t118 32.6237
R1701 GND.n1006 GND.n217 32.5005
R1702 GND.n1006 GND.n1005 32.5005
R1703 GND.n422 GND.n420 30.79
R1704 GND.n420 GND.n419 30.79
R1705 GND.n485 GND.n484 30.79
R1706 GND.n486 GND.n485 30.79
R1707 GND.n428 GND.n421 30.79
R1708 GND.n1024 GND.n1023 30.79
R1709 GND.n1023 GND.n1022 30.79
R1710 GND.t608 GND.t209 29.9395
R1711 GND.n1178 GND.n1177 29.3652
R1712 GND.t22 GND.t623 29.2833
R1713 GND.t41 GND.t581 29.2833
R1714 GND GND.t1 29.0195
R1715 GND.t480 GND 29.0195
R1716 GND.t618 GND 29.0195
R1717 GND.n1190 GND.n1189 28.9887
R1718 GND.n1062 GND.n75 28.9887
R1719 GND.t544 GND.n901 28.4942
R1720 GND.n1194 GND.t314 28.4942
R1721 GND.t64 GND.t30 28.2375
R1722 GND.t59 GND.t26 28.2375
R1723 GND.n1134 GND.t26 27.4531
R1724 GND.t222 GND.n698 26.6966
R1725 GND.n698 GND.t341 26.6966
R1726 GND.t18 GND.n697 26.6966
R1727 GND.n697 GND.t456 26.6966
R1728 GND.n637 GND.t387 26.6966
R1729 GND.n637 GND.t178 26.6966
R1730 GND.n193 GND.n192 26.5914
R1731 GND.t256 GND.n193 26.5914
R1732 GND.t430 GND.t308 26.2229
R1733 GND.t8 GND.t460 26.1458
R1734 GND.n1316 GND.n1315 25.977
R1735 GND.n680 GND.n648 25.977
R1736 GND.n670 GND.n669 25.977
R1737 GND.n1050 GND.n1049 25.4353
R1738 GND.n1051 GND.n1050 25.4353
R1739 GND.n1135 GND.t35 25.3615
R1740 GND.n530 GND.n361 25.224
R1741 GND.n534 GND.n361 25.224
R1742 GND.n536 GND.n535 25.224
R1743 GND.n536 GND.n358 25.224
R1744 GND.n541 GND.n357 25.224
R1745 GND.n545 GND.n357 25.224
R1746 GND.n547 GND.n546 25.224
R1747 GND.n547 GND.n354 25.224
R1748 GND.n552 GND.n353 25.224
R1749 GND.n556 GND.n353 25.224
R1750 GND.n558 GND.n557 25.224
R1751 GND.n558 GND.n350 25.224
R1752 GND.n563 GND.n349 25.224
R1753 GND.n567 GND.n349 25.224
R1754 GND.n569 GND.n568 25.224
R1755 GND.n569 GND.n346 25.224
R1756 GND.n574 GND.n345 25.224
R1757 GND.n578 GND.n345 25.224
R1758 GND.n580 GND.n579 25.224
R1759 GND.n580 GND.n342 25.224
R1760 GND.n585 GND.n341 25.224
R1761 GND.n589 GND.n341 25.224
R1762 GND.n591 GND.n590 25.224
R1763 GND.n591 GND.n338 25.224
R1764 GND.n596 GND.n337 25.224
R1765 GND.n600 GND.n337 25.224
R1766 GND.n602 GND.n601 25.224
R1767 GND.n602 GND.n334 25.224
R1768 GND.n607 GND.n333 25.224
R1769 GND.n611 GND.n333 25.224
R1770 GND.n613 GND.n612 25.224
R1771 GND.n613 GND.n330 25.224
R1772 GND.n624 GND.n331 25.224
R1773 GND.n624 GND.n623 25.224
R1774 GND.n622 GND.n621 25.224
R1775 GND.n621 GND.n618 25.224
R1776 GND.n1387 GND.n1386 25.224
R1777 GND.n1386 GND.n1385 25.224
R1778 GND.n1384 GND.n1383 25.224
R1779 GND.n1383 GND.n5 25.224
R1780 GND.n694 GND.n645 25.1797
R1781 GND.n695 GND.n634 25.1797
R1782 GND.n636 GND.n635 25.1797
R1783 GND.n702 GND.n324 25.1797
R1784 GND.n703 GND.n322 25.1797
R1785 GND.n704 GND.n314 25.1797
R1786 GND.n316 GND.n315 25.1797
R1787 GND.n710 GND.n307 25.1797
R1788 GND.n306 GND.n305 25.1797
R1789 GND.n520 GND.n519 25.1797
R1790 GND.n521 GND.n518 25.1797
R1791 GND.n1127 GND.t624 25.1
R1792 GND.n417 GND.t505 25.0567
R1793 GND.n1353 GND.n1352 24.4711
R1794 GND.n1352 GND.n1351 24.4711
R1795 GND.n1330 GND.n1329 24.4711
R1796 GND.t609 GND.t120 24.3646
R1797 GND.n1317 GND.n1272 24.0946
R1798 GND.n680 GND.n679 24.0946
R1799 GND.n1302 GND.n1292 23.7181
R1800 GND.n1304 GND.n1289 23.7181
R1801 GND.n1324 GND.n29 23.7181
R1802 GND.n1321 GND.n1273 23.7181
R1803 GND.n1360 GND.n1359 23.7181
R1804 GND.n1368 GND.n14 23.7181
R1805 GND.n1358 GND.n17 23.7181
R1806 GND.n1348 GND.n1347 23.7181
R1807 GND.n1339 GND.n1338 23.7181
R1808 GND.n668 GND.n667 23.7181
R1809 GND.n663 GND.n662 23.7181
R1810 GND.n488 GND.n415 23.7181
R1811 GND.n507 GND.n404 23.7181
R1812 GND.n498 GND.n497 23.7181
R1813 GND.n505 GND.n504 23.7181
R1814 GND.n451 GND.n450 23.7181
R1815 GND.n479 GND.n478 23.7181
R1816 GND.n467 GND.n425 23.7181
R1817 GND.n461 GND.n460 23.7181
R1818 GND.n443 GND.n442 23.7181
R1819 GND.n1332 GND.n24 23.3417
R1820 GND.t464 GND.n905 23.1258
R1821 GND.t605 GND.n60 22.7128
R1822 GND.n1041 GND.t337 22.5064
R1823 GND.n1298 GND.n1292 22.2123
R1824 GND.n1304 GND.n1303 22.2123
R1825 GND.n1359 GND.n1358 22.2123
R1826 GND.n1343 GND.n1342 22.2123
R1827 GND.n663 GND.n655 22.2123
R1828 GND.n658 GND.n656 22.2123
R1829 GND.n442 GND.n436 22.2123
R1830 GND.n506 GND.n505 22.2123
R1831 GND.n492 GND.n413 22.2123
R1832 GND.n499 GND.n498 22.2123
R1833 GND.n410 GND.n409 22.2123
R1834 GND.n456 GND.n431 22.2123
R1835 GND.n472 GND.n364 22.2123
R1836 GND.n480 GND.n479 22.2123
R1837 GND.n469 GND.n468 22.2123
R1838 GND.n462 GND.n425 22.2123
R1839 GND.n450 GND.n449 22.2123
R1840 GND.n445 GND.n444 22.2123
R1841 GND.t512 GND.t437 21.9626
R1842 GND.t510 GND.t470 21.9626
R1843 GND.t42 GND.t553 21.9626
R1844 GND.t24 GND.t75 21.9626
R1845 GND.t122 GND.t143 21.7011
R1846 GND.n422 GND 21.0039
R1847 GND.t604 GND.n900 20.8546
R1848 GND.t606 GND.t464 20.8546
R1849 GND.t126 GND.t543 20.8546
R1850 GND.t124 GND.t513 20.8546
R1851 GND.t61 GND.t125 20.8546
R1852 GND.n488 GND 20.7453
R1853 GND GND.n404 20.7453
R1854 GND.n491 GND 20.7453
R1855 GND.n457 GND 20.7453
R1856 GND.n460 GND 20.7453
R1857 GND GND.n514 20.7453
R1858 GND.n535 GND.n534 20.3299
R1859 GND.n546 GND.n545 20.3299
R1860 GND.n557 GND.n556 20.3299
R1861 GND.n568 GND.n567 20.3299
R1862 GND.n579 GND.n578 20.3299
R1863 GND.n590 GND.n589 20.3299
R1864 GND.n601 GND.n600 20.3299
R1865 GND.n612 GND.n611 20.3299
R1866 GND.n623 GND.n622 20.3299
R1867 GND.n1385 GND.n1384 20.3299
R1868 GND.n1354 GND.n1353 19.9534
R1869 GND.n1077 GND.n163 19.8222
R1870 GND.n934 GND.t60 19.4092
R1871 GND.t463 GND.n918 19.2028
R1872 GND.n1331 GND.n1330 19.2005
R1873 GND.n1068 GND.n1067 18.2817
R1874 GND.n1067 GND.n1066 18.2817
R1875 GND.n1065 GND.n1064 18.2817
R1876 GND.n1066 GND.n1065 18.2817
R1877 GND.n993 GND.n992 18.2817
R1878 GND.n994 GND.n993 18.2817
R1879 GND.n996 GND.n995 18.2817
R1880 GND.n995 GND.n994 18.2817
R1881 GND.n987 GND.n986 18.2817
R1882 GND.n986 GND.n985 18.2817
R1883 GND.n968 GND.n967 18.2817
R1884 GND.n985 GND.n968 18.2817
R1885 GND.n1176 GND.n1175 18.2817
R1886 GND.n1175 GND.n1174 18.2817
R1887 GND.n1173 GND.n1172 18.2817
R1888 GND.n1174 GND.n1173 18.2817
R1889 GND.n1188 GND.n1187 18.2817
R1890 GND.n1187 GND.n1186 18.2817
R1891 GND.n86 GND.n80 18.2817
R1892 GND.n87 GND.n80 18.2817
R1893 GND.n231 GND.n78 18.2817
R1894 GND.n1186 GND.n78 18.2817
R1895 GND.n1180 GND.n81 18.2817
R1896 GND.n87 GND.n81 18.2817
R1897 GND.n220 GND.n219 18.2817
R1898 GND.n917 GND.n220 18.2817
R1899 GND.n223 GND.n221 18.2817
R1900 GND.n917 GND.n221 18.2817
R1901 GND.n63 GND.n61 18.2817
R1902 GND.n901 GND.n61 18.2817
R1903 GND.n1199 GND.n62 18.2817
R1904 GND.n901 GND.n62 18.2817
R1905 GND.n1193 GND.n1192 18.2817
R1906 GND.n1194 GND.n1193 18.2817
R1907 GND.n1196 GND.n1195 18.2817
R1908 GND.n1195 GND.n1194 18.2817
R1909 GND.n1054 GND.n1053 18.2817
R1910 GND.n1053 GND.n1052 18.2817
R1911 GND.n184 GND.n183 18.2817
R1912 GND.n1052 GND.n184 18.2817
R1913 GND.t201 GND.t607 18.1704
R1914 GND.n530 GND.n529 17.3181
R1915 GND.n541 GND.n540 17.3181
R1916 GND.n552 GND.n551 17.3181
R1917 GND.n563 GND.n562 17.3181
R1918 GND.n574 GND.n573 17.3181
R1919 GND.n585 GND.n584 17.3181
R1920 GND.n596 GND.n595 17.3181
R1921 GND.n607 GND.n606 17.3181
R1922 GND.n628 GND.n331 17.3181
R1923 GND.n1387 GND.n2 17.3181
R1924 GND.t278 GND.t34 17.2564
R1925 GND.t511 GND.t25 17.2564
R1926 GND.t277 GND.t31 17.2564
R1927 GND.t28 GND.t324 17.2564
R1928 GND.n137 GND.n127 17.2064
R1929 GND.n1101 GND.n127 17.2064
R1930 GND.n1131 GND.n128 17.2064
R1931 GND.n1101 GND.n128 17.2064
R1932 GND.n924 GND.n923 17.2064
R1933 GND.n923 GND.t271 17.2064
R1934 GND.n1081 GND.n1080 15.9492
R1935 GND.n540 GND.n358 15.8123
R1936 GND.n551 GND.n354 15.8123
R1937 GND.n562 GND.n350 15.8123
R1938 GND.n573 GND.n346 15.8123
R1939 GND.n584 GND.n342 15.8123
R1940 GND.n595 GND.n338 15.8123
R1941 GND.n606 GND.n334 15.8123
R1942 GND.n628 GND.n330 15.8123
R1943 GND.n618 GND.n2 15.8123
R1944 GND.n226 GND.t98 15.4862
R1945 GND.n1315 GND.n1287 15.4358
R1946 GND.n1333 GND.n1331 15.4358
R1947 GND.n112 GND.n111 15.0979
R1948 GND.n213 GND.n211 15.0005
R1949 GND.t120 GND.n211 15.0005
R1950 GND.t247 GND.n699 14.708
R1951 GND.t62 GND.t287 14.6603
R1952 GND.t647 GND.t624 14.6419
R1953 GND.t645 GND.t469 14.6419
R1954 GND.t143 GND.t625 14.6419
R1955 GND.t646 GND.t489 14.6419
R1956 GND.t144 GND.t468 14.6419
R1957 GND.t7 GND.t361 14.51
R1958 GND.t614 GND.t634 14.51
R1959 GND.t20 GND.t67 14.51
R1960 GND.t497 GND.t430 14.2473
R1961 GND.t545 GND.n902 14.0409
R1962 GND.t209 GND.n908 14.0409
R1963 GND.t311 GND.t498 14.0409
R1964 GND.t498 GND.n163 13.8344
R1965 GND.n1156 GND.n1155 13.7851
R1966 GND.n1329 GND.n1328 13.5534
R1967 GND.n1114 GND.n1113 13.296
R1968 GND.n1113 GND.n125 13.296
R1969 GND.n375 GND.n368 13.296
R1970 GND.n380 GND.n368 13.296
R1971 GND.n371 GND.n367 13.296
R1972 GND.n369 GND.n367 13.296
R1973 GND.n388 GND.n147 13.296
R1974 GND.n1076 GND.n147 13.296
R1975 GND.n1169 GND.n1168 13.296
R1976 GND.n1168 GND.n1167 13.296
R1977 GND.n1142 GND.n1141 13.296
R1978 GND.n1141 GND.n1140 13.296
R1979 GND.n1165 GND.n1164 13.296
R1980 GND.n1166 GND.n1165 13.296
R1981 GND.n948 GND.n947 13.296
R1982 GND.n947 GND.n946 13.296
R1983 GND.n917 GND.t256 13.215
R1984 GND.n1311 GND.n1287 13.177
R1985 GND.n1354 GND.n17 13.177
R1986 GND.n669 GND.n668 13.177
R1987 GND.n512 GND.n511 13.0995
R1988 GND.n510 GND.n509 13.0995
R1989 GND.n1003 GND.t62 12.802
R1990 GND.n1297 GND.n1293 12.8005
R1991 GND.n1308 GND.n1288 12.8005
R1992 GND.n1343 GND.n21 12.8005
R1993 GND.n1337 GND.n24 12.8005
R1994 GND.n1374 GND.n10 12.8005
R1995 GND.n658 GND.n10 12.8005
R1996 GND.n492 GND.n491 12.8005
R1997 GND.n457 GND.n456 12.8005
R1998 GND.n514 GND.n364 12.8005
R1999 GND.n1040 GND.n1039 12.4473
R2000 GND.n1041 GND.n1040 12.4473
R2001 GND.n922 GND.t609 12.389
R2002 GND.n1069 GND.n1068 12.0476
R2003 GND.n1151 GND.t87 11.8635
R2004 GND.n946 GND.t605 11.3567
R2005 GND.n1298 GND.n1297 11.2946
R2006 GND.n1303 GND.n1302 11.2946
R2007 GND.n1308 GND.n1289 11.2946
R2008 GND.n1311 GND.n1288 11.2946
R2009 GND.n1347 GND.n21 11.2946
R2010 GND.n1338 GND.n1337 11.2946
R2011 GND.n1039 GND.n1038 11.2946
R2012 GND.n1049 GND.n1048 11.2946
R2013 GND.n1025 GND.n1024 11.2946
R2014 GND.n484 GND.n423 10.9181
R2015 GND.t306 GND.t288 10.7372
R2016 GND.n1277 GND.n1275 10.5417
R2017 GND.n1283 GND.n1282 10.5417
R2018 GND.n1348 GND.n20 10.5417
R2019 GND.n1339 GND.n22 10.5417
R2020 GND.n650 GND.n649 10.5417
R2021 GND.n934 GND.t126 10.5308
R2022 GND.n1031 GND.t309 10.5308
R2023 GND.n901 GND.t201 10.3243
R2024 GND.n1003 GND.n1002 10.3243
R2025 GND.n249 GND.n248 10.1749
R2026 GND GND.n423 10.0862
R2027 GND.n483 GND 10.0862
R2028 GND.n1073 GND.n1072 9.91575
R2029 GND.n1074 GND.n1073 9.91575
R2030 GND.n172 GND.n168 9.91575
R2031 GND.n1074 GND.n168 9.91575
R2032 GND.n273 GND.n272 9.32838
R2033 GND.n509 GND.n404 9.3031
R2034 GND.n940 GND.n939 9.3005
R2035 GND.n506 GND.n405 9.3005
R2036 GND.n508 GND.n507 9.3005
R2037 GND.n505 GND.n408 9.3005
R2038 GND.n502 GND.n409 9.3005
R2039 GND.n504 GND.n503 9.3005
R2040 GND.n489 GND.n488 9.3005
R2041 GND.n439 GND.n436 9.3005
R2042 GND.n438 GND.n415 9.3005
R2043 GND.n498 GND.n412 9.3005
R2044 GND.n493 GND.n492 9.3005
R2045 GND.n491 GND.n490 9.3005
R2046 GND.n494 GND.n413 9.3005
R2047 GND.n497 GND.n496 9.3005
R2048 GND.n500 GND.n499 9.3005
R2049 GND.n442 GND.n441 9.3005
R2050 GND.n460 GND.n459 9.3005
R2051 GND.n465 GND.n425 9.3005
R2052 GND.n468 GND.n424 9.3005
R2053 GND.n467 GND.n466 9.3005
R2054 GND.n463 GND.n462 9.3005
R2055 GND.n461 GND.n427 9.3005
R2056 GND.n456 GND.n455 9.3005
R2057 GND.n458 GND.n457 9.3005
R2058 GND.n454 GND.n431 9.3005
R2059 GND.n452 GND.n451 9.3005
R2060 GND.n450 GND.n433 9.3005
R2061 GND.n449 GND.n448 9.3005
R2062 GND.n446 GND.n445 9.3005
R2063 GND.n443 GND.n435 9.3005
R2064 GND.n479 GND.n471 9.3005
R2065 GND.n474 GND.n364 9.3005
R2066 GND.n475 GND.n472 9.3005
R2067 GND.n478 GND.n477 9.3005
R2068 GND.n481 GND.n480 9.3005
R2069 GND.n514 GND.n513 9.3005
R2070 GND.n297 GND.n296 9.3005
R2071 GND.n298 GND.n297 9.3005
R2072 GND.n288 GND.n287 9.3005
R2073 GND.n289 GND.n288 9.3005
R2074 GND.n279 GND.n278 9.3005
R2075 GND.n280 GND.n279 9.3005
R2076 GND.n943 GND.n942 9.3005
R2077 GND.n299 GND.n266 9.3005
R2078 GND.n268 GND.n267 9.3005
R2079 GND.n295 GND.n294 9.3005
R2080 GND.n293 GND.n269 9.3005
R2081 GND.n291 GND.n290 9.3005
R2082 GND.n286 GND.n285 9.3005
R2083 GND.n284 GND.n270 9.3005
R2084 GND.n282 GND.n281 9.3005
R2085 GND.n277 GND.n276 9.3005
R2086 GND.n275 GND.n271 9.3005
R2087 GND.n1216 GND.n1215 9.3005
R2088 GND.n1217 GND.n1216 9.3005
R2089 GND.n1228 GND.n1212 9.3005
R2090 GND.n1229 GND.n1228 9.3005
R2091 GND.n1207 GND.n1206 9.3005
R2092 GND.n1208 GND.n1207 9.3005
R2093 GND.n1243 GND.n56 9.3005
R2094 GND.n1244 GND.n1243 9.3005
R2095 GND.n1254 GND.n51 9.3005
R2096 GND.n1255 GND.n1254 9.3005
R2097 GND.n47 GND.n46 9.3005
R2098 GND.n48 GND.n47 9.3005
R2099 GND.n814 GND.n813 9.3005
R2100 GND.n815 GND.n814 9.3005
R2101 GND.n809 GND.n808 9.3005
R2102 GND.n810 GND.n809 9.3005
R2103 GND.n800 GND.n799 9.3005
R2104 GND.n801 GND.n800 9.3005
R2105 GND.n790 GND.n789 9.3005
R2106 GND.n791 GND.n790 9.3005
R2107 GND.n842 GND.n782 9.3005
R2108 GND.n843 GND.n842 9.3005
R2109 GND.n778 GND.n777 9.3005
R2110 GND.n779 GND.n778 9.3005
R2111 GND.n768 GND.n767 9.3005
R2112 GND.n769 GND.n768 9.3005
R2113 GND.n758 GND.n757 9.3005
R2114 GND.n759 GND.n758 9.3005
R2115 GND.n870 GND.n750 9.3005
R2116 GND.n871 GND.n870 9.3005
R2117 GND.n746 GND.n745 9.3005
R2118 GND.n747 GND.n746 9.3005
R2119 GND.n736 GND.n735 9.3005
R2120 GND.n737 GND.n736 9.3005
R2121 GND.n726 GND.n725 9.3005
R2122 GND.n727 GND.n726 9.3005
R2123 GND.n1219 GND.n1218 9.3005
R2124 GND.n1214 GND.n1213 9.3005
R2125 GND.n1227 GND.n1226 9.3005
R2126 GND.n1231 GND.n1230 9.3005
R2127 GND.n1232 GND.n1210 9.3005
R2128 GND.n1233 GND.n1209 9.3005
R2129 GND.n1205 GND.n1204 9.3005
R2130 GND.n58 GND.n57 9.3005
R2131 GND.n1242 GND.n1241 9.3005
R2132 GND.n1246 GND.n1245 9.3005
R2133 GND.n53 GND.n52 9.3005
R2134 GND.n1253 GND.n1252 9.3005
R2135 GND.n1257 GND.n1256 9.3005
R2136 GND.n1258 GND.n50 9.3005
R2137 GND.n49 GND.n42 9.3005
R2138 GND.n1264 GND.n41 9.3005
R2139 GND.n1265 GND.n40 9.3005
R2140 GND.n1266 GND.n39 9.3005
R2141 GND.n817 GND.n816 9.3005
R2142 GND.n818 GND.n812 9.3005
R2143 GND.n811 GND.n805 9.3005
R2144 GND.n824 GND.n804 9.3005
R2145 GND.n825 GND.n803 9.3005
R2146 GND.n826 GND.n802 9.3005
R2147 GND.n798 GND.n794 9.3005
R2148 GND.n832 GND.n793 9.3005
R2149 GND.n833 GND.n792 9.3005
R2150 GND.n834 GND.n788 9.3005
R2151 GND.n784 GND.n783 9.3005
R2152 GND.n841 GND.n840 9.3005
R2153 GND.n845 GND.n844 9.3005
R2154 GND.n846 GND.n781 9.3005
R2155 GND.n780 GND.n773 9.3005
R2156 GND.n852 GND.n772 9.3005
R2157 GND.n853 GND.n771 9.3005
R2158 GND.n854 GND.n770 9.3005
R2159 GND.n766 GND.n762 9.3005
R2160 GND.n860 GND.n761 9.3005
R2161 GND.n861 GND.n760 9.3005
R2162 GND.n862 GND.n756 9.3005
R2163 GND.n752 GND.n751 9.3005
R2164 GND.n869 GND.n868 9.3005
R2165 GND.n873 GND.n872 9.3005
R2166 GND.n874 GND.n749 9.3005
R2167 GND.n748 GND.n741 9.3005
R2168 GND.n880 GND.n740 9.3005
R2169 GND.n881 GND.n739 9.3005
R2170 GND.n882 GND.n738 9.3005
R2171 GND.n734 GND.n730 9.3005
R2172 GND.n888 GND.n729 9.3005
R2173 GND.n889 GND.n728 9.3005
R2174 GND.n890 GND.n724 9.3005
R2175 GND.n720 GND.n719 9.3005
R2176 GND.n895 GND.n894 9.3005
R2177 GND.n657 GND.n10 9.3005
R2178 GND.n659 GND.n658 9.3005
R2179 GND.n660 GND.n656 9.3005
R2180 GND.n662 GND.n661 9.3005
R2181 GND.n664 GND.n663 9.3005
R2182 GND.n665 GND.n655 9.3005
R2183 GND.n667 GND.n666 9.3005
R2184 GND.n668 GND.n653 9.3005
R2185 GND.n669 GND.n652 9.3005
R2186 GND.n671 GND.n670 9.3005
R2187 GND.n672 GND.n651 9.3005
R2188 GND.n674 GND.n673 9.3005
R2189 GND.n676 GND.n675 9.3005
R2190 GND.n677 GND.n649 9.3005
R2191 GND.n679 GND.n678 9.3005
R2192 GND.n681 GND.n680 9.3005
R2193 GND.n682 GND.n648 9.3005
R2194 GND.n684 GND.n683 9.3005
R2195 GND.n685 GND.n647 9.3005
R2196 GND.n687 GND.n686 9.3005
R2197 GND.n688 GND.n646 9.3005
R2198 GND.n690 GND.n689 9.3005
R2199 GND.n1375 GND.n1374 9.3005
R2200 GND.n1328 GND.n1327 9.3005
R2201 GND.n1335 GND.n24 9.3005
R2202 GND.n1337 GND.n1336 9.3005
R2203 GND.n1347 GND.n1346 9.3005
R2204 GND.n1355 GND.n1354 9.3005
R2205 GND.n1356 GND.n17 9.3005
R2206 GND.n1365 GND.n14 9.3005
R2207 GND.n1368 GND.n1367 9.3005
R2208 GND.n1364 GND.n1363 9.3005
R2209 GND.n1360 GND.n15 9.3005
R2210 GND.n1359 GND.n16 9.3005
R2211 GND.n1358 GND.n1357 9.3005
R2212 GND.n1353 GND.n18 9.3005
R2213 GND.n1352 GND.n19 9.3005
R2214 GND.n1351 GND.n1350 9.3005
R2215 GND.n1349 GND.n1348 9.3005
R2216 GND.n1345 GND.n21 9.3005
R2217 GND.n1344 GND.n1343 9.3005
R2218 GND.n1342 GND.n1341 9.3005
R2219 GND.n1340 GND.n1339 9.3005
R2220 GND.n1338 GND.n23 9.3005
R2221 GND.n1334 GND.n1333 9.3005
R2222 GND.n1330 GND.n26 9.3005
R2223 GND.n1329 GND.n27 9.3005
R2224 GND.n1321 GND.n1320 9.3005
R2225 GND.n1315 GND.n1314 9.3005
R2226 GND.n1290 GND.n1288 9.3005
R2227 GND.n1308 GND.n1307 9.3005
R2228 GND.n1303 GND.n1291 9.3005
R2229 GND.n1299 GND.n1298 9.3005
R2230 GND.n1297 GND.n1296 9.3005
R2231 GND.n1295 GND.n1293 9.3005
R2232 GND.n1300 GND.n1292 9.3005
R2233 GND.n1302 GND.n1301 9.3005
R2234 GND.n1305 GND.n1304 9.3005
R2235 GND.n1306 GND.n1289 9.3005
R2236 GND.n1312 GND.n1311 9.3005
R2237 GND.n1313 GND.n1287 9.3005
R2238 GND.n1316 GND.n1286 9.3005
R2239 GND.n1318 GND.n1317 9.3005
R2240 GND.n1319 GND.n1272 9.3005
R2241 GND.n1285 GND.n1273 9.3005
R2242 GND.n1284 GND.n1283 9.3005
R2243 GND.n1281 GND.n1274 9.3005
R2244 GND.n1280 GND.n1279 9.3005
R2245 GND.n1278 GND.n1277 9.3005
R2246 GND.n1276 GND.n29 9.3005
R2247 GND.n1325 GND.n1324 9.3005
R2248 GND.n1381 GND.n5 9.3005
R2249 GND.n1383 GND.n1382 9.3005
R2250 GND.n1384 GND.n4 9.3005
R2251 GND.n1385 GND.n3 9.3005
R2252 GND.n1386 GND.n1 9.3005
R2253 GND.n1388 GND.n1387 9.3005
R2254 GND.n2 GND.n0 9.3005
R2255 GND.n619 GND.n618 9.3005
R2256 GND.n621 GND.n620 9.3005
R2257 GND.n622 GND.n617 9.3005
R2258 GND.n623 GND.n616 9.3005
R2259 GND.n625 GND.n624 9.3005
R2260 GND.n626 GND.n331 9.3005
R2261 GND.n628 GND.n627 9.3005
R2262 GND.n615 GND.n330 9.3005
R2263 GND.n614 GND.n613 9.3005
R2264 GND.n612 GND.n332 9.3005
R2265 GND.n611 GND.n610 9.3005
R2266 GND.n609 GND.n333 9.3005
R2267 GND.n608 GND.n607 9.3005
R2268 GND.n606 GND.n605 9.3005
R2269 GND.n604 GND.n334 9.3005
R2270 GND.n603 GND.n602 9.3005
R2271 GND.n601 GND.n336 9.3005
R2272 GND.n600 GND.n599 9.3005
R2273 GND.n598 GND.n337 9.3005
R2274 GND.n597 GND.n596 9.3005
R2275 GND.n595 GND.n594 9.3005
R2276 GND.n593 GND.n338 9.3005
R2277 GND.n592 GND.n591 9.3005
R2278 GND.n590 GND.n340 9.3005
R2279 GND.n589 GND.n588 9.3005
R2280 GND.n587 GND.n341 9.3005
R2281 GND.n586 GND.n585 9.3005
R2282 GND.n584 GND.n583 9.3005
R2283 GND.n582 GND.n342 9.3005
R2284 GND.n581 GND.n580 9.3005
R2285 GND.n579 GND.n344 9.3005
R2286 GND.n578 GND.n577 9.3005
R2287 GND.n576 GND.n345 9.3005
R2288 GND.n575 GND.n574 9.3005
R2289 GND.n573 GND.n572 9.3005
R2290 GND.n571 GND.n346 9.3005
R2291 GND.n570 GND.n569 9.3005
R2292 GND.n568 GND.n348 9.3005
R2293 GND.n567 GND.n566 9.3005
R2294 GND.n565 GND.n349 9.3005
R2295 GND.n564 GND.n563 9.3005
R2296 GND.n562 GND.n561 9.3005
R2297 GND.n560 GND.n350 9.3005
R2298 GND.n559 GND.n558 9.3005
R2299 GND.n557 GND.n352 9.3005
R2300 GND.n556 GND.n555 9.3005
R2301 GND.n554 GND.n353 9.3005
R2302 GND.n553 GND.n552 9.3005
R2303 GND.n551 GND.n550 9.3005
R2304 GND.n549 GND.n354 9.3005
R2305 GND.n548 GND.n547 9.3005
R2306 GND.n546 GND.n356 9.3005
R2307 GND.n545 GND.n544 9.3005
R2308 GND.n543 GND.n357 9.3005
R2309 GND.n542 GND.n541 9.3005
R2310 GND.n540 GND.n539 9.3005
R2311 GND.n538 GND.n358 9.3005
R2312 GND.n537 GND.n536 9.3005
R2313 GND.n535 GND.n360 9.3005
R2314 GND.n534 GND.n533 9.3005
R2315 GND.n532 GND.n361 9.3005
R2316 GND.n531 GND.n530 9.3005
R2317 GND.n529 GND.n528 9.3005
R2318 GND.n379 GND.n378 9.14112
R2319 GND.n381 GND.n379 9.14112
R2320 GND.n383 GND.n382 9.14112
R2321 GND.n382 GND.n381 9.14112
R2322 GND.n1321 GND.n1272 9.03579
R2323 GND.n958 GND.n957 8.94409
R2324 GND.t56 GND.t119 8.87896
R2325 GND.n473 GND.t265 8.7005
R2326 GND.n473 GND.t519 8.7005
R2327 GND.n437 GND.t80 8.7005
R2328 GND.n437 GND.t481 8.7005
R2329 GND.n414 GND.t94 8.7005
R2330 GND.n414 GND.t291 8.7005
R2331 GND.n406 GND.t422 8.7005
R2332 GND.n406 GND.t2 8.7005
R2333 GND.n426 GND.t148 8.7005
R2334 GND.n426 GND.t619 8.7005
R2335 GND.n432 GND.t274 8.7005
R2336 GND.n432 GND.t151 8.7005
R2337 GND.n1119 GND.n1118 8.47876
R2338 GND.t27 GND.n1119 8.47876
R2339 GND.n1110 GND.n1109 8.47876
R2340 GND.t488 GND.n1110 8.47876
R2341 GND.n1090 GND.n1089 8.47876
R2342 GND.n1089 GND.t567 8.47876
R2343 GND.n1121 GND.n1120 8.47876
R2344 GND.n1120 GND.t27 8.47876
R2345 GND.n1085 GND.n150 8.47876
R2346 GND.t488 GND.n150 8.47876
R2347 GND.n1088 GND.n1087 8.47876
R2348 GND.t567 GND.n1088 8.47876
R2349 GND.t208 GND.n922 8.46601
R2350 GND.n1002 GND.t306 8.46601
R2351 GND.n1021 GND.t98 8.46601
R2352 GND.n1052 GND.t513 7.64011
R2353 GND.t125 GND.n917 7.64011
R2354 GND.t490 GND.t411 7.3212
R2355 GND.t649 GND.t410 7.3212
R2356 GND.t268 GND.t412 7.3212
R2357 GND.t488 GND.t95 7.3212
R2358 GND.t648 GND.t236 7.3212
R2359 GND.n1126 GND.n1125 7.13465
R2360 GND.n1127 GND.n1126 7.13465
R2361 GND.n1129 GND.n1128 7.13465
R2362 GND.n1128 GND.n1127 7.13465
R2363 GND.t120 GND.n921 7.02068
R2364 GND.n905 GND.t545 6.8142
R2365 GND.n1280 GND.n1275 6.77697
R2366 GND.n1282 GND.n1273 6.77697
R2367 GND.n1351 GND.n20 6.77697
R2368 GND.n1342 GND.n22 6.77697
R2369 GND.n675 GND.n650 6.77697
R2370 GND.n1077 GND.n166 6.44556
R2371 GND.n1094 GND.n148 6.31845
R2372 GND.n946 GND.t339 6.19477
R2373 GND.t60 GND.t606 6.19477
R2374 GND.t543 GND.t608 6.19477
R2375 GND.t287 GND.t210 6.19477
R2376 GND.t553 GND.t0 6.01393
R2377 GND.n1051 GND.t3 5.9883
R2378 GND.n645 GND.t388 5.8005
R2379 GND.n645 GND.t179 5.8005
R2380 GND.n634 GND.t19 5.8005
R2381 GND.n634 GND.t457 5.8005
R2382 GND.n635 GND.t223 5.8005
R2383 GND.n635 GND.t342 5.8005
R2384 GND.n324 GND.t502 5.8005
R2385 GND.n324 GND.t402 5.8005
R2386 GND.n322 GND.t261 5.8005
R2387 GND.n322 GND.t494 5.8005
R2388 GND.n314 GND.t627 5.8005
R2389 GND.n314 GND.t472 5.8005
R2390 GND.n315 GND.t300 5.8005
R2391 GND.n315 GND.t333 5.8005
R2392 GND.n307 GND.t590 5.8005
R2393 GND.n307 GND.t561 5.8005
R2394 GND.n305 GND.t90 5.8005
R2395 GND.n305 GND.t106 5.8005
R2396 GND.n519 GND.t155 5.8005
R2397 GND.n519 GND.t232 5.8005
R2398 GND.n518 GND.t390 5.8005
R2399 GND.n518 GND.t600 5.8005
R2400 GND.n1005 GND.t314 5.78182
R2401 GND.t65 GND.t610 5.36887
R2402 GND.n411 GND.n410 5.21334
R2403 GND.n470 GND.n469 5.21334
R2404 GND.n444 GND.n434 5.21334
R2405 GND.n1042 GND.t546 4.95592
R2406 GND.n1009 GND.n1008 4.89462
R2407 GND.n1014 GND.n1013 4.89462
R2408 GND.n1019 GND.n1018 4.89462
R2409 GND.n938 GND.n936 4.89462
R2410 GND.n932 GND.n931 4.89462
R2411 GND.n402 GND.n383 4.59029
R2412 GND.t521 GND.t463 4.54297
R2413 GND.t210 GND.t337 4.54297
R2414 GND.n1194 GND.t119 4.54297
R2415 GND.n1111 GND.t649 4.44521
R2416 GND.n1377 GND.n1376 4.33704
R2417 GND.n692 GND.n6 4.33704
R2418 GND.t289 GND.t56 4.33649
R2419 GND.n1005 GND.t465 4.33649
R2420 GND.n1153 GND 4.18987
R2421 GND.n105 GND.n104 4.17828
R2422 GND.n103 GND.n102 4.17828
R2423 GND.n403 GND.n402 4.14696
R2424 GND.n1042 GND.n1041 4.13002
R2425 GND.n1327 GND.n1326 4.00641
R2426 GND.t118 GND.n1021 3.92354
R2427 GND.n718 GND.n300 3.71362
R2428 GND.n1155 GND.n1154 3.52871
R2429 GND.n248 GND.n247 3.52871
R2430 GND.t540 GND.t45 3.13794
R2431 GND.n1101 GND.t32 3.13794
R2432 GND.n1326 GND.n1325 3.13461
R2433 GND.n1029 GND.n1028 3.1005
R2434 GND.n1155 GND.n101 3.09574
R2435 GND.n972 GND.n101 3.09574
R2436 GND.n112 GND.n100 3.09574
R2437 GND.n972 GND.n100 3.09574
R2438 GND.n248 GND.n99 2.9255
R2439 GND.n982 GND.n99 2.9255
R2440 GND.n958 GND.n98 2.9255
R2441 GND.n982 GND.n98 2.9255
R2442 GND.n401 GND.n400 2.87229
R2443 GND.n1376 GND 2.85076
R2444 GND GND.n1366 2.85076
R2445 GND GND.n9 2.85076
R2446 GND.n1378 GND.n8 2.82946
R2447 GND.t324 GND.t181 2.61503
R2448 GND.n511 GND.n510 2.5255
R2449 GND.n1112 GND.n148 2.51123
R2450 GND.n1112 GND.n1111 2.51123
R2451 GND.n394 GND.n146 2.51123
R2452 GND.n149 GND.n146 2.51123
R2453 GND.n1037 GND.n198 2.50988
R2454 GND.t308 GND.t311 2.47821
R2455 GND.t313 GND.n166 2.41134
R2456 GND.n402 GND.n401 2.33946
R2457 GND.n1154 GND.n1153 2.33915
R2458 GND.n247 GND.n8 2.33915
R2459 GND.n510 GND.n403 2.33654
R2460 GND.n693 GND.n692 2.2505
R2461 GND.n941 GND.n940 2.23675
R2462 GND.n403 GND.n7 2.20779
R2463 GND.n965 GND.n964 2.13383
R2464 GND.t271 GND.t429 2.06526
R2465 GND.n501 GND.n411 2.04483
R2466 GND.n447 GND.n434 2.04483
R2467 GND.n482 GND.n470 2.04483
R2468 GND.n1380 GND.n6 1.9555
R2469 GND.n1379 GND.n1378 1.94363
R2470 GND.n930 GND.n191 1.92706
R2471 GND.n1045 GND.n191 1.92706
R2472 GND.n898 GND.n897 1.92081
R2473 GND.n899 GND.n898 1.89738
R2474 GND.n216 GND.n205 1.87081
R2475 GND.n912 GND.n911 1.8605
R2476 GND.n928 GND.n927 1.8605
R2477 GND.n938 GND.n937 1.8605
R2478 GND.n1018 GND.n1017 1.8605
R2479 GND.n1034 GND.n1033 1.8605
R2480 GND.n919 GND.n190 1.8605
R2481 GND.n945 GND.t63 1.85878
R2482 GND GND.n644 1.85258
R2483 GND.n642 GND 1.85258
R2484 GND.n640 GND 1.85258
R2485 GND GND.n323 1.85258
R2486 GND GND.n321 1.85258
R2487 GND.n319 GND 1.85258
R2488 GND.n317 GND 1.85258
R2489 GND.n711 GND 1.85258
R2490 GND.n713 GND 1.85258
R2491 GND GND.n301 1.85258
R2492 GND.n1153 GND.n1152 1.84196
R2493 GND.n926 GND.n925 1.788
R2494 GND.n918 GND.t546 1.65231
R2495 GND.t288 GND.n1001 1.65231
R2496 GND GND.n6 1.52425
R2497 GND.n1379 GND.n7 1.48404
R2498 GND.n1027 GND.n205 1.4755
R2499 GND.t53 GND.t187 1.45963
R2500 GND.n908 GND.t65 1.44583
R2501 GND.n1052 GND.n1051 1.44583
R2502 GND.n913 GND.n200 1.3755
R2503 GND.n1022 GND.t286 1.23936
R2504 GND.n1047 GND.n189 1.21613
R2505 GND.n896 GND.n718 1.17175
R2506 GND.n896 GND.n895 1.15253
R2507 GND GND.n693 1.13527
R2508 GND.n1362 GND.n1361 1.12991
R2509 GND.n1378 GND.n1377 1.10279
R2510 GND.n1152 GND.n8 1.0655
R2511 GND.n216 GND.n215 1.04894
R2512 GND.n1015 GND.n1014 1.03383
R2513 GND.n226 GND.t497 1.03288
R2514 GND.n1047 GND.n1046 0.984875
R2515 GND GND.n941 0.977696
R2516 GND.n1046 GND.n1045 0.942687
R2517 GND.n1376 GND.n9 0.872295
R2518 GND.n527 GND.n300 0.857375
R2519 GND.n693 GND.n691 0.856945
R2520 GND.n1366 GND 0.846654
R2521 GND.n1037 GND.n1036 0.839563
R2522 GND.n1010 GND.n215 0.822375
R2523 GND.n1011 GND.n1010 0.822375
R2524 GND.n1361 GND.n14 0.753441
R2525 GND.n941 GND.n896 0.744875
R2526 GND.n931 GND.n930 0.715885
R2527 GND.n1045 GND.n1044 0.715885
R2528 GND.n930 GND.n189 0.711438
R2529 GND.n1326 GND 0.661558
R2530 GND.n521 GND 0.645031
R2531 GND GND.n520 0.645031
R2532 GND.n520 GND 0.645031
R2533 GND.n306 GND 0.645031
R2534 GND GND.n306 0.645031
R2535 GND GND.n710 0.645031
R2536 GND.n710 GND 0.645031
R2537 GND.n316 GND 0.645031
R2538 GND GND.n316 0.645031
R2539 GND.n704 GND 0.645031
R2540 GND.n704 GND 0.645031
R2541 GND GND.n703 0.645031
R2542 GND.n703 GND 0.645031
R2543 GND GND.n702 0.645031
R2544 GND.n702 GND 0.645031
R2545 GND.n636 GND 0.645031
R2546 GND GND.n636 0.645031
R2547 GND.n695 GND 0.645031
R2548 GND.n695 GND 0.645031
R2549 GND GND.n694 0.645031
R2550 GND GND.n1242 0.633946
R2551 GND.n1209 GND 0.633946
R2552 GND GND.n1227 0.633946
R2553 GND.n716 GND.n302 0.625711
R2554 GND.n1010 GND.n1009 0.6205
R2555 GND.n218 GND.n205 0.6205
R2556 GND.t465 GND.t286 0.619928
R2557 GND.n694 GND 0.608898
R2558 GND.n523 GND.n522 0.607197
R2559 GND.n1035 GND.n199 0.59425
R2560 GND.n1011 GND.n207 0.59425
R2561 GND.n1016 GND.n1015 0.568786
R2562 GND.n1152 GND.n1151 0.555206
R2563 GND.n1380 GND.n1379 0.552583
R2564 GND.n527 GND.n7 0.552583
R2565 GND.n1377 GND 0.5405
R2566 GND GND.n1253 0.51148
R2567 GND.n1026 GND.n1025 0.489974
R2568 GND.n217 GND.n216 0.489974
R2569 GND.n214 GND.n199 0.48175
R2570 GND.n1366 GND 0.473256
R2571 GND.n1015 GND.n1011 0.448938
R2572 GND.n192 GND.n191 0.423227
R2573 GND.n1048 GND.n1047 0.423227
R2574 GND.n1027 GND.n1026 0.395812
R2575 GND.n738 GND 0.390703
R2576 GND GND.n869 0.390703
R2577 GND.n770 GND 0.390703
R2578 GND GND.n841 0.390703
R2579 GND.n802 GND 0.390703
R2580 GND GND.n39 0.390703
R2581 GND.n1333 GND.n1332 0.376971
R2582 GND.n925 GND.n924 0.291125
R2583 GND.n1111 GND.n149 0.261953
R2584 GND.t181 GND.t279 0.261953
R2585 GND.n937 GND.n899 0.259875
R2586 GND.n898 GND.n213 0.238962
R2587 GND.n937 GND.n198 0.236438
R2588 GND.n927 GND.n926 0.23175
R2589 GND.n1034 GND.n200 0.23175
R2590 GND.n927 GND.n198 0.230187
R2591 GND.n912 GND.n189 0.230187
R2592 GND.n1035 GND.n1034 0.230187
R2593 GND.n1046 GND.n190 0.230187
R2594 GND.n926 GND.n912 0.228625
R2595 GND.n913 GND.n190 0.228625
R2596 GND.n1036 GND.n1035 0.227062
R2597 GND.n914 GND.n913 0.227062
R2598 GND.n692 GND 0.211237
R2599 GND.n1038 GND.n1037 0.207167
R2600 GND.t256 GND.t3 0.206976
R2601 GND.t429 GND.t208 0.206976
R2602 GND.n921 GND.t521 0.206976
R2603 GND.n1031 GND.t289 0.206976
R2604 GND.n1026 GND.n207 0.198937
R2605 GND.n511 GND.n300 0.196125
R2606 GND.n925 GND.n914 0.186437
R2607 GND.n401 GND.n394 0.164603
R2608 GND.n897 GND.n199 0.164562
R2609 GND.n207 GND.n206 0.159799
R2610 GND.n1028 GND.n1027 0.15675
R2611 GND.n1028 GND.n200 0.155187
R2612 GND.n508 GND.n405 0.120292
R2613 GND.n503 GND.n502 0.120292
R2614 GND.n500 GND.n412 0.120292
R2615 GND.n494 GND.n493 0.120292
R2616 GND.n439 GND.n438 0.120292
R2617 GND.n446 GND.n435 0.120292
R2618 GND.n448 GND.n433 0.120292
R2619 GND.n455 GND.n454 0.120292
R2620 GND.n463 GND.n427 0.120292
R2621 GND.n466 GND.n424 0.120292
R2622 GND.n481 GND.n471 0.120292
R2623 GND.n475 GND.n474 0.120292
R2624 GND.n689 GND.n688 0.120292
R2625 GND.n688 GND.n687 0.120292
R2626 GND.n687 GND.n647 0.120292
R2627 GND.n683 GND.n647 0.120292
R2628 GND.n683 GND.n682 0.120292
R2629 GND.n682 GND.n681 0.120292
R2630 GND.n678 GND.n677 0.120292
R2631 GND.n677 GND.n676 0.120292
R2632 GND.n673 GND.n672 0.120292
R2633 GND.n672 GND.n671 0.120292
R2634 GND.n671 GND.n652 0.120292
R2635 GND.n666 GND.n665 0.120292
R2636 GND.n665 GND.n664 0.120292
R2637 GND.n661 GND.n660 0.120292
R2638 GND.n660 GND.n659 0.120292
R2639 GND.n27 GND.n26 0.120292
R2640 GND.n1334 GND.n26 0.120292
R2641 GND.n1341 GND.n1340 0.120292
R2642 GND.n1350 GND.n1349 0.120292
R2643 GND.n19 GND.n18 0.120292
R2644 GND.n1355 GND.n18 0.120292
R2645 GND.n1357 GND.n16 0.120292
R2646 GND.n1364 GND.n15 0.120292
R2647 GND.n1365 GND.n1364 0.120292
R2648 GND.n1278 GND.n1276 0.120292
R2649 GND.n1279 GND.n1278 0.120292
R2650 GND.n1284 GND.n1274 0.120292
R2651 GND.n1285 GND.n1284 0.120292
R2652 GND.n1318 GND.n1286 0.120292
R2653 GND.n1314 GND.n1286 0.120292
R2654 GND.n1305 GND.n1291 0.120292
R2655 GND.n1300 GND.n1299 0.120292
R2656 GND.n1016 GND.n214 0.115419
R2657 GND GND.n489 0.112479
R2658 GND.n459 GND 0.112479
R2659 GND.n502 GND.n501 0.109875
R2660 GND.n447 GND.n446 0.109875
R2661 GND.n482 GND.n424 0.109875
R2662 GND.n689 GND 0.105969
R2663 GND.n501 GND.n500 0.104667
R2664 GND.n448 GND.n447 0.104667
R2665 GND.n482 GND.n481 0.104667
R2666 GND GND.n1380 0.10425
R2667 GND.n528 GND.n527 0.101125
R2668 GND.n278 GND 0.0866486
R2669 GND.n277 GND.n271 0.0815811
R2670 GND.n286 GND.n270 0.0815811
R2671 GND.n295 GND.n269 0.0815811
R2672 GND.n942 GND.n299 0.0815811
R2673 GND.n895 GND.n719 0.0815811
R2674 GND.n729 GND.n728 0.0815811
R2675 GND.n739 GND.n738 0.0815811
R2676 GND.n749 GND.n748 0.0815811
R2677 GND.n869 GND.n751 0.0815811
R2678 GND.n761 GND.n760 0.0815811
R2679 GND.n771 GND.n770 0.0815811
R2680 GND.n781 GND.n780 0.0815811
R2681 GND.n841 GND.n783 0.0815811
R2682 GND.n793 GND.n792 0.0815811
R2683 GND.n803 GND.n802 0.0815811
R2684 GND.n812 GND.n811 0.0815811
R2685 GND.n40 GND.n39 0.0815811
R2686 GND.n50 GND.n49 0.0815811
R2687 GND.n1253 GND.n52 0.0815811
R2688 GND.n1242 GND.n57 0.0815811
R2689 GND.n1210 GND.n1209 0.0815811
R2690 GND.n1227 GND.n1213 0.0815811
R2691 GND.n287 GND 0.0807365
R2692 GND.n296 GND 0.0807365
R2693 GND.n407 GND.n405 0.0760208
R2694 GND.n495 GND.n494 0.0760208
R2695 GND.n440 GND.n439 0.0760208
R2696 GND.n454 GND.n453 0.0760208
R2697 GND.n464 GND.n463 0.0760208
R2698 GND.n476 GND.n475 0.0760208
R2699 GND GND.n508 0.0603958
R2700 GND.n503 GND 0.0603958
R2701 GND.n496 GND 0.0603958
R2702 GND.n490 GND 0.0603958
R2703 GND.n438 GND 0.0603958
R2704 GND GND.n435 0.0603958
R2705 GND.n452 GND 0.0603958
R2706 GND.n458 GND 0.0603958
R2707 GND GND.n427 0.0603958
R2708 GND.n466 GND 0.0603958
R2709 GND.n477 GND 0.0603958
R2710 GND.n678 GND 0.0603958
R2711 GND.n673 GND 0.0603958
R2712 GND.n653 GND 0.0603958
R2713 GND.n666 GND 0.0603958
R2714 GND.n661 GND 0.0603958
R2715 GND GND.n657 0.0603958
R2716 GND.n1375 GND 0.0603958
R2717 GND GND.n27 0.0603958
R2718 GND.n1335 GND 0.0603958
R2719 GND.n1336 GND 0.0603958
R2720 GND GND.n23 0.0603958
R2721 GND.n1340 GND 0.0603958
R2722 GND.n1344 GND 0.0603958
R2723 GND.n1345 GND 0.0603958
R2724 GND.n1346 GND 0.0603958
R2725 GND.n1349 GND 0.0603958
R2726 GND GND.n19 0.0603958
R2727 GND.n1356 GND 0.0603958
R2728 GND.n1357 GND 0.0603958
R2729 GND GND.n15 0.0603958
R2730 GND.n1367 GND 0.0603958
R2731 GND.n1276 GND 0.0603958
R2732 GND GND.n1274 0.0603958
R2733 GND.n1320 GND 0.0603958
R2734 GND GND.n1319 0.0603958
R2735 GND GND.n1318 0.0603958
R2736 GND GND.n1313 0.0603958
R2737 GND GND.n1312 0.0603958
R2738 GND.n1290 GND 0.0603958
R2739 GND.n1307 GND 0.0603958
R2740 GND GND.n1306 0.0603958
R2741 GND GND.n1305 0.0603958
R2742 GND.n1301 GND 0.0603958
R2743 GND GND.n1300 0.0603958
R2744 GND.n1296 GND 0.0603958
R2745 GND GND.n1295 0.0603958
R2746 GND.n532 GND.n531 0.058
R2747 GND.n533 GND.n532 0.058
R2748 GND.n537 GND.n360 0.058
R2749 GND.n538 GND.n537 0.058
R2750 GND.n543 GND.n542 0.058
R2751 GND.n544 GND.n543 0.058
R2752 GND.n548 GND.n356 0.058
R2753 GND.n549 GND.n548 0.058
R2754 GND.n554 GND.n553 0.058
R2755 GND.n555 GND.n554 0.058
R2756 GND.n559 GND.n352 0.058
R2757 GND.n560 GND.n559 0.058
R2758 GND.n565 GND.n564 0.058
R2759 GND.n566 GND.n565 0.058
R2760 GND.n570 GND.n348 0.058
R2761 GND.n571 GND.n570 0.058
R2762 GND.n576 GND.n575 0.058
R2763 GND.n577 GND.n576 0.058
R2764 GND.n581 GND.n344 0.058
R2765 GND.n582 GND.n581 0.058
R2766 GND.n587 GND.n586 0.058
R2767 GND.n588 GND.n587 0.058
R2768 GND.n592 GND.n340 0.058
R2769 GND.n593 GND.n592 0.058
R2770 GND.n598 GND.n597 0.058
R2771 GND.n599 GND.n598 0.058
R2772 GND.n603 GND.n336 0.058
R2773 GND.n604 GND.n603 0.058
R2774 GND.n609 GND.n608 0.058
R2775 GND.n610 GND.n609 0.058
R2776 GND.n614 GND.n332 0.058
R2777 GND.n615 GND.n614 0.058
R2778 GND.n626 GND.n625 0.058
R2779 GND.n625 GND.n616 0.058
R2780 GND.n620 GND.n617 0.058
R2781 GND.n620 GND.n619 0.058
R2782 GND.n1388 GND.n1 0.058
R2783 GND.n3 GND.n1 0.058
R2784 GND.n1382 GND.n4 0.058
R2785 GND.n1382 GND.n1381 0.058
R2786 GND.n512 GND 0.0577917
R2787 GND.n281 GND.n280 0.0553986
R2788 GND.n290 GND.n289 0.0553986
R2789 GND.n298 GND.n268 0.0553986
R2790 GND.n725 GND.n724 0.0553986
R2791 GND.n735 GND.n734 0.0553986
R2792 GND.n745 GND.n740 0.0553986
R2793 GND.n872 GND.n750 0.0553986
R2794 GND.n757 GND.n756 0.0553986
R2795 GND.n767 GND.n766 0.0553986
R2796 GND.n777 GND.n772 0.0553986
R2797 GND.n844 GND.n782 0.0553986
R2798 GND.n789 GND.n788 0.0553986
R2799 GND.n799 GND.n798 0.0553986
R2800 GND.n808 GND.n804 0.0553986
R2801 GND.n816 GND.n813 0.0553986
R2802 GND.n46 GND.n41 0.0553986
R2803 GND.n1256 GND.n51 0.0553986
R2804 GND.n1245 GND.n56 0.0553986
R2805 GND.n1206 GND.n1205 0.0553986
R2806 GND.n1230 GND.n1212 0.0553986
R2807 GND.n1218 GND.n1215 0.0553986
R2808 GND.n272 GND.n271 0.0545423
R2809 GND.n166 GND.t310 0.0500323
R2810 GND.n408 GND.n407 0.0447708
R2811 GND.n496 GND.n495 0.0447708
R2812 GND.n441 GND.n440 0.0447708
R2813 GND.n453 GND.n452 0.0447708
R2814 GND.n465 GND.n464 0.0447708
R2815 GND.n477 GND.n476 0.0447708
R2816 GND GND.n277 0.0410405
R2817 GND GND.n286 0.0410405
R2818 GND GND.n295 0.0410405
R2819 GND.n942 GND 0.0410405
R2820 GND.n728 GND 0.0410405
R2821 GND.n748 GND 0.0410405
R2822 GND.n760 GND 0.0410405
R2823 GND.n780 GND 0.0410405
R2824 GND.n792 GND 0.0410405
R2825 GND.n811 GND 0.0410405
R2826 GND.n49 GND 0.0410405
R2827 GND GND.n727 0.0351284
R2828 GND GND.n747 0.0351284
R2829 GND GND.n759 0.0351284
R2830 GND GND.n779 0.0351284
R2831 GND GND.n791 0.0351284
R2832 GND GND.n810 0.0351284
R2833 GND GND.n48 0.0351284
R2834 GND.n1244 GND 0.0351284
R2835 GND GND.n1208 0.0351284
R2836 GND.n1229 GND 0.0351284
R2837 GND.n1217 GND 0.0351284
R2838 GND.n501 GND 0.0343542
R2839 GND.n447 GND 0.0343542
R2840 GND.n482 GND 0.0343542
R2841 GND GND.n1345 0.0343542
R2842 GND GND.n653 0.0330521
R2843 GND.n657 GND 0.0330521
R2844 GND GND.n1375 0.0330521
R2845 GND.n1327 GND 0.0330521
R2846 GND GND.n1335 0.0330521
R2847 GND.n1336 GND 0.0330521
R2848 GND GND.n1356 0.0330521
R2849 GND.n1367 GND 0.0330521
R2850 GND.n1325 GND 0.0330521
R2851 GND.n1320 GND 0.0330521
R2852 GND.n1312 GND 0.0330521
R2853 GND.n1307 GND 0.0330521
R2854 GND.n1295 GND 0.0330521
R2855 GND.n531 GND 0.02925
R2856 GND GND.n360 0.02925
R2857 GND.n539 GND 0.02925
R2858 GND.n542 GND 0.02925
R2859 GND GND.n356 0.02925
R2860 GND.n550 GND 0.02925
R2861 GND.n553 GND 0.02925
R2862 GND GND.n352 0.02925
R2863 GND.n561 GND 0.02925
R2864 GND.n564 GND 0.02925
R2865 GND GND.n348 0.02925
R2866 GND.n572 GND 0.02925
R2867 GND.n575 GND 0.02925
R2868 GND GND.n344 0.02925
R2869 GND.n583 GND 0.02925
R2870 GND.n586 GND 0.02925
R2871 GND GND.n340 0.02925
R2872 GND.n594 GND 0.02925
R2873 GND.n597 GND 0.02925
R2874 GND GND.n336 0.02925
R2875 GND.n605 GND 0.02925
R2876 GND.n608 GND 0.02925
R2877 GND GND.n332 0.02925
R2878 GND.n627 GND 0.02925
R2879 GND GND.n626 0.02925
R2880 GND.n617 GND 0.02925
R2881 GND GND.n0 0.02925
R2882 GND GND.n1388 0.02925
R2883 GND.n4 GND 0.02925
R2884 GND.n215 GND 0.0270625
R2885 GND.n280 GND.n270 0.0266824
R2886 GND.n289 GND.n269 0.0266824
R2887 GND.n299 GND.n298 0.0266824
R2888 GND.n725 GND.n719 0.0266824
R2889 GND.n735 GND.n729 0.0266824
R2890 GND.n745 GND.n739 0.0266824
R2891 GND.n750 GND.n749 0.0266824
R2892 GND.n757 GND.n751 0.0266824
R2893 GND.n767 GND.n761 0.0266824
R2894 GND.n777 GND.n771 0.0266824
R2895 GND.n782 GND.n781 0.0266824
R2896 GND.n789 GND.n783 0.0266824
R2897 GND.n799 GND.n793 0.0266824
R2898 GND.n808 GND.n803 0.0266824
R2899 GND.n813 GND.n812 0.0266824
R2900 GND.n46 GND.n40 0.0266824
R2901 GND.n51 GND.n50 0.0266824
R2902 GND.n56 GND.n52 0.0266824
R2903 GND.n1206 GND.n57 0.0266824
R2904 GND.n1212 GND.n1210 0.0266824
R2905 GND.n1215 GND.n1213 0.0266824
R2906 GND GND.n9 0.026141
R2907 GND GND.n737 0.0249932
R2908 GND.n871 GND 0.0249932
R2909 GND GND.n769 0.0249932
R2910 GND.n843 GND 0.0249932
R2911 GND GND.n801 0.0249932
R2912 GND.n815 GND 0.0249932
R2913 GND.n1255 GND 0.0249932
R2914 GND GND.n408 0.0239375
R2915 GND GND.n412 0.0239375
R2916 GND.n493 GND 0.0239375
R2917 GND.n490 GND 0.0239375
R2918 GND.n489 GND 0.0239375
R2919 GND.n441 GND 0.0239375
R2920 GND.n433 GND 0.0239375
R2921 GND.n455 GND 0.0239375
R2922 GND GND.n458 0.0239375
R2923 GND.n459 GND 0.0239375
R2924 GND GND.n465 0.0239375
R2925 GND GND.n471 0.0239375
R2926 GND.n474 GND 0.0239375
R2927 GND.n513 GND 0.0239375
R2928 GND.n664 GND 0.0239375
R2929 GND.n659 GND 0.0239375
R2930 GND.n23 GND 0.0239375
R2931 GND GND.n1344 0.0239375
R2932 GND.n1346 GND 0.0239375
R2933 GND.n16 GND 0.0239375
R2934 GND GND.n1290 0.0239375
R2935 GND.n1306 GND 0.0239375
R2936 GND GND.n1291 0.0239375
R2937 GND.n1301 GND 0.0239375
R2938 GND.n1299 GND 0.0239375
R2939 GND.n1296 GND 0.0239375
R2940 GND.n676 GND 0.0226354
R2941 GND.n1341 GND 0.0226354
R2942 GND.n1350 GND 0.0226354
R2943 GND GND.n1285 0.0226354
R2944 GND.n509 GND 0.0213333
R2945 GND.n681 GND 0.0213333
R2946 GND GND.n652 0.0213333
R2947 GND GND.n1334 0.0213333
R2948 GND GND.n1355 0.0213333
R2949 GND GND.n1365 0.0213333
R2950 GND.n1319 GND 0.0213333
R2951 GND.n1314 GND 0.0213333
R2952 GND.n1313 GND 0.0213333
R2953 GND.n501 GND 0.0194732
R2954 GND.n447 GND 0.0194732
R2955 GND GND.n482 0.0194732
R2956 GND.n1279 GND 0.016125
R2957 GND.n528 GND 0.016125
R2958 GND.n539 GND 0.016125
R2959 GND.n550 GND 0.016125
R2960 GND.n561 GND 0.016125
R2961 GND.n572 GND 0.016125
R2962 GND.n583 GND 0.016125
R2963 GND.n594 GND 0.016125
R2964 GND.n605 GND 0.016125
R2965 GND.n627 GND 0.016125
R2966 GND GND.n0 0.016125
R2967 GND.n691 GND 0.0148229
R2968 GND.n940 GND.n899 0.01175
R2969 GND.n1017 GND.n199 0.011346
R2970 GND.n533 GND 0.011125
R2971 GND GND.n538 0.011125
R2972 GND.n544 GND 0.011125
R2973 GND GND.n549 0.011125
R2974 GND.n555 GND 0.011125
R2975 GND GND.n560 0.011125
R2976 GND.n566 GND 0.011125
R2977 GND GND.n571 0.011125
R2978 GND.n577 GND 0.011125
R2979 GND GND.n582 0.011125
R2980 GND.n588 GND 0.011125
R2981 GND GND.n593 0.011125
R2982 GND.n599 GND 0.011125
R2983 GND GND.n604 0.011125
R2984 GND.n610 GND 0.011125
R2985 GND GND.n615 0.011125
R2986 GND GND.n616 0.011125
R2987 GND.n619 GND 0.011125
R2988 GND GND.n3 0.011125
R2989 GND.n1381 GND 0.011125
R2990 GND.n1017 GND.n1016 0.00646529
R2991 GND.n281 GND.n278 0.00641216
R2992 GND.n290 GND.n287 0.00641216
R2993 GND.n296 GND.n268 0.00641216
R2994 GND.n727 GND.n724 0.00641216
R2995 GND.n737 GND.n734 0.00641216
R2996 GND.n747 GND.n740 0.00641216
R2997 GND.n872 GND.n871 0.00641216
R2998 GND.n759 GND.n756 0.00641216
R2999 GND.n769 GND.n766 0.00641216
R3000 GND.n779 GND.n772 0.00641216
R3001 GND.n844 GND.n843 0.00641216
R3002 GND.n791 GND.n788 0.00641216
R3003 GND.n801 GND.n798 0.00641216
R3004 GND.n810 GND.n804 0.00641216
R3005 GND.n816 GND.n815 0.00641216
R3006 GND.n48 GND.n41 0.00641216
R3007 GND.n1256 GND.n1255 0.00641216
R3008 GND.n1245 GND.n1244 0.00641216
R3009 GND.n1208 GND.n1205 0.00641216
R3010 GND.n1230 GND.n1229 0.00641216
R3011 GND.n1218 GND.n1217 0.00641216
R3012 GND.n513 GND.n512 0.00310417
R3013 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t5 222.043
R3014 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t3 222.043
R3015 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n27 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t1 140.061
R3016 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n28 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t0 139.566
R3017 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t8 126.178
R3018 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t24 124.9
R3019 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t19 124.9
R3020 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t14 124.9
R3021 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t13 124.9
R3022 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t7 124.9
R3023 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t23 124.9
R3024 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t22 124.9
R3025 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t18 124.9
R3026 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t17 124.9
R3027 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t12 124.9
R3028 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t11 124.9
R3029 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t6 124.9
R3030 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t28 124.9
R3031 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t10 124.9
R3032 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t9 124.9
R3033 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t26 124.9
R3034 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t25 124.9
R3035 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t21 124.9
R3036 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t20 124.9
R3037 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t16 124.9
R3038 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t15 124.9
R3039 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t4 108.754
R3040 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n25 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t2 108.365
R3041 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t27 20.8855
R3042 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 9.08711
R3043 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n26 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n25 7.91883
R3044 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n27 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n26 5.02291
R3045 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n21 3.41379
R3046 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n28 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n27 3.40258
R3047 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n19 1.27824
R3048 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n17 1.27824
R3049 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n15 1.27824
R3050 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n13 1.27824
R3051 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n11 1.27824
R3052 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n9 1.27824
R3053 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n7 1.27824
R3054 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n5 1.27824
R3055 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n3 1.27824
R3056 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n1 1.27824
R3057 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R3058 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n18 0.391454
R3059 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R3060 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n16 0.391454
R3061 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R3062 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n14 0.391454
R3063 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R3064 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n12 0.391454
R3065 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R3066 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n10 0.391454
R3067 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R3068 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n8 0.391454
R3069 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R3070 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n6 0.391454
R3071 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R3072 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n4 0.391454
R3073 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R3074 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n2 0.391454
R3075 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.391454
R3076 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n0 0.391454
R3077 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n25 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n24 0.310917
R3078 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n26 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n22 0.270394
R3079 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n20 0.266454
R3080 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n23 0.224458
R3081 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n28 0.063
R3082 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.0498421
R3083 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t1 227.856
R3084 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n2 152.333
R3085 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t3 140.382
R3086 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t4 114.031
R3087 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t0 83.3993
R3088 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.t2 81.5883
R3089 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n3 14.4422
R3090 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n1 7.56882
R3091 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n0 5.08175
R3092 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R3093 a_42781_10934.t0 a_42781_10934.t1 114.052
R3094 top_segment_2_0.DEC2[1].n0 top_segment_2_0.DEC2[1].t1 334.771
R3095 top_segment_2_0.DEC2[1].n5 top_segment_2_0.DEC2[1].t16 213.218
R3096 top_segment_2_0.DEC2[1].n13 top_segment_2_0.DEC2[1].t13 213.218
R3097 top_segment_2_0.DEC2[1].n18 top_segment_2_0.DEC2[1].t24 213.218
R3098 top_segment_2_0.DEC2[1] top_segment_2_0.DEC2[1].t20 212.899
R3099 top_segment_2_0.DEC2[1].n10 top_segment_2_0.DEC2[1].t11 212.554
R3100 top_segment_2_0.DEC2[1].n9 top_segment_2_0.DEC2[1].t8 212.554
R3101 top_segment_2_0.DEC2[1].n8 top_segment_2_0.DEC2[1].t3 212.554
R3102 top_segment_2_0.DEC2[1].n7 top_segment_2_0.DEC2[1].t22 212.554
R3103 top_segment_2_0.DEC2[1].n6 top_segment_2_0.DEC2[1].t9 212.554
R3104 top_segment_2_0.DEC2[1].n5 top_segment_2_0.DEC2[1].t19 212.554
R3105 top_segment_2_0.DEC2[1].n13 top_segment_2_0.DEC2[1].t10 212.554
R3106 top_segment_2_0.DEC2[1].n14 top_segment_2_0.DEC2[1].t5 212.554
R3107 top_segment_2_0.DEC2[1].n15 top_segment_2_0.DEC2[1].t2 212.554
R3108 top_segment_2_0.DEC2[1].n16 top_segment_2_0.DEC2[1].t23 212.554
R3109 top_segment_2_0.DEC2[1].n17 top_segment_2_0.DEC2[1].t6 212.554
R3110 top_segment_2_0.DEC2[1].n4 top_segment_2_0.DEC2[1].t15 208.054
R3111 top_segment_2_0.DEC2[1].n12 top_segment_2_0.DEC2[1].t12 208.054
R3112 top_segment_2_0.DEC2[1].n19 top_segment_2_0.DEC2[1].t18 208.054
R3113 top_segment_2_0.DEC2[1].n23 top_segment_2_0.DEC2[1].n22 152
R3114 top_segment_2_0.DEC2[1].n3 top_segment_2_0.DEC2[1].t4 131.306
R3115 top_segment_2_0.DEC2[1].n1 top_segment_2_0.DEC2[1].t17 126.278
R3116 top_segment_2_0.DEC2[1].n1 top_segment_2_0.DEC2[1].t7 125.566
R3117 top_segment_2_0.DEC2[1].n22 top_segment_2_0.DEC2[1].t21 114.031
R3118 top_segment_2_0.DEC2[1].n0 top_segment_2_0.DEC2[1].t0 87.8231
R3119 top_segment_2_0.DEC2[1].n22 top_segment_2_0.DEC2[1].t14 81.5883
R3120 top_segment_2_0.DEC2[1] top_segment_2_0.DEC2[1].n21 34.7422
R3121 top_segment_2_0.DEC2[1].n21 top_segment_2_0.DEC2[1].n4 31.4317
R3122 top_segment_2_0.DEC2[1].n21 top_segment_2_0.DEC2[1].n20 28.8753
R3123 top_segment_2_0.DEC2[1].n24 top_segment_2_0.DEC2[1] 14.6403
R3124 top_segment_2_0.DEC2[1] top_segment_2_0.DEC2[1].n23 11.4706
R3125 top_segment_2_0.DEC2[1] top_segment_2_0.DEC2[1].n3 5.12863
R3126 top_segment_2_0.DEC2[1].n4 top_segment_2_0.DEC2[1] 4.82021
R3127 top_segment_2_0.DEC2[1].n2 top_segment_2_0.DEC2[1].n1 4.68383
R3128 top_segment_2_0.DEC2[1].n12 top_segment_2_0.DEC2[1].n11 4.5005
R3129 top_segment_2_0.DEC2[1].n19 top_segment_2_0.DEC2[1].n18 4.5005
R3130 top_segment_2_0.DEC2[1].n23 top_segment_2_0.DEC2[1] 4.48881
R3131 top_segment_2_0.DEC2[1].n20 top_segment_2_0.DEC2[1].n19 2.63367
R3132 top_segment_2_0.DEC2[1] top_segment_2_0.DEC2[1].n24 1.01821
R3133 top_segment_2_0.DEC2[1].n24 top_segment_2_0.DEC2[1] 0.7755
R3134 top_segment_2_0.DEC2[1].n6 top_segment_2_0.DEC2[1].n5 0.663962
R3135 top_segment_2_0.DEC2[1].n7 top_segment_2_0.DEC2[1].n6 0.663962
R3136 top_segment_2_0.DEC2[1].n8 top_segment_2_0.DEC2[1].n7 0.663962
R3137 top_segment_2_0.DEC2[1].n9 top_segment_2_0.DEC2[1].n8 0.663962
R3138 top_segment_2_0.DEC2[1].n10 top_segment_2_0.DEC2[1].n9 0.663962
R3139 top_segment_2_0.DEC2[1].n11 top_segment_2_0.DEC2[1].n10 0.663962
R3140 top_segment_2_0.DEC2[1].n18 top_segment_2_0.DEC2[1].n17 0.663962
R3141 top_segment_2_0.DEC2[1].n17 top_segment_2_0.DEC2[1].n16 0.663962
R3142 top_segment_2_0.DEC2[1].n16 top_segment_2_0.DEC2[1].n15 0.663962
R3143 top_segment_2_0.DEC2[1].n15 top_segment_2_0.DEC2[1].n14 0.663962
R3144 top_segment_2_0.DEC2[1].n14 top_segment_2_0.DEC2[1].n13 0.663962
R3145 top_segment_2_0.DEC2[1].n2 top_segment_2_0.DEC2[1].n0 0.608192
R3146 top_segment_2_0.DEC2[1].n20 top_segment_2_0.DEC2[1].n12 0.34425
R3147 top_segment_2_0.DEC2[1].n11 top_segment_2_0.DEC2[1] 0.269731
R3148 top_segment_2_0.DEC2[1].n3 top_segment_2_0.DEC2[1].n2 0.177583
R3149 a_26719_5238.n2 a_26719_5238.t2 247.918
R3150 a_26719_5238.n0 a_26719_5238.t1 245.935
R3151 a_26719_5238.n1 a_26719_5238.t4 245.381
R3152 a_26719_5238.n0 a_26719_5238.t3 239.267
R3153 a_26719_5238.t0 a_26719_5238.n2 239.267
R3154 a_26719_5238.n1 a_26719_5238.n0 6.24633
R3155 a_26719_5238.n2 a_26719_5238.n1 0.7755
R3156 top_segment_1_0.rseg_1_v3_1.v19 top_segment_1_0.rseg_1_v3_1.v19.t0 245.726
R3157 top_segment_1_0.rseg_1_v3_1.v19.n0 top_segment_1_0.rseg_1_v3_1.v19.t1 10.6701
R3158 top_segment_1_0.rseg_1_v3_1.v19.n0 top_segment_1_0.rseg_1_v3_1.v19.t2 10.5739
R3159 top_segment_1_0.rseg_1_v3_1.v19 top_segment_1_0.rseg_1_v3_1.v19.n0 1.51759
R3160 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 272.038
R3161 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t0 258.846
R3162 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t3 230.363
R3163 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n0 224.776
R3164 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t4 158.064
R3165 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n1 152.292
R3166 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t2 26.5955
R3167 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.t1 26.5955
R3168 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 24.0946
R3169 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n2 20.0033
R3170 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 6.4005
R3171 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 3.76521
R3172 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n4 3.03935
R3173 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 2.30266
R3174 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n3 1.50638
R3175 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y.n5 0.921363
R3176 VDD.n238 VDD.t67 674.802
R3177 VDD.n84 VDD.n83 674.766
R3178 VDD.n142 VDD.n115 674.766
R3179 VDD.n440 VDD.t98 633.369
R3180 VDD.t169 VDD.n276 553.428
R3181 VDD.t182 VDD.n81 465.683
R3182 VDD.n277 VDD 432.123
R3183 VDD.n313 VDD.t69 420.43
R3184 VDD.n439 VDD.t144 420.25
R3185 VDD.t88 VDD.n15 420.25
R3186 VDD.t192 VDD.n19 420.25
R3187 VDD.t90 VDD.n23 420.25
R3188 VDD.t113 VDD.n27 420.25
R3189 VDD.t49 VDD.n31 420.25
R3190 VDD.t41 VDD.n35 420.25
R3191 VDD.t35 VDD.n39 420.25
R3192 VDD.n43 VDD.t25 420.25
R3193 VDD.n83 VDD.t157 414.33
R3194 VDD.n142 VDD.t29 414.33
R3195 VDD.t107 VDD 411.372
R3196 VDD VDD.n141 401.233
R3197 VDD VDD.t213 369.938
R3198 VDD.t63 VDD 369.938
R3199 VDD.t217 VDD 369.938
R3200 VDD.t80 VDD 369.938
R3201 VDD.t56 VDD 369.938
R3202 VDD.t139 VDD 369.938
R3203 VDD.t119 VDD 369.938
R3204 VDD.t86 VDD 369.938
R3205 VDD.t82 VDD 369.938
R3206 VDD VDD.t123 369.938
R3207 VDD VDD.t153 366.978
R3208 VDD.t159 VDD 366.978
R3209 VDD.t103 VDD 361.06
R3210 VDD.t179 VDD 361.06
R3211 VDD.t96 VDD 361.06
R3212 VDD VDD.t221 361.06
R3213 VDD VDD.t117 361.06
R3214 VDD VDD.t142 361.06
R3215 VDD VDD.t37 361.06
R3216 VDD VDD.t10 361.06
R3217 VDD VDD.t0 361.06
R3218 VDD VDD.t21 361.06
R3219 VDD.t6 VDD 361.06
R3220 VDD.n218 VDD.t18 340.301
R3221 VDD.n298 VDD.t201 340.301
R3222 VDD.n201 VDD.t156 336.416
R3223 VDD.n307 VDD.n208 327.377
R3224 VDD.n228 VDD.n227 320.976
R3225 VDD.n223 VDD.n221 320.976
R3226 VDD.n325 VDD.n324 318.305
R3227 VDD.n300 VDD.n212 318.305
R3228 VDD.n191 VDD.n190 318.303
R3229 VDD VDD.t169 313.707
R3230 VDD.n183 VDD.n160 313.575
R3231 VDD.n154 VDD.n153 278.858
R3232 VDD.n155 VDD.n153 278.858
R3233 VDD.n332 VDD.n153 278.858
R3234 VDD.n330 VDD.n153 278.858
R3235 VDD.n164 VDD.n163 278.858
R3236 VDD.n163 VDD.n162 278.858
R3237 VDD.n163 VDD.n152 278.858
R3238 VDD.n81 VDD 270.827
R3239 VDD.n85 VDD 270.827
R3240 VDD.n82 VDD 270.827
R3241 VDD.n114 VDD 270.827
R3242 VDD.n143 VDD 270.827
R3243 VDD.n161 VDD.n152 269.485
R3244 VDD.n332 VDD.n331 269.485
R3245 VDD.n162 VDD.n161 269.485
R3246 VDD.n331 VDD.n155 269.485
R3247 VDD.n164 VDD.n161 269.485
R3248 VDD.n331 VDD.n154 269.485
R3249 VDD.n331 VDD.n330 269.485
R3250 VDD.n81 VDD.n80 267.296
R3251 VDD.n86 VDD.n85 267.296
R3252 VDD.n82 VDD.n54 267.296
R3253 VDD.n114 VDD.n113 267.296
R3254 VDD.n144 VDD.n143 267.296
R3255 VDD.n344 VDD.t124 255.905
R3256 VDD.n42 VDD.t26 255.905
R3257 VDD.n355 VDD.t83 255.905
R3258 VDD.n38 VDD.t36 255.905
R3259 VDD.n366 VDD.t87 255.905
R3260 VDD.n34 VDD.t42 255.905
R3261 VDD.n377 VDD.t120 255.905
R3262 VDD.n30 VDD.t50 255.905
R3263 VDD.n388 VDD.t140 255.905
R3264 VDD.n26 VDD.t114 255.905
R3265 VDD.n399 VDD.t57 255.905
R3266 VDD.n22 VDD.t91 255.905
R3267 VDD.n410 VDD.t81 255.905
R3268 VDD.n18 VDD.t193 255.905
R3269 VDD.n421 VDD.t218 255.905
R3270 VDD.n14 VDD.t89 255.905
R3271 VDD.n432 VDD.t64 255.905
R3272 VDD.n3 VDD.t145 255.905
R3273 VDD.n8 VDD.t214 255.905
R3274 VDD.n441 VDD.t99 255.905
R3275 VDD.n189 VDD.t181 255.905
R3276 VDD.n270 VDD.t170 255.905
R3277 VDD.n203 VDD.t146 255.905
R3278 VDD.n195 VDD.t51 255.904
R3279 VDD.n203 VDD.t70 255.904
R3280 VDD.n340 VDD.t126 252.95
R3281 VDD.n345 VDD.t28 252.95
R3282 VDD.n351 VDD.t9 252.95
R3283 VDD.n356 VDD.t46 252.95
R3284 VDD.n362 VDD.t3 252.95
R3285 VDD.n367 VDD.t24 252.95
R3286 VDD.n373 VDD.t122 252.95
R3287 VDD.n378 VDD.t203 252.95
R3288 VDD.n384 VDD.t110 252.95
R3289 VDD.n389 VDD.t116 252.95
R3290 VDD.n395 VDD.t77 252.95
R3291 VDD.n400 VDD.t93 252.95
R3292 VDD.n406 VDD.t79 252.95
R3293 VDD.n411 VDD.t195 252.95
R3294 VDD.n417 VDD.t220 252.95
R3295 VDD.n422 VDD.t167 252.95
R3296 VDD.n428 VDD.t66 252.95
R3297 VDD.n433 VDD.t150 252.95
R3298 VDD.n4 VDD.t216 252.95
R3299 VDD.n7 VDD.t101 252.95
R3300 VDD.n210 VDD.t59 250.722
R3301 VDD.n187 VDD.t131 249.901
R3302 VDD.n181 VDD.t168 249.52
R3303 VDD.n298 VDD.t133 249.52
R3304 VDD.n329 VDD.t44 249.387
R3305 VDD.n167 VDD.t134 249.363
R3306 VDD.n177 VDD.t173 249.363
R3307 VDD.n258 VDD.t7 249.363
R3308 VDD.n263 VDD.t160 249.363
R3309 VDD.n247 VDD.t22 249.363
R3310 VDD.n235 VDD.t154 249.363
R3311 VDD.n56 VDD.t183 249.362
R3312 VDD.n74 VDD.t104 249.362
R3313 VDD.n69 VDD.t180 249.362
R3314 VDD.n66 VDD.t97 249.362
R3315 VDD.n92 VDD.t158 249.362
R3316 VDD.n97 VDD.t222 249.362
R3317 VDD.n102 VDD.t118 249.362
R3318 VDD.n107 VDD.t143 249.362
R3319 VDD.n48 VDD.t30 249.362
R3320 VDD.n125 VDD.t38 249.362
R3321 VDD.n130 VDD.t11 249.362
R3322 VDD.n135 VDD.t1 249.362
R3323 VDD.n167 VDD.t196 249.362
R3324 VDD.n177 VDD.t141 249.362
R3325 VDD.n301 VDD.t72 249.362
R3326 VDD.n283 VDD.t164 249.062
R3327 VDD.n219 VDD.t185 249.062
R3328 VDD.n294 VDD.t152 248.929
R3329 VDD.t105 VDD.t182 248.599
R3330 VDD.t33 VDD.t103 248.599
R3331 VDD.t52 VDD.t179 248.599
R3332 VDD.t39 VDD.t96 248.599
R3333 VDD.t157 VDD.t207 248.599
R3334 VDD.t221 VDD.t205 248.599
R3335 VDD.t117 VDD.t19 248.599
R3336 VDD.t142 VDD.t177 248.599
R3337 VDD.t29 VDD.t61 248.599
R3338 VDD.t37 VDD.t12 248.599
R3339 VDD.t10 VDD.t111 248.599
R3340 VDD.t0 VDD.t94 248.599
R3341 VDD.t98 VDD.t100 248.599
R3342 VDD.t213 VDD.t215 248.599
R3343 VDD.t149 VDD.t144 248.599
R3344 VDD.t65 VDD.t63 248.599
R3345 VDD.t166 VDD.t88 248.599
R3346 VDD.t219 VDD.t217 248.599
R3347 VDD.t194 VDD.t192 248.599
R3348 VDD.t78 VDD.t80 248.599
R3349 VDD.t92 VDD.t90 248.599
R3350 VDD.t76 VDD.t56 248.599
R3351 VDD.t115 VDD.t113 248.599
R3352 VDD.t109 VDD.t139 248.599
R3353 VDD.t202 VDD.t49 248.599
R3354 VDD.t121 VDD.t119 248.599
R3355 VDD.t23 VDD.t41 248.599
R3356 VDD.t2 VDD.t86 248.599
R3357 VDD.t45 VDD.t35 248.599
R3358 VDD.t8 VDD.t82 248.599
R3359 VDD.t25 VDD.t27 248.599
R3360 VDD.t123 VDD.t125 248.599
R3361 VDD.t153 VDD.t190 248.599
R3362 VDD.t21 VDD.t127 248.599
R3363 VDD.t209 VDD.t159 248.599
R3364 VDD.t197 VDD.t6 248.599
R3365 VDD.n170 VDD.t223 247.394
R3366 VDD.n175 VDD.t138 247.394
R3367 VDD.n230 VDD.t198 247.394
R3368 VDD.n259 VDD.t210 247.394
R3369 VDD.n232 VDD.t128 247.394
R3370 VDD.n246 VDD.t191 247.394
R3371 VDD.n283 VDD.t85 247.394
R3372 VDD.n219 VDD.t32 247.394
R3373 VDD.n75 VDD.t106 247.394
R3374 VDD.n59 VDD.t34 247.394
R3375 VDD.n67 VDD.t53 247.394
R3376 VDD.n55 VDD.t40 247.394
R3377 VDD.n96 VDD.t208 247.394
R3378 VDD.n101 VDD.t206 247.394
R3379 VDD.n106 VDD.t20 247.394
R3380 VDD.n49 VDD.t178 247.394
R3381 VDD.n124 VDD.t62 247.394
R3382 VDD.n129 VDD.t13 247.394
R3383 VDD.n134 VDD.t112 247.394
R3384 VDD.n116 VDD.t95 247.394
R3385 VDD.n170 VDD.t135 247.394
R3386 VDD.n175 VDD.t15 247.394
R3387 VDD.n181 VDD.t16 247.394
R3388 VDD.n299 VDD.t55 247.394
R3389 VDD.n288 VDD.t189 245.178
R3390 VDD.n217 VDD.t172 245.178
R3391 VDD.n302 VDD.t130 245.178
R3392 VDD.n158 VDD.t165 245.178
R3393 VDD.n268 VDD.t108 243.512
R3394 VDD.n239 VDD.t68 243.512
R3395 VDD.n289 VDD.t212 243.508
R3396 VDD.n282 VDD 230.766
R3397 VDD VDD.n439 221.964
R3398 VDD.n15 VDD 221.964
R3399 VDD.n19 VDD 221.964
R3400 VDD.n23 VDD 221.964
R3401 VDD.n27 VDD 221.964
R3402 VDD.n31 VDD 221.964
R3403 VDD.n35 VDD 221.964
R3404 VDD.n39 VDD 221.964
R3405 VDD.n43 VDD 221.964
R3406 VDD.n84 VDD 219.004
R3407 VDD.n115 VDD 219.004
R3408 VDD.n276 VDD 219.004
R3409 VDD.n295 VDD.n294 213.119
R3410 VDD.n308 VDD.n207 213.119
R3411 VDD.n439 VDD.n438 213.119
R3412 VDD.n427 VDD.n15 213.119
R3413 VDD.n416 VDD.n19 213.119
R3414 VDD.n405 VDD.n23 213.119
R3415 VDD.n394 VDD.n27 213.119
R3416 VDD.n383 VDD.n31 213.119
R3417 VDD.n372 VDD.n35 213.119
R3418 VDD.n361 VDD.n39 213.119
R3419 VDD.n350 VDD.n43 213.119
R3420 VDD.n276 VDD.n275 213.119
R3421 VDD.t67 VDD.t224 213.084
R3422 VDD.t60 VDD.t107 213.084
R3423 VDD.n297 VDD.n296 209.368
R3424 VDD.n312 VDD.n311 209.368
R3425 VDD VDD.t105 207.166
R3426 VDD VDD.t33 207.166
R3427 VDD VDD.t52 207.166
R3428 VDD VDD.t39 207.166
R3429 VDD.t207 VDD 207.166
R3430 VDD.t205 VDD 207.166
R3431 VDD.t19 VDD 207.166
R3432 VDD.t177 VDD 207.166
R3433 VDD.t61 VDD 207.166
R3434 VDD.t12 VDD 207.166
R3435 VDD.t111 VDD 207.166
R3436 VDD.t94 VDD 207.166
R3437 VDD.t190 VDD 207.166
R3438 VDD.t127 VDD 207.166
R3439 VDD VDD.t209 207.166
R3440 VDD VDD.t197 207.166
R3441 VDD.t71 VDD 206.45
R3442 VDD.t100 VDD 198.287
R3443 VDD.t215 VDD 198.287
R3444 VDD VDD.t149 198.287
R3445 VDD VDD.t65 198.287
R3446 VDD VDD.t166 198.287
R3447 VDD VDD.t219 198.287
R3448 VDD VDD.t194 198.287
R3449 VDD VDD.t78 198.287
R3450 VDD VDD.t92 198.287
R3451 VDD VDD.t76 198.287
R3452 VDD VDD.t115 198.287
R3453 VDD VDD.t109 198.287
R3454 VDD VDD.t202 198.287
R3455 VDD VDD.t121 198.287
R3456 VDD VDD.t23 198.287
R3457 VDD VDD.t2 198.287
R3458 VDD VDD.t45 198.287
R3459 VDD VDD.t8 198.287
R3460 VDD.t27 VDD 198.287
R3461 VDD.t125 VDD 198.287
R3462 VDD.t224 VDD 189.409
R3463 VDD VDD.t60 189.409
R3464 VDD.t69 VDD 177.916
R3465 VDD.t147 VDD.t174 140.989
R3466 VDD.t54 VDD.t71 140.989
R3467 VDD.t211 VDD.t151 140.989
R3468 VDD.t161 VDD.t171 134.276
R3469 VDD.t4 VDD.t31 134.276
R3470 VDD.t188 VDD.t136 134.276
R3471 VDD.t84 VDD.t47 134.276
R3472 VDD VDD.n312 125.883
R3473 VDD VDD.n295 124.206
R3474 VDD VDD.t129 107.421
R3475 VDD VDD.t132 107.421
R3476 VDD.t184 VDD 107.421
R3477 VDD VDD.t163 107.421
R3478 VDD.t174 VDD.n207 100.707
R3479 VDD.n296 VDD.t161 100.707
R3480 VDD VDD.t186 97.3503
R3481 VDD.n312 VDD.t155 93.9934
R3482 VDD VDD.t17 90.6365
R3483 VDD.n295 VDD.t151 80.5659
R3484 VDD.n165 VDD.n154 76.0729
R3485 VDD.n155 VDD.n151 76.0729
R3486 VDD.n333 VDD.n332 76.0729
R3487 VDD.n330 VDD.n329 76.0729
R3488 VDD.n165 VDD.n164 76.0728
R3489 VDD.n162 VDD.n151 76.0728
R3490 VDD.n333 VDD.n152 76.0728
R3491 VDD.t58 VDD.t147 72.1736
R3492 VDD.t136 VDD 70.4952
R3493 VDD.t129 VDD.t58 68.8168
R3494 VDD.t200 VDD 67.1383
R3495 VDD.n207 VDD.t155 60.4245
R3496 VDD.n296 VDD.t200 60.4245
R3497 VDD.n143 VDD.n142 51.3536
R3498 VDD.n115 VDD.n114 51.3536
R3499 VDD.n83 VDD.n82 51.3536
R3500 VDD.n85 VDD.n84 51.3536
R3501 VDD.n161 VDD 48.6651
R3502 VDD.n318 VDD.n317 43.9358
R3503 VDD.t132 VDD 43.6401
R3504 VDD.n160 VDD.t73 38.4155
R3505 VDD.n190 VDD.t75 38.4155
R3506 VDD.n324 VDD.t204 38.4155
R3507 VDD.n212 VDD.t176 38.4155
R3508 VDD.n331 VDD 36.603
R3509 VDD.n318 VDD.n197 34.6358
R3510 VDD.n322 VDD.n197 34.6358
R3511 VDD.n323 VDD.n322 34.6358
R3512 VDD.n264 VDD.n252 34.6358
R3513 VDD.n271 VDD.n231 34.6358
R3514 VDD.n241 VDD.n240 34.6358
R3515 VDD.n204 VDD.n199 34.6358
R3516 VDD.n311 VDD.n200 34.6358
R3517 VDD.n297 VDD.n217 33.5064
R3518 VDD.n183 VDD.n182 33.1299
R3519 VDD.n289 VDD.n288 33.1299
R3520 VDD.n141 VDD.n140 32.4116
R3521 VDD.n284 VDD.n228 30.8711
R3522 VDD.n224 VDD.n223 30.8711
R3523 VDD.n191 VDD.n156 27.4829
R3524 VDD.n325 VDD.n323 27.4829
R3525 VDD.t17 VDD.t211 26.8556
R3526 VDD.n160 VDD.t74 26.5955
R3527 VDD.n190 VDD.t102 26.5955
R3528 VDD.n324 VDD.t199 26.5955
R3529 VDD.n227 VDD.t137 26.5955
R3530 VDD.n227 VDD.t48 26.5955
R3531 VDD.n221 VDD.t162 26.5955
R3532 VDD.n221 VDD.t5 26.5955
R3533 VDD.n208 VDD.t175 26.5955
R3534 VDD.n208 VDD.t148 26.5955
R3535 VDD.n212 VDD.t187 26.5955
R3536 VDD.n76 VDD.n56 25.977
R3537 VDD.n74 VDD.n73 25.977
R3538 VDD.n69 VDD.n68 25.977
R3539 VDD.n66 VDD.n65 25.977
R3540 VDD.n92 VDD.n53 25.977
R3541 VDD.n97 VDD.n52 25.977
R3542 VDD.n102 VDD.n51 25.977
R3543 VDD.n108 VDD.n107 25.977
R3544 VDD.n120 VDD.n48 25.977
R3545 VDD.n125 VDD.n119 25.977
R3546 VDD.n130 VDD.n118 25.977
R3547 VDD.n136 VDD.n135 25.977
R3548 VDD.n171 VDD.n167 25.977
R3549 VDD.n177 VDD.n176 25.977
R3550 VDD.n188 VDD.n187 25.977
R3551 VDD.n258 VDD.n254 25.977
R3552 VDD.n263 VDD.n253 25.977
R3553 VDD.n248 VDD.n247 25.977
R3554 VDD.n245 VDD.n235 25.977
R3555 VDD.n344 VDD.n45 25.224
R3556 VDD.n340 VDD.n45 25.224
R3557 VDD.n346 VDD.n42 25.224
R3558 VDD.n346 VDD.n345 25.224
R3559 VDD.n355 VDD.n41 25.224
R3560 VDD.n351 VDD.n41 25.224
R3561 VDD.n357 VDD.n38 25.224
R3562 VDD.n357 VDD.n356 25.224
R3563 VDD.n366 VDD.n37 25.224
R3564 VDD.n362 VDD.n37 25.224
R3565 VDD.n368 VDD.n34 25.224
R3566 VDD.n368 VDD.n367 25.224
R3567 VDD.n377 VDD.n33 25.224
R3568 VDD.n373 VDD.n33 25.224
R3569 VDD.n379 VDD.n30 25.224
R3570 VDD.n379 VDD.n378 25.224
R3571 VDD.n388 VDD.n29 25.224
R3572 VDD.n384 VDD.n29 25.224
R3573 VDD.n390 VDD.n26 25.224
R3574 VDD.n390 VDD.n389 25.224
R3575 VDD.n399 VDD.n25 25.224
R3576 VDD.n395 VDD.n25 25.224
R3577 VDD.n401 VDD.n22 25.224
R3578 VDD.n401 VDD.n400 25.224
R3579 VDD.n410 VDD.n21 25.224
R3580 VDD.n406 VDD.n21 25.224
R3581 VDD.n412 VDD.n18 25.224
R3582 VDD.n412 VDD.n411 25.224
R3583 VDD.n421 VDD.n17 25.224
R3584 VDD.n417 VDD.n17 25.224
R3585 VDD.n423 VDD.n14 25.224
R3586 VDD.n423 VDD.n422 25.224
R3587 VDD.n432 VDD.n13 25.224
R3588 VDD.n428 VDD.n13 25.224
R3589 VDD.n434 VDD.n3 25.224
R3590 VDD.n434 VDD.n433 25.224
R3591 VDD.n9 VDD.n8 25.224
R3592 VDD.n9 VDD.n4 25.224
R3593 VDD.n441 VDD.n2 25.224
R3594 VDD.n7 VDD.n2 25.224
R3595 VDD.n80 VDD.n79 25.1591
R3596 VDD.n87 VDD.n86 25.1591
R3597 VDD.n91 VDD.n54 25.1591
R3598 VDD.n113 VDD.n112 25.1591
R3599 VDD.n145 VDD.n144 25.1591
R3600 VDD.n76 VDD.n75 24.4711
R3601 VDD.n73 VDD.n59 24.4711
R3602 VDD.n68 VDD.n67 24.4711
R3603 VDD.n65 VDD.n55 24.4711
R3604 VDD.n96 VDD.n53 24.4711
R3605 VDD.n101 VDD.n52 24.4711
R3606 VDD.n106 VDD.n51 24.4711
R3607 VDD.n108 VDD.n49 24.4711
R3608 VDD.n124 VDD.n120 24.4711
R3609 VDD.n129 VDD.n119 24.4711
R3610 VDD.n134 VDD.n118 24.4711
R3611 VDD.n136 VDD.n116 24.4711
R3612 VDD.n171 VDD.n170 24.4711
R3613 VDD.n176 VDD.n175 24.4711
R3614 VDD.n182 VDD.n181 24.4711
R3615 VDD.n254 VDD.n230 24.4711
R3616 VDD.n259 VDD.n253 24.4711
R3617 VDD.n269 VDD.n268 24.4711
R3618 VDD.n248 VDD.n232 24.4711
R3619 VDD.n246 VDD.n245 24.4711
R3620 VDD.n284 VDD.n283 24.4711
R3621 VDD.n307 VDD.n306 24.4711
R3622 VDD.n224 VDD.n219 24.4711
R3623 VDD.n329 VDD.n156 23.7181
R3624 VDD.n329 VDD.n328 23.7181
R3625 VDD.n264 VDD.n263 23.7181
R3626 VDD.n275 VDD.n231 23.7181
R3627 VDD.n241 VDD.n235 23.7181
R3628 VDD.n313 VDD.n199 23.7181
R3629 VDD.n187 VDD.n158 22.9652
R3630 VDD.n290 VDD.n218 22.9652
R3631 VDD.n298 VDD.n297 22.9652
R3632 VDD.n308 VDD.n201 22.5887
R3633 VDD.n302 VDD.n301 22.5887
R3634 VDD.n163 VDD.t43 21.2133
R3635 VDD.t14 VDD.n153 21.2133
R3636 VDD.n308 VDD.n307 21.0829
R3637 VDD.n345 VDD.n344 20.3299
R3638 VDD.n356 VDD.n355 20.3299
R3639 VDD.n367 VDD.n366 20.3299
R3640 VDD.n378 VDD.n377 20.3299
R3641 VDD.n389 VDD.n388 20.3299
R3642 VDD.n400 VDD.n399 20.3299
R3643 VDD.n411 VDD.n410 20.3299
R3644 VDD.n422 VDD.n421 20.3299
R3645 VDD.n433 VDD.n432 20.3299
R3646 VDD.n8 VDD.n7 20.3299
R3647 VDD.t186 VDD.t54 20.1418
R3648 VDD.n268 VDD.n252 19.9534
R3649 VDD.n240 VDD.n239 19.9534
R3650 VDD.n301 VDD.n300 18.824
R3651 VDD.n306 VDD.n210 18.4476
R3652 VDD.t43 VDD.n161 17.4699
R3653 VDD.n331 VDD.t14 17.4699
R3654 VDD.n350 VDD.n42 17.3181
R3655 VDD.n361 VDD.n38 17.3181
R3656 VDD.n372 VDD.n34 17.3181
R3657 VDD.n383 VDD.n30 17.3181
R3658 VDD.n394 VDD.n26 17.3181
R3659 VDD.n405 VDD.n22 17.3181
R3660 VDD.n416 VDD.n18 17.3181
R3661 VDD.n427 VDD.n14 17.3181
R3662 VDD.n438 VDD.n3 17.3181
R3663 VDD.n441 VDD.n440 17.3181
R3664 VDD.n303 VDD.n210 16.1887
R3665 VDD.n351 VDD.n350 15.8123
R3666 VDD.n362 VDD.n361 15.8123
R3667 VDD.n373 VDD.n372 15.8123
R3668 VDD.n384 VDD.n383 15.8123
R3669 VDD.n395 VDD.n394 15.8123
R3670 VDD.n406 VDD.n405 15.8123
R3671 VDD.n417 VDD.n416 15.8123
R3672 VDD.n428 VDD.n427 15.8123
R3673 VDD.n438 VDD.n4 15.8123
R3674 VDD.n80 VDD 15.0074
R3675 VDD.n86 VDD 15.0074
R3676 VDD VDD.n54 15.0074
R3677 VDD.n113 VDD 15.0074
R3678 VDD.n144 VDD 15.0074
R3679 VDD.n294 VDD.n218 14.3064
R3680 VDD.n300 VDD.n299 14.3064
R3681 VDD.n299 VDD.n298 14.3064
R3682 VDD.n239 VDD.n238 13.5534
R3683 VDD.n79 VDD.n56 12.8005
R3684 VDD.n75 VDD.n74 12.8005
R3685 VDD.n69 VDD.n59 12.8005
R3686 VDD.n67 VDD.n66 12.8005
R3687 VDD.n87 VDD.n55 12.8005
R3688 VDD.n92 VDD.n91 12.8005
R3689 VDD.n97 VDD.n96 12.8005
R3690 VDD.n102 VDD.n101 12.8005
R3691 VDD.n107 VDD.n106 12.8005
R3692 VDD.n112 VDD.n49 12.8005
R3693 VDD.n145 VDD.n48 12.8005
R3694 VDD.n125 VDD.n124 12.8005
R3695 VDD.n130 VDD.n129 12.8005
R3696 VDD.n135 VDD.n134 12.8005
R3697 VDD.n140 VDD.n116 12.8005
R3698 VDD.n333 VDD.n151 12.8005
R3699 VDD.n170 VDD.n151 12.8005
R3700 VDD.n175 VDD.n167 12.8005
R3701 VDD.n177 VDD.n165 12.8005
R3702 VDD.n181 VDD.n165 12.8005
R3703 VDD.n277 VDD.n230 12.8005
R3704 VDD.n259 VDD.n258 12.8005
R3705 VDD.n275 VDD.n232 12.8005
R3706 VDD.n247 VDD.n246 12.8005
R3707 VDD.n283 VDD.n282 12.8005
R3708 VDD.n294 VDD.n219 12.8005
R3709 VDD.n89 VDD.n47 11.6828
R3710 VDD.n148 VDD.n147 11.6828
R3711 VDD.n271 VDD.n270 10.5417
R3712 VDD.n204 VDD.n203 10.5417
R3713 VDD.n337 VDD 9.79446
R3714 VDD.n79 VDD 9.32654
R3715 VDD.n140 VDD.n139 9.3005
R3716 VDD.n138 VDD.n116 9.3005
R3717 VDD.n137 VDD.n136 9.3005
R3718 VDD.n135 VDD.n117 9.3005
R3719 VDD.n134 VDD.n133 9.3005
R3720 VDD.n132 VDD.n118 9.3005
R3721 VDD.n131 VDD.n130 9.3005
R3722 VDD.n129 VDD.n128 9.3005
R3723 VDD.n127 VDD.n119 9.3005
R3724 VDD.n126 VDD.n125 9.3005
R3725 VDD.n124 VDD.n123 9.3005
R3726 VDD.n122 VDD.n120 9.3005
R3727 VDD.n121 VDD.n48 9.3005
R3728 VDD.n146 VDD.n145 9.3005
R3729 VDD.n112 VDD.n111 9.3005
R3730 VDD.n110 VDD.n49 9.3005
R3731 VDD.n109 VDD.n108 9.3005
R3732 VDD.n107 VDD.n50 9.3005
R3733 VDD.n106 VDD.n105 9.3005
R3734 VDD.n104 VDD.n51 9.3005
R3735 VDD.n103 VDD.n102 9.3005
R3736 VDD.n101 VDD.n100 9.3005
R3737 VDD.n99 VDD.n52 9.3005
R3738 VDD.n98 VDD.n97 9.3005
R3739 VDD.n96 VDD.n95 9.3005
R3740 VDD.n94 VDD.n53 9.3005
R3741 VDD.n93 VDD.n92 9.3005
R3742 VDD.n91 VDD.n90 9.3005
R3743 VDD.n88 VDD.n87 9.3005
R3744 VDD.n63 VDD.n55 9.3005
R3745 VDD.n65 VDD.n64 9.3005
R3746 VDD.n66 VDD.n62 9.3005
R3747 VDD.n67 VDD.n61 9.3005
R3748 VDD.n68 VDD.n60 9.3005
R3749 VDD.n70 VDD.n69 9.3005
R3750 VDD.n71 VDD.n59 9.3005
R3751 VDD.n73 VDD.n72 9.3005
R3752 VDD.n74 VDD.n58 9.3005
R3753 VDD.n75 VDD.n57 9.3005
R3754 VDD.n77 VDD.n76 9.3005
R3755 VDD.n78 VDD.n56 9.3005
R3756 VDD.n238 VDD.n198 9.3005
R3757 VDD.n239 VDD.n237 9.3005
R3758 VDD.n243 VDD.n235 9.3005
R3759 VDD.n246 VDD.n234 9.3005
R3760 VDD.n247 VDD.n233 9.3005
R3761 VDD.n250 VDD.n232 9.3005
R3762 VDD.n275 VDD.n274 9.3005
R3763 VDD.n268 VDD.n267 9.3005
R3764 VDD.n263 VDD.n262 9.3005
R3765 VDD.n260 VDD.n259 9.3005
R3766 VDD.n258 VDD.n257 9.3005
R3767 VDD.n255 VDD.n230 9.3005
R3768 VDD.n278 VDD.n277 9.3005
R3769 VDD.n256 VDD.n254 9.3005
R3770 VDD.n261 VDD.n253 9.3005
R3771 VDD.n265 VDD.n264 9.3005
R3772 VDD.n266 VDD.n252 9.3005
R3773 VDD.n269 VDD.n251 9.3005
R3774 VDD.n272 VDD.n271 9.3005
R3775 VDD.n273 VDD.n231 9.3005
R3776 VDD.n249 VDD.n248 9.3005
R3777 VDD.n245 VDD.n244 9.3005
R3778 VDD.n242 VDD.n241 9.3005
R3779 VDD.n240 VDD.n236 9.3005
R3780 VDD.n314 VDD.n313 9.3005
R3781 VDD.n311 VDD.n310 9.3005
R3782 VDD.n304 VDD.n303 9.3005
R3783 VDD.n300 VDD.n213 9.3005
R3784 VDD.n298 VDD.n215 9.3005
R3785 VDD.n297 VDD.n216 9.3005
R3786 VDD.n222 VDD.n220 9.3005
R3787 VDD.n226 VDD.n219 9.3005
R3788 VDD.n294 VDD.n293 9.3005
R3789 VDD.n291 VDD.n290 9.3005
R3790 VDD.n287 VDD.n286 9.3005
R3791 VDD.n283 VDD.n229 9.3005
R3792 VDD.n282 VDD.n281 9.3005
R3793 VDD.n285 VDD.n284 9.3005
R3794 VDD.n292 VDD.n218 9.3005
R3795 VDD.n225 VDD.n224 9.3005
R3796 VDD.n299 VDD.n214 9.3005
R3797 VDD.n301 VDD.n211 9.3005
R3798 VDD.n306 VDD.n305 9.3005
R3799 VDD.n307 VDD.n209 9.3005
R3800 VDD.n309 VDD.n308 9.3005
R3801 VDD.n206 VDD.n200 9.3005
R3802 VDD.n205 VDD.n204 9.3005
R3803 VDD.n202 VDD.n199 9.3005
R3804 VDD.n326 VDD.n325 9.3005
R3805 VDD.n329 VDD.n194 9.3005
R3806 VDD.n185 VDD.n184 9.3005
R3807 VDD.n181 VDD.n180 9.3005
R3808 VDD.n179 VDD.n165 9.3005
R3809 VDD.n178 VDD.n177 9.3005
R3810 VDD.n175 VDD.n174 9.3005
R3811 VDD.n173 VDD.n167 9.3005
R3812 VDD.n170 VDD.n169 9.3005
R3813 VDD.n168 VDD.n151 9.3005
R3814 VDD.n334 VDD.n333 9.3005
R3815 VDD.n172 VDD.n171 9.3005
R3816 VDD.n176 VDD.n166 9.3005
R3817 VDD.n182 VDD.n159 9.3005
R3818 VDD.n187 VDD.n186 9.3005
R3819 VDD.n188 VDD.n157 9.3005
R3820 VDD.n192 VDD.n191 9.3005
R3821 VDD.n193 VDD.n156 9.3005
R3822 VDD.n328 VDD.n327 9.3005
R3823 VDD.n323 VDD.n196 9.3005
R3824 VDD.n322 VDD.n321 9.3005
R3825 VDD.n320 VDD.n197 9.3005
R3826 VDD.n319 VDD.n318 9.3005
R3827 VDD.n440 VDD.n0 9.3005
R3828 VDD.n7 VDD.n6 9.3005
R3829 VDD.n11 VDD.n4 9.3005
R3830 VDD.n438 VDD.n437 9.3005
R3831 VDD.n433 VDD.n12 9.3005
R3832 VDD.n429 VDD.n428 9.3005
R3833 VDD.n427 VDD.n426 9.3005
R3834 VDD.n422 VDD.n16 9.3005
R3835 VDD.n418 VDD.n417 9.3005
R3836 VDD.n416 VDD.n415 9.3005
R3837 VDD.n411 VDD.n20 9.3005
R3838 VDD.n407 VDD.n406 9.3005
R3839 VDD.n405 VDD.n404 9.3005
R3840 VDD.n400 VDD.n24 9.3005
R3841 VDD.n396 VDD.n395 9.3005
R3842 VDD.n394 VDD.n393 9.3005
R3843 VDD.n389 VDD.n28 9.3005
R3844 VDD.n385 VDD.n384 9.3005
R3845 VDD.n383 VDD.n382 9.3005
R3846 VDD.n378 VDD.n32 9.3005
R3847 VDD.n374 VDD.n373 9.3005
R3848 VDD.n372 VDD.n371 9.3005
R3849 VDD.n367 VDD.n36 9.3005
R3850 VDD.n363 VDD.n362 9.3005
R3851 VDD.n361 VDD.n360 9.3005
R3852 VDD.n356 VDD.n40 9.3005
R3853 VDD.n352 VDD.n351 9.3005
R3854 VDD.n350 VDD.n349 9.3005
R3855 VDD.n345 VDD.n44 9.3005
R3856 VDD.n341 VDD.n340 9.3005
R3857 VDD.n342 VDD.n45 9.3005
R3858 VDD.n344 VDD.n343 9.3005
R3859 VDD.n347 VDD.n346 9.3005
R3860 VDD.n348 VDD.n42 9.3005
R3861 VDD.n353 VDD.n41 9.3005
R3862 VDD.n355 VDD.n354 9.3005
R3863 VDD.n358 VDD.n357 9.3005
R3864 VDD.n359 VDD.n38 9.3005
R3865 VDD.n364 VDD.n37 9.3005
R3866 VDD.n366 VDD.n365 9.3005
R3867 VDD.n369 VDD.n368 9.3005
R3868 VDD.n370 VDD.n34 9.3005
R3869 VDD.n375 VDD.n33 9.3005
R3870 VDD.n377 VDD.n376 9.3005
R3871 VDD.n380 VDD.n379 9.3005
R3872 VDD.n381 VDD.n30 9.3005
R3873 VDD.n386 VDD.n29 9.3005
R3874 VDD.n388 VDD.n387 9.3005
R3875 VDD.n391 VDD.n390 9.3005
R3876 VDD.n392 VDD.n26 9.3005
R3877 VDD.n397 VDD.n25 9.3005
R3878 VDD.n399 VDD.n398 9.3005
R3879 VDD.n402 VDD.n401 9.3005
R3880 VDD.n403 VDD.n22 9.3005
R3881 VDD.n408 VDD.n21 9.3005
R3882 VDD.n410 VDD.n409 9.3005
R3883 VDD.n413 VDD.n412 9.3005
R3884 VDD.n414 VDD.n18 9.3005
R3885 VDD.n419 VDD.n17 9.3005
R3886 VDD.n421 VDD.n420 9.3005
R3887 VDD.n424 VDD.n423 9.3005
R3888 VDD.n425 VDD.n14 9.3005
R3889 VDD.n430 VDD.n13 9.3005
R3890 VDD.n432 VDD.n431 9.3005
R3891 VDD.n435 VDD.n434 9.3005
R3892 VDD.n436 VDD.n3 9.3005
R3893 VDD.n10 VDD.n9 9.3005
R3894 VDD.n8 VDD.n5 9.3005
R3895 VDD.n2 VDD.n1 9.3005
R3896 VDD.n442 VDD.n441 9.3005
R3897 VDD.n189 VDD.n188 8.28285
R3898 VDD.n328 VDD.n195 8.28285
R3899 VDD.n270 VDD.n269 8.28285
R3900 VDD.n203 VDD.n200 8.28285
R3901 VDD.n141 VDD 7.34877
R3902 VDD.t171 VDD.t4 6.71428
R3903 VDD.t31 VDD.t184 6.71428
R3904 VDD.t47 VDD.t188 6.71428
R3905 VDD.t163 VDD.t84 6.71428
R3906 VDD.n150 VDD.n47 6.09998
R3907 VDD.n336 VDD.n335 4.33704
R3908 VDD VDD.n46 4.10787
R3909 VDD.n315 VDD.n198 3.76683
R3910 VDD.n287 VDD.n228 3.76521
R3911 VDD.n223 VDD.n222 3.76521
R3912 VDD.n279 VDD 3.09034
R3913 VDD VDD.n280 3.09034
R3914 VDD.n335 VDD 3.09034
R3915 VDD.n315 VDD.n314 2.89503
R3916 VDD.n317 VDD.n316 2.89503
R3917 VDD.n150 VDD.n149 2.34946
R3918 VDD.n339 VDD.n338 2.34946
R3919 VDD VDD.n46 2.27784
R3920 VDD.n338 VDD.n337 2.24112
R3921 VDD.n339 VDD.n46 2.16789
R3922 VDD.n149 VDD.n148 1.91476
R3923 VDD.n337 VDD.n336 1.82316
R3924 VDD.n338 VDD.n150 1.73404
R3925 VDD.n184 VDD.n183 1.50638
R3926 VDD.n184 VDD.n158 1.12991
R3927 VDD.n288 VDD.n287 1.12991
R3928 VDD.n311 VDD.n201 1.12991
R3929 VDD.n303 VDD.n302 1.12991
R3930 VDD.n222 VDD.n217 1.12991
R3931 VDD.n148 VDD.n47 1.12238
R3932 VDD.n316 VDD.n315 0.872295
R3933 VDD.n280 VDD.n279 0.872295
R3934 VDD VDD.n339 0.647576
R3935 VDD.n149 VDD.n0 0.643669
R3936 VDD.n335 VDD 0.462038
R3937 VDD.n280 VDD 0.410756
R3938 VDD.n191 VDD.n189 0.376971
R3939 VDD.n325 VDD.n195 0.376971
R3940 VDD.n290 VDD.n289 0.376971
R3941 VDD.n336 VDD 0.302844
R3942 VDD.n316 VDD 0.229667
R3943 VDD.n78 VDD.n77 0.120292
R3944 VDD.n77 VDD.n57 0.120292
R3945 VDD.n72 VDD.n58 0.120292
R3946 VDD.n72 VDD.n71 0.120292
R3947 VDD.n70 VDD.n60 0.120292
R3948 VDD.n61 VDD.n60 0.120292
R3949 VDD.n64 VDD.n62 0.120292
R3950 VDD.n64 VDD.n63 0.120292
R3951 VDD.n94 VDD.n93 0.120292
R3952 VDD.n95 VDD.n94 0.120292
R3953 VDD.n99 VDD.n98 0.120292
R3954 VDD.n100 VDD.n99 0.120292
R3955 VDD.n104 VDD.n103 0.120292
R3956 VDD.n105 VDD.n104 0.120292
R3957 VDD.n109 VDD.n50 0.120292
R3958 VDD.n110 VDD.n109 0.120292
R3959 VDD.n122 VDD.n121 0.120292
R3960 VDD.n123 VDD.n122 0.120292
R3961 VDD.n127 VDD.n126 0.120292
R3962 VDD.n128 VDD.n127 0.120292
R3963 VDD.n132 VDD.n131 0.120292
R3964 VDD.n133 VDD.n132 0.120292
R3965 VDD.n137 VDD.n117 0.120292
R3966 VDD.n138 VDD.n137 0.120292
R3967 VDD.n237 VDD.n236 0.120292
R3968 VDD.n242 VDD.n236 0.120292
R3969 VDD.n244 VDD.n243 0.120292
R3970 VDD.n244 VDD.n234 0.120292
R3971 VDD.n249 VDD.n233 0.120292
R3972 VDD.n250 VDD.n249 0.120292
R3973 VDD.n273 VDD.n272 0.120292
R3974 VDD.n272 VDD.n251 0.120292
R3975 VDD.n267 VDD.n266 0.120292
R3976 VDD.n266 VDD.n265 0.120292
R3977 VDD.n262 VDD.n261 0.120292
R3978 VDD.n261 VDD.n260 0.120292
R3979 VDD.n257 VDD.n256 0.120292
R3980 VDD.n256 VDD.n255 0.120292
R3981 VDD.n205 VDD.n202 0.120292
R3982 VDD.n206 VDD.n205 0.120292
R3983 VDD.n305 VDD.n209 0.120292
R3984 VDD.n305 VDD.n304 0.120292
R3985 VDD.n213 VDD.n211 0.120292
R3986 VDD.n214 VDD.n213 0.120292
R3987 VDD.n225 VDD.n220 0.120292
R3988 VDD.n226 VDD.n225 0.120292
R3989 VDD.n292 VDD.n291 0.120292
R3990 VDD.n286 VDD.n285 0.120292
R3991 VDD.n285 VDD.n229 0.120292
R3992 VDD.n320 VDD.n319 0.120292
R3993 VDD.n321 VDD.n320 0.120292
R3994 VDD.n326 VDD.n196 0.120292
R3995 VDD.n327 VDD.n326 0.120292
R3996 VDD.n193 VDD.n192 0.120292
R3997 VDD.n192 VDD.n157 0.120292
R3998 VDD.n185 VDD.n159 0.120292
R3999 VDD.n180 VDD.n159 0.120292
R4000 VDD.n178 VDD.n166 0.120292
R4001 VDD.n174 VDD.n166 0.120292
R4002 VDD.n173 VDD.n172 0.120292
R4003 VDD.n172 VDD.n169 0.120292
R4004 VDD.n90 VDD 0.11899
R4005 VDD VDD.n146 0.11899
R4006 VDD.n319 VDD 0.109875
R4007 VDD VDD.n196 0.104667
R4008 VDD.n147 VDD 0.09425
R4009 VDD.n89 VDD 0.078625
R4010 VDD.n442 VDD.n1 0.072375
R4011 VDD.n6 VDD.n1 0.072375
R4012 VDD.n10 VDD.n5 0.072375
R4013 VDD.n11 VDD.n10 0.072375
R4014 VDD.n436 VDD.n435 0.072375
R4015 VDD.n435 VDD.n12 0.072375
R4016 VDD.n431 VDD.n430 0.072375
R4017 VDD.n430 VDD.n429 0.072375
R4018 VDD.n425 VDD.n424 0.072375
R4019 VDD.n424 VDD.n16 0.072375
R4020 VDD.n420 VDD.n419 0.072375
R4021 VDD.n419 VDD.n418 0.072375
R4022 VDD.n414 VDD.n413 0.072375
R4023 VDD.n413 VDD.n20 0.072375
R4024 VDD.n409 VDD.n408 0.072375
R4025 VDD.n408 VDD.n407 0.072375
R4026 VDD.n403 VDD.n402 0.072375
R4027 VDD.n402 VDD.n24 0.072375
R4028 VDD.n398 VDD.n397 0.072375
R4029 VDD.n397 VDD.n396 0.072375
R4030 VDD.n392 VDD.n391 0.072375
R4031 VDD.n391 VDD.n28 0.072375
R4032 VDD.n387 VDD.n386 0.072375
R4033 VDD.n386 VDD.n385 0.072375
R4034 VDD.n381 VDD.n380 0.072375
R4035 VDD.n380 VDD.n32 0.072375
R4036 VDD.n376 VDD.n375 0.072375
R4037 VDD.n375 VDD.n374 0.072375
R4038 VDD.n370 VDD.n369 0.072375
R4039 VDD.n369 VDD.n36 0.072375
R4040 VDD.n365 VDD.n364 0.072375
R4041 VDD.n364 VDD.n363 0.072375
R4042 VDD.n359 VDD.n358 0.072375
R4043 VDD.n358 VDD.n40 0.072375
R4044 VDD.n354 VDD.n353 0.072375
R4045 VDD.n353 VDD.n352 0.072375
R4046 VDD.n348 VDD.n347 0.072375
R4047 VDD.n347 VDD.n44 0.072375
R4048 VDD.n343 VDD.n342 0.072375
R4049 VDD.n342 VDD.n341 0.072375
R4050 VDD VDD.n78 0.0603958
R4051 VDD.n58 VDD 0.0603958
R4052 VDD VDD.n70 0.0603958
R4053 VDD.n62 VDD 0.0603958
R4054 VDD.n88 VDD 0.0603958
R4055 VDD.n93 VDD 0.0603958
R4056 VDD.n98 VDD 0.0603958
R4057 VDD.n103 VDD 0.0603958
R4058 VDD VDD.n50 0.0603958
R4059 VDD.n111 VDD 0.0603958
R4060 VDD.n121 VDD 0.0603958
R4061 VDD.n126 VDD 0.0603958
R4062 VDD.n131 VDD 0.0603958
R4063 VDD VDD.n117 0.0603958
R4064 VDD.n139 VDD 0.0603958
R4065 VDD.n237 VDD 0.0603958
R4066 VDD.n243 VDD 0.0603958
R4067 VDD VDD.n233 0.0603958
R4068 VDD.n274 VDD 0.0603958
R4069 VDD VDD.n273 0.0603958
R4070 VDD.n267 VDD 0.0603958
R4071 VDD.n262 VDD 0.0603958
R4072 VDD.n257 VDD 0.0603958
R4073 VDD.n278 VDD 0.0603958
R4074 VDD.n202 VDD 0.0603958
R4075 VDD.n310 VDD 0.0603958
R4076 VDD VDD.n309 0.0603958
R4077 VDD.n209 VDD 0.0603958
R4078 VDD.n211 VDD 0.0603958
R4079 VDD.n215 VDD 0.0603958
R4080 VDD.n216 VDD 0.0603958
R4081 VDD.n220 VDD 0.0603958
R4082 VDD.n293 VDD 0.0603958
R4083 VDD VDD.n292 0.0603958
R4084 VDD.n286 VDD 0.0603958
R4085 VDD.n281 VDD 0.0603958
R4086 VDD VDD.n194 0.0603958
R4087 VDD VDD.n193 0.0603958
R4088 VDD.n186 VDD 0.0603958
R4089 VDD VDD.n185 0.0603958
R4090 VDD VDD.n179 0.0603958
R4091 VDD VDD.n178 0.0603958
R4092 VDD VDD.n173 0.0603958
R4093 VDD VDD.n168 0.0603958
R4094 VDD.n334 VDD 0.0603958
R4095 VDD VDD.n89 0.0408646
R4096 VDD.n274 VDD 0.0382604
R4097 VDD.n279 VDD 0.0365577
R4098 VDD VDD.n442 0.0364375
R4099 VDD VDD.n5 0.0364375
R4100 VDD.n437 VDD 0.0364375
R4101 VDD VDD.n436 0.0364375
R4102 VDD.n431 VDD 0.0364375
R4103 VDD.n426 VDD 0.0364375
R4104 VDD VDD.n425 0.0364375
R4105 VDD.n420 VDD 0.0364375
R4106 VDD.n415 VDD 0.0364375
R4107 VDD VDD.n414 0.0364375
R4108 VDD.n409 VDD 0.0364375
R4109 VDD.n404 VDD 0.0364375
R4110 VDD VDD.n403 0.0364375
R4111 VDD.n398 VDD 0.0364375
R4112 VDD.n393 VDD 0.0364375
R4113 VDD VDD.n392 0.0364375
R4114 VDD.n387 VDD 0.0364375
R4115 VDD.n382 VDD 0.0364375
R4116 VDD VDD.n381 0.0364375
R4117 VDD.n376 VDD 0.0364375
R4118 VDD.n371 VDD 0.0364375
R4119 VDD VDD.n370 0.0364375
R4120 VDD.n365 VDD 0.0364375
R4121 VDD.n360 VDD 0.0364375
R4122 VDD VDD.n359 0.0364375
R4123 VDD.n354 VDD 0.0364375
R4124 VDD.n349 VDD 0.0364375
R4125 VDD VDD.n348 0.0364375
R4126 VDD.n343 VDD 0.0364375
R4127 VDD VDD.n198 0.03175
R4128 VDD VDD.n278 0.03175
R4129 VDD.n314 VDD 0.03175
R4130 VDD.n310 VDD 0.03175
R4131 VDD.n309 VDD 0.03175
R4132 VDD VDD.n216 0.03175
R4133 VDD.n293 VDD 0.03175
R4134 VDD.n281 VDD 0.03175
R4135 VDD.n179 VDD 0.03175
R4136 VDD.n168 VDD 0.03175
R4137 VDD VDD.n334 0.03175
R4138 VDD VDD.n88 0.0265417
R4139 VDD.n90 VDD 0.0265417
R4140 VDD.n111 VDD 0.0265417
R4141 VDD.n146 VDD 0.0265417
R4142 VDD.n139 VDD 0.0265417
R4143 VDD.n147 VDD 0.0252396
R4144 VDD VDD.n57 0.0239375
R4145 VDD.n71 VDD 0.0239375
R4146 VDD VDD.n61 0.0239375
R4147 VDD.n63 VDD 0.0239375
R4148 VDD.n95 VDD 0.0239375
R4149 VDD.n100 VDD 0.0239375
R4150 VDD.n105 VDD 0.0239375
R4151 VDD VDD.n110 0.0239375
R4152 VDD.n123 VDD 0.0239375
R4153 VDD.n128 VDD 0.0239375
R4154 VDD.n133 VDD 0.0239375
R4155 VDD VDD.n138 0.0239375
R4156 VDD.n234 VDD 0.0239375
R4157 VDD VDD.n250 0.0239375
R4158 VDD.n260 VDD 0.0239375
R4159 VDD.n255 VDD 0.0239375
R4160 VDD VDD.n214 0.0239375
R4161 VDD.n291 VDD 0.0239375
R4162 VDD.n174 VDD 0.0239375
R4163 VDD.n169 VDD 0.0239375
R4164 VDD VDD.n251 0.0226354
R4165 VDD VDD.n206 0.0226354
R4166 VDD.n327 VDD 0.0226354
R4167 VDD VDD.n157 0.0226354
R4168 VDD VDD.n242 0.0213333
R4169 VDD.n265 VDD 0.0213333
R4170 VDD.n304 VDD 0.0213333
R4171 VDD VDD.n215 0.0213333
R4172 VDD VDD.n226 0.0213333
R4173 VDD VDD.n229 0.0213333
R4174 VDD.n194 VDD 0.0213333
R4175 VDD.n186 VDD 0.0213333
R4176 VDD.n180 VDD 0.0213333
R4177 VDD VDD.n0 0.01925
R4178 VDD.n437 VDD 0.01925
R4179 VDD.n426 VDD 0.01925
R4180 VDD.n415 VDD 0.01925
R4181 VDD.n404 VDD 0.01925
R4182 VDD.n393 VDD 0.01925
R4183 VDD.n382 VDD 0.01925
R4184 VDD.n371 VDD 0.01925
R4185 VDD.n360 VDD 0.01925
R4186 VDD.n349 VDD 0.01925
R4187 VDD.n321 VDD 0.016125
R4188 VDD.n6 VDD 0.0137813
R4189 VDD VDD.n11 0.0137813
R4190 VDD VDD.n12 0.0137813
R4191 VDD.n429 VDD 0.0137813
R4192 VDD VDD.n16 0.0137813
R4193 VDD.n418 VDD 0.0137813
R4194 VDD VDD.n20 0.0137813
R4195 VDD.n407 VDD 0.0137813
R4196 VDD VDD.n24 0.0137813
R4197 VDD.n396 VDD 0.0137813
R4198 VDD VDD.n28 0.0137813
R4199 VDD.n385 VDD 0.0137813
R4200 VDD VDD.n32 0.0137813
R4201 VDD.n374 VDD 0.0137813
R4202 VDD VDD.n36 0.0137813
R4203 VDD.n363 VDD 0.0137813
R4204 VDD VDD.n40 0.0137813
R4205 VDD.n352 VDD 0.0137813
R4206 VDD VDD.n44 0.0137813
R4207 VDD.n341 VDD 0.0137813
R4208 VDD.n317 VDD 0.0109167
R4209 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t0 230.71
R4210 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t5 230.576
R4211 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t4 230.155
R4212 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t7 230.155
R4213 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n7 205.28
R4214 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t9 158.275
R4215 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t6 157.856
R4216 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t8 157.856
R4217 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n8 153.067
R4218 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n2 152
R4219 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n0 152
R4220 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t1 135.947
R4221 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n11 67.4857
R4222 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n10 44.0818
R4223 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n6 33.5064
R4224 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t2 26.5955
R4225 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t3 26.5955
R4226 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n5 23.9017
R4227 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n9 19.3316
R4228 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 16.4149
R4229 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n1 12.2559
R4230 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n3 11.0199
R4231 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 5.6005
R4232 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n4 5.0505
R4233 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 2.10199
R4234 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 2.10199
R4235 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.05675
R4236 top_segment_3_0.b[5].n2 top_segment_3_0.b[5].n1 863.124
R4237 top_segment_3_0.b[5].n1 top_segment_3_0.b[5].n0 585
R4238 top_segment_3_0.b[5] top_segment_3_0.b[5].t0 495.469
R4239 top_segment_3_0.b[5].n6 top_segment_3_0.b[5].t4 217.555
R4240 top_segment_3_0.b[5].n6 top_segment_3_0.b[5].t6 216.893
R4241 top_segment_3_0.b[5].n5 top_segment_3_0.b[5].t5 216.893
R4242 top_segment_3_0.b[5].n4 top_segment_3_0.b[5].t2 216.893
R4243 top_segment_3_0.b[5].n8 top_segment_3_0.b[5].t3 212.393
R4244 top_segment_3_0.b[5].n3 top_segment_3_0.b[5].t1 141.189
R4245 top_segment_3_0.b[5].n1 top_segment_3_0.b[5].t0 140.738
R4246 top_segment_3_0.b[5] top_segment_3_0.b[5].n8 90.6776
R4247 top_segment_3_0.b[5].n9 top_segment_3_0.b[5] 14.3755
R4248 top_segment_3_0.b[5].n2 top_segment_3_0.b[5] 11.6369
R4249 top_segment_3_0.b[5].n0 top_segment_3_0.b[5] 10.1408
R4250 top_segment_3_0.b[5] top_segment_3_0.b[5].n9 8.53383
R4251 top_segment_3_0.b[5] top_segment_3_0.b[5].n3 7.94225
R4252 top_segment_3_0.b[5].n3 top_segment_3_0.b[5] 6.14988
R4253 top_segment_3_0.b[5].n9 top_segment_3_0.b[5] 5.81868
R4254 top_segment_3_0.b[5].n8 top_segment_3_0.b[5].n7 4.5005
R4255 top_segment_3_0.b[5].n0 top_segment_3_0.b[5] 2.16154
R4256 top_segment_3_0.b[5] top_segment_3_0.b[5].n2 0.665435
R4257 top_segment_3_0.b[5].n5 top_segment_3_0.b[5].n4 0.663962
R4258 top_segment_3_0.b[5].n7 top_segment_3_0.b[5].n5 0.663962
R4259 top_segment_3_0.b[5].n7 top_segment_3_0.b[5].n6 0.663962
R4260 top_segment_3_0.b[5].n4 top_segment_3_0.b[5] 0.325019
R4261 a_15695_17684.n0 a_15695_17684.t2 670.792
R4262 a_15695_17684.n0 a_15695_17684.t1 666.963
R4263 a_15695_17684.t0 a_15695_17684.n0 665.304
R4264 a_13061_17684.n0 a_13061_17684.t2 671.227
R4265 a_13061_17684.n0 a_13061_17684.t1 665.75
R4266 a_13061_17684.t0 a_13061_17684.n0 665.298
R4267 VDDH.n31 VDDH.n18 5941.3
R4268 VDDH.n673 VDDH.n31 5941.3
R4269 VDDH.n692 VDDH.n18 5939.4
R4270 VDDH.n7 VDDH.n5 5352.3
R4271 VDDH.n433 VDDH.n429 4436.17
R4272 VDDH.n433 VDDH.n430 4436.17
R4273 VDDH.n435 VDDH.n429 4436.17
R4274 VDDH.n435 VDDH.n430 4436.17
R4275 VDDH.n676 VDDH.n675 4157.2
R4276 VDDH.n281 VDDH.n277 3638.5
R4277 VDDH.n300 VDDH.n277 3638.5
R4278 VDDH.n342 VDDH.n317 3298.14
R4279 VDDH.n345 VDDH.n317 3296.17
R4280 VDDH.n345 VDDH.n318 2942.38
R4281 VDDH.n352 VDDH.n310 2942.38
R4282 VDDH.n354 VDDH.n305 2942.38
R4283 VDDH.n355 VDDH.n305 2942.38
R4284 VDDH.n351 VDDH.n310 2942.38
R4285 VDDH.n342 VDDH.n319 2940.41
R4286 VDDH.n677 VDDH.n676 2855.7
R4287 VDDH.n62 VDDH.n33 2705.6
R4288 VDDH.n297 VDDH.n280 2692.3
R4289 VDDH.n517 VDDH.n378 2671.14
R4290 VDDH.n519 VDDH.n378 2671.14
R4291 VDDH.n519 VDDH.n516 2671.14
R4292 VDDH.n517 VDDH.n516 2671.14
R4293 VDDH.n441 VDDH.n413 2671.14
R4294 VDDH.n441 VDDH.n414 2671.14
R4295 VDDH.n443 VDDH.n413 2671.14
R4296 VDDH.n443 VDDH.n414 2671.14
R4297 VDDH.n422 VDDH.n418 2671.14
R4298 VDDH.n424 VDDH.n418 2671.14
R4299 VDDH.n424 VDDH.n420 2671.14
R4300 VDDH.n422 VDDH.n420 2671.14
R4301 VDDH.n508 VDDH.n383 2671.14
R4302 VDDH.n508 VDDH.n384 2671.14
R4303 VDDH.n510 VDDH.n383 2671.14
R4304 VDDH.n510 VDDH.n384 2671.14
R4305 VDDH.n501 VDDH.n388 2671.14
R4306 VDDH.n501 VDDH.n389 2671.14
R4307 VDDH.n499 VDDH.n389 2671.14
R4308 VDDH.n499 VDDH.n388 2671.14
R4309 VDDH.n454 VDDH.n448 2671.14
R4310 VDDH.n454 VDDH.n450 2671.14
R4311 VDDH.n452 VDDH.n450 2671.14
R4312 VDDH.n452 VDDH.n448 2671.14
R4313 VDDH.n461 VDDH.n407 2671.14
R4314 VDDH.n461 VDDH.n408 2671.14
R4315 VDDH.n463 VDDH.n408 2671.14
R4316 VDDH.n463 VDDH.n407 2671.14
R4317 VDDH.n494 VDDH.n394 2671.14
R4318 VDDH.n494 VDDH.n395 2671.14
R4319 VDDH.n492 VDDH.n395 2671.14
R4320 VDDH.n492 VDDH.n394 2671.14
R4321 VDDH.n483 VDDH.n399 2671.14
R4322 VDDH.n483 VDDH.n400 2671.14
R4323 VDDH.n485 VDDH.n400 2671.14
R4324 VDDH.n485 VDDH.n399 2671.14
R4325 VDDH.n474 VDDH.n467 2671.14
R4326 VDDH.n474 VDDH.n468 2671.14
R4327 VDDH.n472 VDDH.n468 2671.14
R4328 VDDH.n472 VDDH.n467 2671.14
R4329 VDDH.n353 VDDH.n352 2588.59
R4330 VDDH.n354 VDDH.n353 2588.59
R4331 VDDH.n351 VDDH.n308 2588.59
R4332 VDDH.n355 VDDH.n308 2588.59
R4333 VDDH.n297 VDDH.n278 2513.7
R4334 VDDH.n14 VDDH.n7 2129.9
R4335 VDDH.n695 VDDH.n14 2069.1
R4336 VDDH.n278 VDDH.n5 1983.6
R4337 VDDH.n627 VDDH.n81 1881
R4338 VDDH.n627 VDDH.n82 1881
R4339 VDDH.n596 VDDH.n82 1881
R4340 VDDH.n596 VDDH.n148 1881
R4341 VDDH.n576 VDDH.n148 1881
R4342 VDDH.n576 VDDH.n166 1881
R4343 VDDH.n553 VDDH.n166 1881
R4344 VDDH.n553 VDDH.n231 1881
R4345 VDDH.n539 VDDH.n231 1881
R4346 VDDH.n539 VDDH.n538 1881
R4347 VDDH.n333 VDDH.n327 1857.41
R4348 VDDH.n332 VDDH.n327 1857.41
R4349 VDDH.n674 VDDH.n13 1506.3
R4350 VDDH.n337 VDDH.n318 1503.62
R4351 VDDH.n337 VDDH.n325 1503.62
R4352 VDDH.n333 VDDH.n325 1503.62
R4353 VDDH.n338 VDDH.n319 1503.62
R4354 VDDH.n338 VDDH.n322 1503.62
R4355 VDDH.n332 VDDH.n322 1503.62
R4356 VDDH.n675 VDDH.n19 1407.9
R4357 VDDH.n685 VDDH.n30 1182.12
R4358 VDDH.n30 VDDH.n20 1182.12
R4359 VDDH.n691 VDDH.n20 1181.74
R4360 VDDH.n281 VDDH.n280 986.101
R4361 VDDH.n300 VDDH.n278 986.101
R4362 VDDH.n426 VDDH.n415 883.577
R4363 VDDH.n445 VDDH.n411 883.577
R4364 VDDH.n432 VDDH.n416 854.212
R4365 VDDH.n432 VDDH.n431 854.212
R4366 VDDH.n684 VDDH.n683 823.718
R4367 VDDH.n436 VDDH.n428 781.929
R4368 VDDH.n437 VDDH.n436 781.929
R4369 VDDH.t74 VDDH.t40 740.356
R4370 VDDH.n703 VDDH.n702 725.46
R4371 VDDH.n364 VDDH.n363 720.942
R4372 VDDH.n364 VDDH.n276 720.942
R4373 VDDH.n675 VDDH.n674 720.101
R4374 VDDH.n523 VDDH.t224 667.769
R4375 VDDH.n341 VDDH.n315 636.236
R4376 VDDH.t122 VDDH.t240 583.548
R4377 VDDH.t187 VDDH.t197 583.548
R4378 VDDH.t92 VDDH.t186 583.548
R4379 VDDH.n358 VDDH.n304 568.095
R4380 VDDH.n684 VDDH.n680 564.33
R4381 VDDH.n346 VDDH.n316 563.577
R4382 VDDH.n341 VDDH.n340 563.201
R4383 VDDH.t209 VDDH.t69 552.236
R4384 VDDH.n667 VDDH.n34 536.095
R4385 VDDH.n63 VDDH.n34 536.095
R4386 VDDH.n296 VDDH.n283 533.46
R4387 VDDH.t29 VDDH.t164 523.162
R4388 VDDH.t274 VDDH.t221 523.162
R4389 VDDH.t75 VDDH.t9 523.162
R4390 VDDH.t2 VDDH.t27 523.162
R4391 VDDH.t207 VDDH.t305 523.162
R4392 VDDH.t310 VDDH.t175 523.162
R4393 VDDH.n421 VDDH.n417 516.141
R4394 VDDH.n507 VDDH.n381 516.141
R4395 VDDH.n460 VDDH.n406 516.141
R4396 VDDH.n464 VDDH.n406 516.141
R4397 VDDH.n471 VDDH.n469 516.141
R4398 VDDH.n521 VDDH.n377 516.141
R4399 VDDH.n521 VDDH.n520 516.141
R4400 VDDH.n16 VDDH.n14 513
R4401 VDDH.n674 VDDH.n16 511.101
R4402 VDDH.n541 VDDH.t301 499.882
R4403 VDDH.n263 VDDH.t272 499.882
R4404 VDDH.n230 VDDH.t0 499.882
R4405 VDDH.n536 VDDH.t65 499.882
R4406 VDDH.n313 VDDH.n312 495.812
R4407 VDDH.n312 VDDH.n304 495.812
R4408 VDDH.n350 VDDH.n349 495.812
R4409 VDDH.n350 VDDH.n307 495.812
R4410 VDDH.n356 VDDH.n307 495.812
R4411 VDDH.n357 VDDH.n356 495.812
R4412 VDDH VDDH.n313 490.166
R4413 VDDH.n677 VDDH.n13 489.267
R4414 VDDH.n295 VDDH.n4 486.776
R4415 VDDH.n695 VDDH.n13 486.401
R4416 VDDH.t275 VDDH.t111 475
R4417 VDDH.t165 VDDH.t189 475
R4418 VDDH.t190 VDDH.t188 475
R4419 VDDH.t37 VDDH.t43 475
R4420 VDDH.t43 VDDH.t48 475
R4421 VDDH.t176 VDDH.t284 475
R4422 VDDH.t277 VDDH.t237 475
R4423 VDDH.t56 VDDH.t280 475
R4424 VDDH.n440 VDDH.n415 443.86
R4425 VDDH.n419 VDDH.n409 443.86
R4426 VDDH.n419 VDDH.n411 443.86
R4427 VDDH.n445 VDDH.n444 443.86
R4428 VDDH.n444 VDDH.n386 443.86
R4429 VDDH.n455 VDDH.n447 443.86
R4430 VDDH.n502 VDDH.n387 443.86
R4431 VDDH.n507 VDDH.n506 443.86
R4432 VDDH.n465 VDDH.n464 443.86
R4433 VDDH.n451 VDDH.n404 443.86
R4434 VDDH.n451 VDDH.n401 443.86
R4435 VDDH.n498 VDDH.n391 443.86
R4436 VDDH.n498 VDDH.n497 443.86
R4437 VDDH.n511 VDDH.n382 443.86
R4438 VDDH.n512 VDDH.n511 443.86
R4439 VDDH.n471 VDDH.n470 443.86
R4440 VDDH.n486 VDDH.n398 443.86
R4441 VDDH.n487 VDDH.n486 443.86
R4442 VDDH.n491 VDDH.n488 443.86
R4443 VDDH.n491 VDDH.n490 443.86
R4444 VDDH.n520 VDDH.n379 443.86
R4445 VDDH.t94 VDDH.t108 431.25
R4446 VDDH.t117 VDDH.t94 431.25
R4447 VDDH.t119 VDDH.t117 431.25
R4448 VDDH.t93 VDDH.t116 431.25
R4449 VDDH.t116 VDDH.t95 431.25
R4450 VDDH.t95 VDDH.t96 431.25
R4451 VDDH.t113 VDDH.t112 431.25
R4452 VDDH.t267 VDDH.t113 431.25
R4453 VDDH.t111 VDDH.t267 431.25
R4454 VDDH.t276 VDDH.t275 431.25
R4455 VDDH.t166 VDDH.t276 431.25
R4456 VDDH.t189 VDDH.t190 431.25
R4457 VDDH.t188 VDDH.t37 431.25
R4458 VDDH.t239 VDDH.t70 431.25
R4459 VDDH.t73 VDDH.t239 431.25
R4460 VDDH.t98 VDDH.t73 431.25
R4461 VDDH.t71 VDDH.t72 431.25
R4462 VDDH.t72 VDDH.t97 431.25
R4463 VDDH.t97 VDDH.t238 431.25
R4464 VDDH.t99 VDDH.t282 431.25
R4465 VDDH.t103 VDDH.t99 431.25
R4466 VDDH.t104 VDDH.t103 431.25
R4467 VDDH.t102 VDDH.t91 431.25
R4468 VDDH.t285 VDDH.t102 431.25
R4469 VDDH.t283 VDDH.t285 431.25
R4470 VDDH.t105 VDDH.t107 431.25
R4471 VDDH.t106 VDDH.t105 431.25
R4472 VDDH.t121 VDDH.t106 431.25
R4473 VDDH.t110 VDDH.t118 431.25
R4474 VDDH.t118 VDDH.t120 431.25
R4475 VDDH.t120 VDDH.t109 431.25
R4476 VDDH.t126 VDDH.t203 431.25
R4477 VDDH.t297 VDDH.t126 431.25
R4478 VDDH.t299 VDDH.t297 431.25
R4479 VDDH.t295 VDDH.t296 431.25
R4480 VDDH.t296 VDDH.t298 431.25
R4481 VDDH.t298 VDDH.t124 431.25
R4482 VDDH.t136 VDDH.t128 431.25
R4483 VDDH.t138 VDDH.t136 431.25
R4484 VDDH.t132 VDDH.t138 431.25
R4485 VDDH.t308 VDDH.t137 431.25
R4486 VDDH.t137 VDDH.t131 431.25
R4487 VDDH.t131 VDDH.t133 431.25
R4488 VDDH.t142 VDDH.t223 431.25
R4489 VDDH.t225 VDDH.t142 431.25
R4490 VDDH.t227 VDDH.t225 431.25
R4491 VDDH.t228 VDDH.t144 431.25
R4492 VDDH.t144 VDDH.t145 431.25
R4493 VDDH.t145 VDDH.t191 431.25
R4494 VDDH.t125 VDDH.t123 431.25
R4495 VDDH.t300 VDDH.t125 431.25
R4496 VDDH.t200 VDDH.t300 431.25
R4497 VDDH.t202 VDDH.t198 431.25
R4498 VDDH.t198 VDDH.t199 431.25
R4499 VDDH.t199 VDDH.t201 431.25
R4500 VDDH.t139 VDDH.t309 431.25
R4501 VDDH.t135 VDDH.t139 431.25
R4502 VDDH.t134 VDDH.t135 431.25
R4503 VDDH.t127 VDDH.t129 431.25
R4504 VDDH.t129 VDDH.t130 431.25
R4505 VDDH.t130 VDDH.t140 431.25
R4506 VDDH.t193 VDDH.t143 431.25
R4507 VDDH.t195 VDDH.t193 431.25
R4508 VDDH.t196 VDDH.t195 431.25
R4509 VDDH.t192 VDDH.t194 431.25
R4510 VDDH.t194 VDDH.t226 431.25
R4511 VDDH.t226 VDDH.t222 431.25
R4512 VDDH.t284 VDDH.t90 431.25
R4513 VDDH.t237 VDDH.t176 431.25
R4514 VDDH.t280 VDDH.t281 431.25
R4515 VDDH.t58 VDDH.t56 431.25
R4516 VDDH.t57 VDDH.t58 431.25
R4517 VDDH.t52 VDDH.t55 431.25
R4518 VDDH.t54 VDDH.t52 431.25
R4519 VDDH.t54 VDDH.t51 431.25
R4520 VDDH.t53 VDDH.t51 431.25
R4521 VDDH.t64 VDDH.t141 431.25
R4522 VDDH.t59 VDDH.t64 431.25
R4523 VDDH.t59 VDDH.t61 431.25
R4524 VDDH.t61 VDDH.t60 431.25
R4525 VDDH.t213 VDDH.t217 431.25
R4526 VDDH.t210 VDDH.t213 431.25
R4527 VDDH.t216 VDDH.t210 431.25
R4528 VDDH.t220 VDDH.t216 431.25
R4529 VDDH.t220 VDDH.t218 431.25
R4530 VDDH.t218 VDDH.t214 431.25
R4531 VDDH.t214 VDDH.t219 431.25
R4532 VDDH.t219 VDDH.t215 431.25
R4533 VDDH.t34 VDDH.t179 431.25
R4534 VDDH.t179 VDDH.t35 431.25
R4535 VDDH.t35 VDDH.t33 431.25
R4536 VDDH.t178 VDDH.t33 431.25
R4537 VDDH.t178 VDDH.t307 431.25
R4538 VDDH.t307 VDDH.t177 431.25
R4539 VDDH.t177 VDDH.t36 431.25
R4540 VDDH.t36 VDDH.t306 431.25
R4541 VDDH.n347 VDDH.n346 428.048
R4542 VDDH.n702 VDDH.n6 422.024
R4543 VDDH.n697 VDDH.n6 409.976
R4544 VDDH.n503 VDDH.n502 406.589
R4545 VDDH.n704 VDDH.n4 397.93
R4546 VDDH.t108 VDDH.n516 379.062
R4547 VDDH.t96 VDDH.n378 379.062
R4548 VDDH.t112 VDDH.n429 379.062
R4549 VDDH.t48 VDDH.n430 379.062
R4550 VDDH.t70 VDDH.n413 379.062
R4551 VDDH.t238 VDDH.n414 379.062
R4552 VDDH.t282 VDDH.n422 379.062
R4553 VDDH.n424 VDDH.t283 379.062
R4554 VDDH.t107 VDDH.n383 379.062
R4555 VDDH.t109 VDDH.n384 379.062
R4556 VDDH.t203 VDDH.n388 379.062
R4557 VDDH.t124 VDDH.n389 379.062
R4558 VDDH.t128 VDDH.n448 379.062
R4559 VDDH.t133 VDDH.n450 379.062
R4560 VDDH.t223 VDDH.n407 379.062
R4561 VDDH.t191 VDDH.n408 379.062
R4562 VDDH.t123 VDDH.n394 379.062
R4563 VDDH.t201 VDDH.n395 379.062
R4564 VDDH.t309 VDDH.n399 379.062
R4565 VDDH.t140 VDDH.n400 379.062
R4566 VDDH.t143 VDDH.n467 379.062
R4567 VDDH.t222 VDDH.n468 379.062
R4568 VDDH.t90 VDDH.n317 379.062
R4569 VDDH.t60 VDDH.n327 379.062
R4570 VDDH.t217 VDDH.n310 379.062
R4571 VDDH.t306 VDDH.n305 379.062
R4572 VDDH.t69 VDDH.t229 378.611
R4573 VDDH.t240 VDDH.t158 378.611
R4574 VDDH.t169 VDDH.t122 378.611
R4575 VDDH.t197 VDDH.t81 378.611
R4576 VDDH.t150 VDDH.t187 378.611
R4577 VDDH.t186 VDDH.t288 378.611
R4578 VDDH.t160 VDDH.t92 378.611
R4579 VDDH.t156 VDDH.t303 378.611
R4580 VDDH.n427 VDDH.n417 371.2
R4581 VDDH.n458 VDDH.n457 368.942
R4582 VDDH.n465 VDDH.n404 368.942
R4583 VDDH.n331 VDDH.n330 360.283
R4584 VDDH.n323 VDDH.n318 353.793
R4585 VDDH.n323 VDDH.n319 353.793
R4586 VDDH.n328 VDDH.n325 353.793
R4587 VDDH.n328 VDDH.n322 353.793
R4588 VDDH.n353 VDDH.n309 353.793
R4589 VDDH.n309 VDDH.n308 353.793
R4590 VDDH.n439 VDDH.n438 352.377
R4591 VDDH.n466 VDDH.n465 343.341
R4592 VDDH.n476 VDDH.n404 343.341
R4593 VDDH.n479 VDDH.n401 343.341
R4594 VDDH.n481 VDDH.n391 343.341
R4595 VDDH.n497 VDDH.n496 343.341
R4596 VDDH.n393 VDDH.n382 343.341
R4597 VDDH.n478 VDDH.n477 339.954
R4598 VDDH.n470 VDDH.n398 339.954
R4599 VDDH.n704 VDDH.n703 339.954
R4600 VDDH.n324 VDDH.t57 332.812
R4601 VDDH.t55 VDDH.n324 332.812
R4602 VDDH.n329 VDDH.t53 332.812
R4603 VDDH.t141 VDDH.n329 332.812
R4604 VDDH.t215 VDDH.n314 332.812
R4605 VDDH.n314 VDDH.t34 332.812
R4606 VDDH.n459 VDDH.n409 332.8
R4607 VDDH.n456 VDDH.n411 332.8
R4608 VDDH.n446 VDDH.n445 332.8
R4609 VDDH.n503 VDDH.n386 332.8
R4610 VDDH.n38 VDDH.t290 330.12
R4611 VDDH.n50 VDDH.t78 330.12
R4612 VDDH.n69 VDDH.t292 330.12
R4613 VDDH.n71 VDDH.t77 330.12
R4614 VDDH.n35 VDDH.t185 330.12
R4615 VDDH.n36 VDDH.t293 330.12
R4616 VDDH.n665 VDDH.t79 330.12
R4617 VDDH.n664 VDDH.t182 330.12
R4618 VDDH.n663 VDDH.t80 330.12
R4619 VDDH.n662 VDDH.t42 330.12
R4620 VDDH.n660 VDDH.t183 330.12
R4621 VDDH.n659 VDDH.t291 330.12
R4622 VDDH.n653 VDDH.n41 321.882
R4623 VDDH.n58 VDDH.n43 321.882
R4624 VDDH.n650 VDDH.n48 321.882
R4625 VDDH.n640 VDDH.n45 321.882
R4626 VDDH.n249 VDDH.n248 321.882
R4627 VDDH.n262 VDDH.n252 321.882
R4628 VDDH.n237 VDDH.n236 321.882
R4629 VDDH.n568 VDDH.n208 321.882
R4630 VDDH.n225 VDDH.n208 321.882
R4631 VDDH.n225 VDDH.n221 321.882
R4632 VDDH.n222 VDDH.n221 321.882
R4633 VDDH.n556 VDDH.n222 321.882
R4634 VDDH.n161 VDDH.n160 321.882
R4635 VDDH.n162 VDDH.n161 321.882
R4636 VDDH.n573 VDDH.n162 321.882
R4637 VDDH.n573 VDDH.n572 321.882
R4638 VDDH.n572 VDDH.n206 321.882
R4639 VDDH.n187 VDDH.n177 321.882
R4640 VDDH.n187 VDDH.n171 321.882
R4641 VDDH.n192 VDDH.n171 321.882
R4642 VDDH.n192 VDDH.n168 321.882
R4643 VDDH.n201 VDDH.n168 321.882
R4644 VDDH.n604 VDDH.n141 321.882
R4645 VDDH.n151 VDDH.n141 321.882
R4646 VDDH.n593 VDDH.n151 321.882
R4647 VDDH.n593 VDDH.n152 321.882
R4648 VDDH.n174 VDDH.n152 321.882
R4649 VDDH.n619 VDDH.n119 321.882
R4650 VDDH.n136 VDDH.n119 321.882
R4651 VDDH.n136 VDDH.n132 321.882
R4652 VDDH.n133 VDDH.n132 321.882
R4653 VDDH.n607 VDDH.n133 321.882
R4654 VDDH.n76 VDDH.n75 321.882
R4655 VDDH.n77 VDDH.n76 321.882
R4656 VDDH.n624 VDDH.n77 321.882
R4657 VDDH.n624 VDDH.n623 321.882
R4658 VDDH.n623 VDDH.n117 321.882
R4659 VDDH.n98 VDDH.n89 321.882
R4660 VDDH.n98 VDDH.n87 321.882
R4661 VDDH.n103 VDDH.n87 321.882
R4662 VDDH.n103 VDDH.n84 321.882
R4663 VDDH.n112 VDDH.n84 321.882
R4664 VDDH.n535 VDDH.n268 321.882
R4665 VDDH.n393 VDDH.n380 320
R4666 VDDH.n469 VDDH.n466 313.224
R4667 VDDH.n401 VDDH.n391 310.966
R4668 VDDH.n481 VDDH.n480 306.825
R4669 VDDH.n480 VDDH.n392 297.788
R4670 VDDH.n488 VDDH.n487 297.788
R4671 VDDH.n514 VDDH.n513 295.154
R4672 VDDH.n682 VDDH.n12 294.767
R4673 VDDH.n280 VDDH.n19 292.601
R4674 VDDH.n683 VDDH.n21 288.753
R4675 VDDH.n340 VDDH.n339 288
R4676 VDDH.n339 VDDH.n321 288
R4677 VDDH.n331 VDDH.n321 288
R4678 VDDH.n336 VDDH.n316 288
R4679 VDDH.n336 VDDH.n335 288
R4680 VDDH.n335 VDDH.n334 288
R4681 VDDH.n506 VDDH.n504 284.613
R4682 VDDH.n497 VDDH.n382 284.613
R4683 VDDH.n496 VDDH.n392 283.106
R4684 VDDH.n434 VDDH.t166 281.25
R4685 VDDH.n457 VDDH.n456 277.836
R4686 VDDH.n477 VDDH.n476 277.836
R4687 VDDH.n447 VDDH.n446 273.695
R4688 VDDH.n514 VDDH.n380 272.565
R4689 VDDH.n490 VDDH.n379 272.565
R4690 VDDH.n652 VDDH.n40 271.068
R4691 VDDH.n60 VDDH.n44 271.068
R4692 VDDH.n647 VDDH.n47 271.068
R4693 VDDH.n639 VDDH.n46 271.068
R4694 VDDH.n543 VDDH.n542 271.068
R4695 VDDH.n253 VDDH.n251 271.068
R4696 VDDH.n239 VDDH.n238 271.068
R4697 VDDH.n528 VDDH.n267 271.068
R4698 VDDH.n349 VDDH.n347 270.307
R4699 VDDH.n357 VDDH.n306 270.307
R4700 VDDH.n316 VDDH.n307 270.307
R4701 VDDH.n479 VDDH.n478 269.93
R4702 VDDH.n657 VDDH.t304 252.982
R4703 VDDH.n55 VDDH.t181 252.982
R4704 VDDH.n66 VDDH.t6 252.982
R4705 VDDH.n644 VDDH.t89 252.982
R4706 VDDH.n94 VDDH.t212 252.982
R4707 VDDH.n108 VDDH.t47 252.982
R4708 VDDH.n629 VDDH.t63 252.982
R4709 VDDH.n126 VDDH.t31 252.982
R4710 VDDH.n614 VDDH.t279 252.982
R4711 VDDH.n144 VDDH.t115 252.982
R4712 VDDH.n599 VDDH.t101 252.982
R4713 VDDH.n588 VDDH.t11 252.982
R4714 VDDH.n183 VDDH.t269 252.982
R4715 VDDH.n197 VDDH.t4 252.982
R4716 VDDH.n578 VDDH.t39 252.982
R4717 VDDH.n215 VDDH.t206 252.982
R4718 VDDH.n563 VDDH.t50 252.982
R4719 VDDH.n243 VDDH.t68 252.982
R4720 VDDH.n550 VDDH.t1 252.982
R4721 VDDH.n257 VDDH.t273 252.982
R4722 VDDH.n270 VDDH.t302 252.982
R4723 VDDH.n531 VDDH.t66 252.982
R4724 VDDH.n692 VDDH.n19 248.9
R4725 VDDH.n459 VDDH.n458 240.941
R4726 VDDH.n428 VDDH.n427 236.8
R4727 VDDH.n439 VDDH.n437 236.8
R4728 VDDH.n343 VDDH.t281 235.939
R4729 VDDH.n330 VDDH.n306 232.66
R4730 VDDH.n28 VDDH.t149 227.737
R4731 VDDH.n672 VDDH.t184 226.81
R4732 VDDH.n513 VDDH 225.882
R4733 VDDH.n518 VDDH.t119 215.625
R4734 VDDH.n518 VDDH.t93 215.625
R4735 VDDH.n442 VDDH.t98 215.625
R4736 VDDH.n442 VDDH.t71 215.625
R4737 VDDH.n423 VDDH.t104 215.625
R4738 VDDH.t91 VDDH.n423 215.625
R4739 VDDH.n509 VDDH.t121 215.625
R4740 VDDH.n509 VDDH.t110 215.625
R4741 VDDH.n500 VDDH.t299 215.625
R4742 VDDH.n500 VDDH.t295 215.625
R4743 VDDH.n453 VDDH.t132 215.625
R4744 VDDH.n453 VDDH.t308 215.625
R4745 VDDH.n462 VDDH.t227 215.625
R4746 VDDH.n462 VDDH.t228 215.625
R4747 VDDH.n493 VDDH.t200 215.625
R4748 VDDH.n493 VDDH.t202 215.625
R4749 VDDH.n484 VDDH.t134 215.625
R4750 VDDH.n484 VDDH.t127 215.625
R4751 VDDH.n473 VDDH.t196 215.625
R4752 VDDH.n473 VDDH.t192 215.625
R4753 VDDH.n347 VDDH.n315 207.812
R4754 VDDH.n460 VDDH.n459 202.918
R4755 VDDH.n475 VDDH.n466 202.918
R4756 VDDH.n301 VDDH.n4 200.282
R4757 VDDH.n283 VDDH.n282 200.282
R4758 VDDH.n266 VDDH.n265 200.111
R4759 VDDH.n247 VDDH.n246 200.111
R4760 VDDH.n259 VDDH.n254 200.111
R4761 VDDH.n552 VDDH.n232 200.111
R4762 VDDH.n561 VDDH.n218 200.111
R4763 VDDH.n577 VDDH.n165 200.111
R4764 VDDH.n181 VDDH.n180 200.111
R4765 VDDH.n597 VDDH.n147 200.111
R4766 VDDH.n612 VDDH.n129 200.111
R4767 VDDH.n628 VDDH.n80 200.111
R4768 VDDH.n92 VDDH.n91 200.111
R4769 VDDH.n344 VDDH.t277 193.75
R4770 VDDH.n96 VDDH.n89 191.167
R4771 VDDH.t229 VDDH.n554 189.305
R4772 VDDH.n554 VDDH.t158 189.305
R4773 VDDH.n264 VDDH.t169 189.305
R4774 VDDH.t81 VDDH.n264 189.305
R4775 VDDH.n540 VDDH.t150 189.305
R4776 VDDH.n540 VDDH.t288 189.305
R4777 VDDH.n537 VDDH.t160 189.305
R4778 VDDH.n537 VDDH.t156 189.305
R4779 VDDH.n544 VDDH.n249 185
R4780 VDDH.n545 VDDH.n248 185
R4781 VDDH.n541 VDDH.n248 185
R4782 VDDH.n260 VDDH.n252 185
R4783 VDDH.n262 VDDH.n261 185
R4784 VDDH.n263 VDDH.n262 185
R4785 VDDH.n237 VDDH.n234 185
R4786 VDDH.n236 VDDH.n235 185
R4787 VDDH.n236 VDDH.n230 185
R4788 VDDH.n112 VDDH.n111 185
R4789 VDDH.n113 VDDH.n112 185
R4790 VDDH.n85 VDDH.n84 185
R4791 VDDH.n84 VDDH.n83 185
R4792 VDDH.n104 VDDH.n103 185
R4793 VDDH.n103 VDDH.n102 185
R4794 VDDH.n87 VDDH.n86 185
R4795 VDDH.n100 VDDH.n87 185
R4796 VDDH.n98 VDDH.n97 185
R4797 VDDH.n99 VDDH.n98 185
R4798 VDDH.n89 VDDH.n88 185
R4799 VDDH.n121 VDDH.n117 185
R4800 VDDH.n621 VDDH.n117 185
R4801 VDDH.n623 VDDH.n118 185
R4802 VDDH.n623 VDDH.n622 185
R4803 VDDH.n624 VDDH.n78 185
R4804 VDDH.n625 VDDH.n624 185
R4805 VDDH.n632 VDDH.n77 185
R4806 VDDH.n116 VDDH.n77 185
R4807 VDDH.n633 VDDH.n76 185
R4808 VDDH.n115 VDDH.n76 185
R4809 VDDH.n634 VDDH.n75 185
R4810 VDDH.n114 VDDH.n75 185
R4811 VDDH.n608 VDDH.n607 185
R4812 VDDH.n607 VDDH.n606 185
R4813 VDDH.n609 VDDH.n133 185
R4814 VDDH.n140 VDDH.n133 185
R4815 VDDH.n610 VDDH.n132 185
R4816 VDDH.n139 VDDH.n132 185
R4817 VDDH.n136 VDDH.n131 185
R4818 VDDH.n137 VDDH.n136 185
R4819 VDDH.n120 VDDH.n119 185
R4820 VDDH.n135 VDDH.n119 185
R4821 VDDH.n619 VDDH.n618 185
R4822 VDDH.n620 VDDH.n619 185
R4823 VDDH.n174 VDDH.n173 185
R4824 VDDH.n175 VDDH.n174 185
R4825 VDDH.n154 VDDH.n152 185
R4826 VDDH.n172 VDDH.n152 185
R4827 VDDH.n593 VDDH.n592 185
R4828 VDDH.n594 VDDH.n593 185
R4829 VDDH.n153 VDDH.n151 185
R4830 VDDH.n151 VDDH.n150 185
R4831 VDDH.n142 VDDH.n141 185
R4832 VDDH.n149 VDDH.n141 185
R4833 VDDH.n604 VDDH.n603 185
R4834 VDDH.n605 VDDH.n604 185
R4835 VDDH.n201 VDDH.n200 185
R4836 VDDH.n202 VDDH.n201 185
R4837 VDDH.n169 VDDH.n168 185
R4838 VDDH.n168 VDDH.n167 185
R4839 VDDH.n193 VDDH.n192 185
R4840 VDDH.n192 VDDH.n191 185
R4841 VDDH.n171 VDDH.n170 185
R4842 VDDH.n189 VDDH.n171 185
R4843 VDDH.n187 VDDH.n186 185
R4844 VDDH.n188 VDDH.n187 185
R4845 VDDH.n178 VDDH.n177 185
R4846 VDDH.n177 VDDH.n176 185
R4847 VDDH.n210 VDDH.n206 185
R4848 VDDH.n570 VDDH.n206 185
R4849 VDDH.n572 VDDH.n207 185
R4850 VDDH.n572 VDDH.n571 185
R4851 VDDH.n573 VDDH.n163 185
R4852 VDDH.n574 VDDH.n573 185
R4853 VDDH.n581 VDDH.n162 185
R4854 VDDH.n205 VDDH.n162 185
R4855 VDDH.n582 VDDH.n161 185
R4856 VDDH.n204 VDDH.n161 185
R4857 VDDH.n583 VDDH.n160 185
R4858 VDDH.n203 VDDH.n160 185
R4859 VDDH.n557 VDDH.n556 185
R4860 VDDH.n556 VDDH.n555 185
R4861 VDDH.n558 VDDH.n222 185
R4862 VDDH.n229 VDDH.n222 185
R4863 VDDH.n559 VDDH.n221 185
R4864 VDDH.n228 VDDH.n221 185
R4865 VDDH.n225 VDDH.n220 185
R4866 VDDH.n226 VDDH.n225 185
R4867 VDDH.n209 VDDH.n208 185
R4868 VDDH.n224 VDDH.n208 185
R4869 VDDH.n568 VDDH.n567 185
R4870 VDDH.n569 VDDH.n568 185
R4871 VDDH.n535 VDDH.n534 185
R4872 VDDH.n536 VDDH.n535 185
R4873 VDDH.n529 VDDH.n268 185
R4874 VDDH.n641 VDDH.n640 185
R4875 VDDH.n72 VDDH.n45 185
R4876 VDDH.n651 VDDH.n45 185
R4877 VDDH.n648 VDDH.n48 185
R4878 VDDH.n650 VDDH.n649 185
R4879 VDDH.n651 VDDH.n650 185
R4880 VDDH.n59 VDDH.n58 185
R4881 VDDH.n51 VDDH.n43 185
R4882 VDDH.n651 VDDH.n43 185
R4883 VDDH.n654 VDDH.n653 185
R4884 VDDH.n41 VDDH.n39 185
R4885 VDDH.n651 VDDH.n41 185
R4886 VDDH.t44 VDDH.t148 179.685
R4887 VDDH.t44 VDDH.n671 175.309
R4888 VDDH.n482 VDDH.n479 173.929
R4889 VDDH.t40 VDDH.t7 168.685
R4890 VDDH.t76 VDDH.t8 168.685
R4891 VDDH.n456 VDDH.n455 166.024
R4892 VDDH.n476 VDDH.n475 166.024
R4893 VDDH.n440 VDDH.n439 163.766
R4894 VDDH.n496 VDDH.n495 160.754
R4895 VDDH.n42 VDDH.t76 158.225
R4896 VDDH.n683 VDDH.n682 152.471
R4897 VDDH.n434 VDDH.t165 150
R4898 VDDH.n513 VDDH.n377 148.707
R4899 VDDH.n651 VDDH.t5 144.494
R4900 VDDH.n9 VDDH.t245 139.454
R4901 VDDH.n2 VDDH.t258 139.454
R4902 VDDH.n303 VDDH.t248 139.454
R4903 VDDH.n290 VDDH.t255 139.454
R4904 VDDH.n288 VDDH.t264 139.454
R4905 VDDH.n24 VDDH.t241 139.454
R4906 VDDH.n26 VDDH.t252 139.454
R4907 VDDH.n369 VDDH.t261 139.454
R4908 VDDH.n482 VDDH.n481 137.036
R4909 VDDH.n361 VDDH.t251 135.362
R4910 VDDH.n8 VDDH.t247 135.312
R4911 VDDH.n8 VDDH.t246 135.312
R4912 VDDH.n1 VDDH.t260 135.312
R4913 VDDH.n1 VDDH.t259 135.312
R4914 VDDH.n287 VDDH.t265 135.312
R4915 VDDH.n287 VDDH.t266 135.312
R4916 VDDH.n289 VDDH.t257 135.312
R4917 VDDH.n23 VDDH.t244 135.312
R4918 VDDH.n23 VDDH.t243 135.312
R4919 VDDH.n25 VDDH.t253 135.312
R4920 VDDH.n25 VDDH.t254 135.312
R4921 VDDH.n370 VDDH.t262 135.312
R4922 VDDH.n302 VDDH.t250 135.312
R4923 VDDH.n286 VDDH.t256 134.712
R4924 VDDH.n286 VDDH.t20 134.712
R4925 VDDH.n292 VDDH.t17 134.712
R4926 VDDH.n292 VDDH.t26 134.712
R4927 VDDH.n284 VDDH.t13 134.712
R4928 VDDH.n284 VDDH.t22 134.712
R4929 VDDH.n367 VDDH.t23 134.712
R4930 VDDH.n367 VDDH.t263 134.712
R4931 VDDH.n273 VDDH.t25 134.712
R4932 VDDH.n273 VDDH.t18 134.712
R4933 VDDH.n274 VDDH.t15 134.712
R4934 VDDH.n274 VDDH.t19 134.712
R4935 VDDH.n670 VDDH.n669 129.44
R4936 VDDH.n334 VDDH.n306 127.624
R4937 VDDH.n671 VDDH.t32 125.675
R4938 VDDH.n495 VDDH.n393 123.859
R4939 VDDH VDDH.n512 117.46
R4940 VDDH.t21 VDDH.t242 113.218
R4941 VDDH.t24 VDDH.t12 113.218
R4942 VDDH.t14 VDDH.t16 113.218
R4943 VDDH.t249 VDDH.t14 113.218
R4944 VDDH.n681 VDDH.n6 106.541
R4945 VDDH.n682 VDDH.n681 106.165
R4946 VDDH.n279 VDDH.t21 105.088
R4947 VDDH.t41 VDDH.n668 102.35
R4948 VDDH.n696 VDDH.n12 101.272
R4949 VDDH.t28 VDDH.t74 100.906
R4950 VDDH.t180 VDDH.t41 100.906
R4951 VDDH.t16 VDDH.n298 99.0655
R4952 VDDH.n678 VDDH.n12 96.9471
R4953 VDDH.t32 VDDH.t204 95.9301
R4954 VDDH.t294 VDDH.t184 95.9301
R4955 VDDH.n113 VDDH.n83 92.2149
R4956 VDDH.n622 VDDH.n621 92.2149
R4957 VDDH.n606 VDDH.n140 92.2149
R4958 VDDH.n175 VDDH.n172 92.2149
R4959 VDDH.n202 VDDH.n167 92.2149
R4960 VDDH.n571 VDDH.n570 92.2149
R4961 VDDH.n555 VDDH.n229 92.2149
R4962 VDDH.n88 VDDH.t211 89.3332
R4963 VDDH.t62 VDDH.n114 89.3332
R4964 VDDH.n620 VDDH.t278 89.3332
R4965 VDDH.n605 VDDH.t100 89.3332
R4966 VDDH.n176 VDDH.t268 89.3332
R4967 VDDH.t38 VDDH.n203 89.3332
R4968 VDDH.n569 VDDH.t49 89.3332
R4969 VDDH.n542 VDDH.n249 86.068
R4970 VDDH.n252 VDDH.n251 86.068
R4971 VDDH.n238 VDDH.n237 86.068
R4972 VDDH.n268 VDDH.n267 86.068
R4973 VDDH.n640 VDDH.n46 86.068
R4974 VDDH.n48 VDDH.n47 86.068
R4975 VDDH.n58 VDDH.n44 86.068
R4976 VDDH.n653 VDDH.n652 86.068
R4977 VDDH.n88 VDDH.t45 84.5303
R4978 VDDH.n114 VDDH.t29 84.5303
R4979 VDDH.t221 VDDH.n620 84.5303
R4980 VDDH.t9 VDDH.n605 84.5303
R4981 VDDH.n176 VDDH.t2 84.5303
R4982 VDDH.n203 VDDH.t207 84.5303
R4983 VDDH.t175 VDDH.n569 84.5303
R4984 VDDH.n32 VDDH.t7 84.3432
R4985 VDDH.t8 VDDH.n32 84.3432
R4986 VDDH.t164 VDDH.n113 82.6092
R4987 VDDH.n621 VDDH.t274 82.6092
R4988 VDDH.n606 VDDH.t75 82.6092
R4989 VDDH.t27 VDDH.n175 82.6092
R4990 VDDH.t305 VDDH.n202 82.6092
R4991 VDDH.n570 VDDH.t310 82.6092
R4992 VDDH.n555 VDDH.t209 82.6092
R4993 VDDH.n694 VDDH.t155 82.5045
R4994 VDDH.t154 VDDH.n693 82.5045
R4995 VDDH.t204 VDDH.n670 81.8009
R4996 VDDH.n348 VDDH 77.9299
R4997 VDDH.t155 VDDH.t154 77.6867
R4998 VDDH.t242 VDDH.n17 72.869
R4999 VDDH.n299 VDDH.t249 72.869
R5000 VDDH.n427 VDDH.n426 72.6593
R5001 VDDH.n437 VDDH.n416 72.2828
R5002 VDDH.n431 VDDH.n428 72.2828
R5003 VDDH.n438 VDDH.n386 72.2828
R5004 VDDH.n426 VDDH.n425 72.2828
R5005 VDDH.n425 VDDH.n411 72.2828
R5006 VDDH.n421 VDDH.n409 72.2828
R5007 VDDH.n415 VDDH.n412 72.2828
R5008 VDDH.n445 VDDH.n412 72.2828
R5009 VDDH.n512 VDDH.n381 72.2828
R5010 VDDH.n504 VDDH.n385 72.2828
R5011 VDDH.n497 VDDH.n385 72.2828
R5012 VDDH.n390 VDDH.n387 72.2828
R5013 VDDH.n391 VDDH.n390 72.2828
R5014 VDDH.n449 VDDH.n447 72.2828
R5015 VDDH.n449 VDDH.n401 72.2828
R5016 VDDH.n457 VDDH.n410 72.2828
R5017 VDDH.n410 VDDH.n404 72.2828
R5018 VDDH.n458 VDDH.n405 72.2828
R5019 VDDH.n465 VDDH.n405 72.2828
R5020 VDDH.n506 VDDH.n505 72.2828
R5021 VDDH.n505 VDDH.n382 72.2828
R5022 VDDH.n489 VDDH.n380 72.2828
R5023 VDDH.n490 VDDH.n489 72.2828
R5024 VDDH.n396 VDDH.n392 72.2828
R5025 VDDH.n488 VDDH.n396 72.2828
R5026 VDDH.n480 VDDH.n397 72.2828
R5027 VDDH.n487 VDDH.n397 72.2828
R5028 VDDH.n478 VDDH.n402 72.2828
R5029 VDDH.n402 VDDH.n398 72.2828
R5030 VDDH.n477 VDDH.n403 72.2828
R5031 VDDH.n470 VDDH.n403 72.2828
R5032 VDDH.n515 VDDH.n514 72.2828
R5033 VDDH.n515 VDDH.n379 72.2828
R5034 VDDH.n335 VDDH.n326 72.2828
R5035 VDDH.n326 VDDH.n321 72.2828
R5036 VDDH.n320 VDDH.n316 72.2828
R5037 VDDH.n340 VDDH.n320 72.2828
R5038 VDDH.n349 VDDH.n348 72.2828
R5039 VDDH.n312 VDDH.n311 72.2828
R5040 VDDH.n311 VDDH.n307 72.2828
R5041 VDDH.n358 VDDH.n357 72.2828
R5042 VDDH.n651 VDDH.n42 66.0363
R5043 VDDH.n299 VDDH.n5 63.1385
R5044 VDDH.n100 VDDH.t83 59.5556
R5045 VDDH.n116 VDDH.t270 59.5556
R5046 VDDH.n137 VDDH.t233 59.5556
R5047 VDDH.n150 VDDH.t87 59.5556
R5048 VDDH.n189 VDDH.t173 59.5556
R5049 VDDH.n205 VDDH.t286 59.5556
R5050 VDDH.n226 VDDH.t231 59.5556
R5051 VDDH.n283 VDDH.n21 57.977
R5052 VDDH.n102 VDDH.t171 57.6345
R5053 VDDH.n625 VDDH.t152 57.6345
R5054 VDDH.t162 VDDH.n139 57.6345
R5055 VDDH.n594 VDDH.t85 57.6345
R5056 VDDH.n191 VDDH.t167 57.6345
R5057 VDDH.n574 VDDH.t146 57.6345
R5058 VDDH.t235 VDDH.n228 57.6345
R5059 VDDH.n694 VDDH.n15 55.8602
R5060 VDDH.n691 VDDH.n21 54.2123
R5061 VDDH.n371 VDDH.n370 52.8457
R5062 VDDH.n11 VDDH.n10 50.7802
R5063 VDDH.n698 VDDH.n11 50.7802
R5064 VDDH.n32 VDDH.t28 50.4534
R5065 VDDH.n542 VDDH.n541 49.4675
R5066 VDDH.n263 VDDH.n251 49.4675
R5067 VDDH.n238 VDDH.n230 49.4675
R5068 VDDH.n536 VDDH.n267 49.4675
R5069 VDDH.n651 VDDH.n46 49.4675
R5070 VDDH.n651 VDDH.n47 49.4675
R5071 VDDH.n651 VDDH.n44 49.4675
R5072 VDDH.n652 VDDH.n651 49.4675
R5073 VDDH.n102 VDDH.n101 47.0682
R5074 VDDH.n626 VDDH.n625 47.0682
R5075 VDDH.n139 VDDH.n138 47.0682
R5076 VDDH.n595 VDDH.n594 47.0682
R5077 VDDH.n191 VDDH.n190 47.0682
R5078 VDDH.n575 VDDH.n574 47.0682
R5079 VDDH.n228 VDDH.n227 47.0682
R5080 VDDH.n693 VDDH.n17 46.3713
R5081 VDDH.n430 VDDH.n416 46.2505
R5082 VDDH.n431 VDDH.n429 46.2505
R5083 VDDH.n438 VDDH.n414 46.2505
R5084 VDDH.n425 VDDH.n424 46.2505
R5085 VDDH.n422 VDDH.n421 46.2505
R5086 VDDH.n413 VDDH.n412 46.2505
R5087 VDDH.n384 VDDH.n381 46.2505
R5088 VDDH.n389 VDDH.n385 46.2505
R5089 VDDH.n390 VDDH.n388 46.2505
R5090 VDDH.n450 VDDH.n449 46.2505
R5091 VDDH.n448 VDDH.n410 46.2505
R5092 VDDH.n408 VDDH.n405 46.2505
R5093 VDDH.n407 VDDH.n406 46.2505
R5094 VDDH.n505 VDDH.n383 46.2505
R5095 VDDH.n489 VDDH.n395 46.2505
R5096 VDDH.n396 VDDH.n394 46.2505
R5097 VDDH.n400 VDDH.n397 46.2505
R5098 VDDH.n402 VDDH.n399 46.2505
R5099 VDDH.n468 VDDH.n403 46.2505
R5100 VDDH.n469 VDDH.n467 46.2505
R5101 VDDH.n516 VDDH.n515 46.2505
R5102 VDDH.n521 VDDH.n378 46.2505
R5103 VDDH.n323 VDDH.n320 46.2505
R5104 VDDH.n324 VDDH.n323 46.2505
R5105 VDDH.n328 VDDH.n326 46.2505
R5106 VDDH.n329 VDDH.n328 46.2505
R5107 VDDH.n330 VDDH.n327 46.2505
R5108 VDDH.n317 VDDH.n315 46.2505
R5109 VDDH.n348 VDDH.n310 46.2505
R5110 VDDH.n311 VDDH.n309 46.2505
R5111 VDDH.n314 VDDH.n309 46.2505
R5112 VDDH.n358 VDDH.n305 46.2505
R5113 VDDH.n101 VDDH.n100 45.1471
R5114 VDDH.n626 VDDH.n116 45.1471
R5115 VDDH.n138 VDDH.n137 45.1471
R5116 VDDH.n595 VDDH.n150 45.1471
R5117 VDDH.n190 VDDH.n189 45.1471
R5118 VDDH.n575 VDDH.n205 45.1471
R5119 VDDH.n227 VDDH.n226 45.1471
R5120 VDDH.n446 VDDH.n387 37.2711
R5121 VDDH.n504 VDDH.n503 37.2711
R5122 VDDH.n654 VDDH.n39 36.1417
R5123 VDDH.n654 VDDH.n40 36.1417
R5124 VDDH.n59 VDDH.n51 36.1417
R5125 VDDH.n60 VDDH.n59 36.1417
R5126 VDDH.n649 VDDH.n648 36.1417
R5127 VDDH.n648 VDDH.n647 36.1417
R5128 VDDH.n545 VDDH.n544 36.1417
R5129 VDDH.n544 VDDH.n543 36.1417
R5130 VDDH.n261 VDDH.n260 36.1417
R5131 VDDH.n260 VDDH.n253 36.1417
R5132 VDDH.n235 VDDH.n234 36.1417
R5133 VDDH.n239 VDDH.n234 36.1417
R5134 VDDH.n567 VDDH.n209 36.1417
R5135 VDDH.n220 VDDH.n209 36.1417
R5136 VDDH.n559 VDDH.n220 36.1417
R5137 VDDH.n559 VDDH.n558 36.1417
R5138 VDDH.n558 VDDH.n557 36.1417
R5139 VDDH.n583 VDDH.n582 36.1417
R5140 VDDH.n582 VDDH.n581 36.1417
R5141 VDDH.n581 VDDH.n163 36.1417
R5142 VDDH.n207 VDDH.n163 36.1417
R5143 VDDH.n210 VDDH.n207 36.1417
R5144 VDDH.n186 VDDH.n178 36.1417
R5145 VDDH.n186 VDDH.n170 36.1417
R5146 VDDH.n193 VDDH.n170 36.1417
R5147 VDDH.n193 VDDH.n169 36.1417
R5148 VDDH.n200 VDDH.n169 36.1417
R5149 VDDH.n603 VDDH.n142 36.1417
R5150 VDDH.n153 VDDH.n142 36.1417
R5151 VDDH.n592 VDDH.n153 36.1417
R5152 VDDH.n592 VDDH.n154 36.1417
R5153 VDDH.n173 VDDH.n154 36.1417
R5154 VDDH.n618 VDDH.n120 36.1417
R5155 VDDH.n131 VDDH.n120 36.1417
R5156 VDDH.n610 VDDH.n131 36.1417
R5157 VDDH.n610 VDDH.n609 36.1417
R5158 VDDH.n609 VDDH.n608 36.1417
R5159 VDDH.n634 VDDH.n633 36.1417
R5160 VDDH.n633 VDDH.n632 36.1417
R5161 VDDH.n632 VDDH.n78 36.1417
R5162 VDDH.n118 VDDH.n78 36.1417
R5163 VDDH.n121 VDDH.n118 36.1417
R5164 VDDH.n97 VDDH.n86 36.1417
R5165 VDDH.n104 VDDH.n86 36.1417
R5166 VDDH.n104 VDDH.n85 36.1417
R5167 VDDH.n111 VDDH.n85 36.1417
R5168 VDDH.n529 VDDH.n528 36.1417
R5169 VDDH.n534 VDDH.n529 36.1417
R5170 VDDH.n641 VDDH.n72 36.1417
R5171 VDDH.n641 VDDH.n639 36.1417
R5172 VDDH.n669 VDDH.n32 35.5918
R5173 VDDH.t83 VDDH.n99 32.6598
R5174 VDDH.t270 VDDH.n115 32.6598
R5175 VDDH.t233 VDDH.n135 32.6598
R5176 VDDH.t87 VDDH.n149 32.6598
R5177 VDDH.t173 VDDH.n188 32.6598
R5178 VDDH.t286 VDDH.n204 32.6598
R5179 VDDH.t231 VDDH.n224 32.6598
R5180 VDDH.t171 VDDH.t46 31.6992
R5181 VDDH.t30 VDDH.t152 31.6992
R5182 VDDH.t114 VDDH.t162 31.6992
R5183 VDDH.t10 VDDH.t85 31.6992
R5184 VDDH.t167 VDDH.t3 31.6992
R5185 VDDH.t205 VDDH.t146 31.6992
R5186 VDDH.t67 VDDH.t235 31.6992
R5187 VDDH.n265 VDDH.t161 27.6955
R5188 VDDH.n265 VDDH.t157 27.6955
R5189 VDDH.n246 VDDH.t151 27.6955
R5190 VDDH.n246 VDDH.t289 27.6955
R5191 VDDH.n254 VDDH.t170 27.6955
R5192 VDDH.n254 VDDH.t82 27.6955
R5193 VDDH.n232 VDDH.t230 27.6955
R5194 VDDH.n232 VDDH.t159 27.6955
R5195 VDDH.n218 VDDH.t232 27.6955
R5196 VDDH.n218 VDDH.t236 27.6955
R5197 VDDH.n165 VDDH.t287 27.6955
R5198 VDDH.n165 VDDH.t147 27.6955
R5199 VDDH.n180 VDDH.t174 27.6955
R5200 VDDH.n180 VDDH.t168 27.6955
R5201 VDDH.n147 VDDH.t88 27.6955
R5202 VDDH.n147 VDDH.t86 27.6955
R5203 VDDH.n129 VDDH.t234 27.6955
R5204 VDDH.n129 VDDH.t163 27.6955
R5205 VDDH.n80 VDDH.t271 27.6955
R5206 VDDH.n80 VDDH.t153 27.6955
R5207 VDDH.n91 VDDH.t84 27.6955
R5208 VDDH.n91 VDDH.t172 27.6955
R5209 VDDH.n696 VDDH.n695 23.1255
R5210 VDDH.n695 VDDH.n694 23.1255
R5211 VDDH.n681 VDDH.n16 23.1255
R5212 VDDH.n693 VDDH.n16 23.1255
R5213 VDDH.n359 VDDH.n358 20.252
R5214 VDDH.n668 VDDH.n667 19.4051
R5215 VDDH.n92 VDDH.n81 16.2626
R5216 VDDH.n628 VDDH.n627 16.2626
R5217 VDDH.n612 VDDH.n82 16.2626
R5218 VDDH.n597 VDDH.n596 16.2626
R5219 VDDH.n181 VDDH.n148 16.2626
R5220 VDDH.n577 VDDH.n576 16.2626
R5221 VDDH.n561 VDDH.n166 16.2626
R5222 VDDH.n553 VDDH.n552 16.2626
R5223 VDDH.n259 VDDH.n231 16.2626
R5224 VDDH.n539 VDDH.n247 16.2626
R5225 VDDH.n538 VDDH.n266 16.2626
R5226 VDDH.n101 VDDH.n81 15.4172
R5227 VDDH.n627 VDDH.n626 15.4172
R5228 VDDH.n138 VDDH.n82 15.4172
R5229 VDDH.n596 VDDH.n595 15.4172
R5230 VDDH.n190 VDDH.n148 15.4172
R5231 VDDH.n576 VDDH.n575 15.4172
R5232 VDDH.n227 VDDH.n166 15.4172
R5233 VDDH.n554 VDDH.n553 15.4172
R5234 VDDH.n264 VDDH.n231 15.4172
R5235 VDDH.n540 VDDH.n539 15.4172
R5236 VDDH.n538 VDDH.n537 15.4172
R5237 VDDH.n669 VDDH.t180 14.8631
R5238 VDDH.n522 VDDH.n521 14.4353
R5239 VDDH.n298 VDDH.t24 14.1526
R5240 VDDH.n670 VDDH.t294 14.1297
R5241 VDDH.n301 VDDH.n300 11.563
R5242 VDDH.n300 VDDH.n299 11.563
R5243 VDDH.n282 VDDH.n281 11.563
R5244 VDDH.n281 VDDH.n17 11.563
R5245 VDDH.n676 VDDH.n673 11.4005
R5246 VDDH.n541 VDDH.n540 11.31
R5247 VDDH.n264 VDDH.n263 11.31
R5248 VDDH.n554 VDDH.n230 11.31
R5249 VDDH.n537 VDDH.n536 11.31
R5250 VDDH.n680 VDDH.n678 11.2946
R5251 VDDH.n296 VDDH.n295 11.2946
R5252 VDDH.n677 VDDH.n15 10.9826
R5253 VDDH.n523 VDDH.t208 10.5739
R5254 VDDH.n63 VDDH.n62 9.73734
R5255 VDDH.n62 VDDH.n42 9.73734
R5256 VDDH.n34 VDDH.n33 9.73734
R5257 VDDH.n668 VDDH.n33 9.66826
R5258 VDDH.n531 VDDH.n530 9.3005
R5259 VDDH.n532 VDDH.n531 9.3005
R5260 VDDH.n534 VDDH.n533 9.3005
R5261 VDDH.n529 VDDH.n266 9.3005
R5262 VDDH.n528 VDDH.n527 9.3005
R5263 VDDH.n270 VDDH.n269 9.3005
R5264 VDDH.n271 VDDH.n270 9.3005
R5265 VDDH.n543 VDDH.n250 9.3005
R5266 VDDH.n544 VDDH.n247 9.3005
R5267 VDDH.n546 VDDH.n545 9.3005
R5268 VDDH.n258 VDDH.n257 9.3005
R5269 VDDH.n257 VDDH.n256 9.3005
R5270 VDDH.n255 VDDH.n253 9.3005
R5271 VDDH.n260 VDDH.n259 9.3005
R5272 VDDH.n261 VDDH.n241 9.3005
R5273 VDDH.n551 VDDH.n550 9.3005
R5274 VDDH.n550 VDDH.n549 9.3005
R5275 VDDH.n240 VDDH.n239 9.3005
R5276 VDDH.n552 VDDH.n234 9.3005
R5277 VDDH.n235 VDDH.n233 9.3005
R5278 VDDH.n243 VDDH.n242 9.3005
R5279 VDDH.n244 VDDH.n243 9.3005
R5280 VDDH.n564 VDDH.n563 9.3005
R5281 VDDH.n563 VDDH.n562 9.3005
R5282 VDDH.n557 VDDH.n223 9.3005
R5283 VDDH.n558 VDDH.n219 9.3005
R5284 VDDH.n560 VDDH.n559 9.3005
R5285 VDDH.n220 VDDH.n217 9.3005
R5286 VDDH.n565 VDDH.n209 9.3005
R5287 VDDH.n567 VDDH.n566 9.3005
R5288 VDDH.n215 VDDH.n214 9.3005
R5289 VDDH.n216 VDDH.n215 9.3005
R5290 VDDH.n578 VDDH.n164 9.3005
R5291 VDDH.n579 VDDH.n578 9.3005
R5292 VDDH.n211 VDDH.n210 9.3005
R5293 VDDH.n213 VDDH.n207 9.3005
R5294 VDDH.n212 VDDH.n163 9.3005
R5295 VDDH.n581 VDDH.n580 9.3005
R5296 VDDH.n582 VDDH.n159 9.3005
R5297 VDDH.n584 VDDH.n583 9.3005
R5298 VDDH.n197 VDDH.n196 9.3005
R5299 VDDH.n198 VDDH.n197 9.3005
R5300 VDDH.n184 VDDH.n183 9.3005
R5301 VDDH.n183 VDDH.n182 9.3005
R5302 VDDH.n200 VDDH.n199 9.3005
R5303 VDDH.n195 VDDH.n169 9.3005
R5304 VDDH.n194 VDDH.n193 9.3005
R5305 VDDH.n179 VDDH.n170 9.3005
R5306 VDDH.n186 VDDH.n185 9.3005
R5307 VDDH.n178 VDDH.n156 9.3005
R5308 VDDH.n589 VDDH.n588 9.3005
R5309 VDDH.n588 VDDH.n587 9.3005
R5310 VDDH.n600 VDDH.n599 9.3005
R5311 VDDH.n599 VDDH.n598 9.3005
R5312 VDDH.n173 VDDH.n155 9.3005
R5313 VDDH.n590 VDDH.n154 9.3005
R5314 VDDH.n592 VDDH.n591 9.3005
R5315 VDDH.n153 VDDH.n146 9.3005
R5316 VDDH.n601 VDDH.n142 9.3005
R5317 VDDH.n603 VDDH.n602 9.3005
R5318 VDDH.n144 VDDH.n143 9.3005
R5319 VDDH.n145 VDDH.n144 9.3005
R5320 VDDH.n615 VDDH.n614 9.3005
R5321 VDDH.n614 VDDH.n613 9.3005
R5322 VDDH.n608 VDDH.n134 9.3005
R5323 VDDH.n609 VDDH.n130 9.3005
R5324 VDDH.n611 VDDH.n610 9.3005
R5325 VDDH.n131 VDDH.n128 9.3005
R5326 VDDH.n616 VDDH.n120 9.3005
R5327 VDDH.n618 VDDH.n617 9.3005
R5328 VDDH.n126 VDDH.n125 9.3005
R5329 VDDH.n127 VDDH.n126 9.3005
R5330 VDDH.n629 VDDH.n79 9.3005
R5331 VDDH.n630 VDDH.n629 9.3005
R5332 VDDH.n122 VDDH.n121 9.3005
R5333 VDDH.n124 VDDH.n118 9.3005
R5334 VDDH.n123 VDDH.n78 9.3005
R5335 VDDH.n632 VDDH.n631 9.3005
R5336 VDDH.n633 VDDH.n74 9.3005
R5337 VDDH.n635 VDDH.n634 9.3005
R5338 VDDH.n108 VDDH.n107 9.3005
R5339 VDDH.n109 VDDH.n108 9.3005
R5340 VDDH.n95 VDDH.n94 9.3005
R5341 VDDH.n94 VDDH.n93 9.3005
R5342 VDDH.n111 VDDH.n110 9.3005
R5343 VDDH.n106 VDDH.n85 9.3005
R5344 VDDH.n105 VDDH.n104 9.3005
R5345 VDDH.n90 VDDH.n86 9.3005
R5346 VDDH.n645 VDDH.n644 9.3005
R5347 VDDH.n644 VDDH.n643 9.3005
R5348 VDDH.n66 VDDH.n65 9.3005
R5349 VDDH.n67 VDDH.n66 9.3005
R5350 VDDH.n55 VDDH.n54 9.3005
R5351 VDDH.n56 VDDH.n55 9.3005
R5352 VDDH.n658 VDDH.n657 9.3005
R5353 VDDH.n657 VDDH.n656 9.3005
R5354 VDDH.n647 VDDH.n646 9.3005
R5355 VDDH.n648 VDDH.n68 9.3005
R5356 VDDH.n649 VDDH.n49 9.3005
R5357 VDDH.n61 VDDH.n60 9.3005
R5358 VDDH.n59 VDDH.n57 9.3005
R5359 VDDH.n52 VDDH.n51 9.3005
R5360 VDDH.n53 VDDH.n40 9.3005
R5361 VDDH.n655 VDDH.n654 9.3005
R5362 VDDH.n39 VDDH.n37 9.3005
R5363 VDDH.n639 VDDH.n638 9.3005
R5364 VDDH.n642 VDDH.n641 9.3005
R5365 VDDH.n72 VDDH.n70 9.3005
R5366 VDDH.n332 VDDH.n331 9.2505
R5367 VDDH.t59 VDDH.n332 9.2505
R5368 VDDH.n339 VDDH.n338 9.2505
R5369 VDDH.n338 VDDH.t54 9.2505
R5370 VDDH.n334 VDDH.n333 9.2505
R5371 VDDH.n333 VDDH.t59 9.2505
R5372 VDDH.n337 VDDH.n336 9.2505
R5373 VDDH.t54 VDDH.n337 9.2505
R5374 VDDH.t12 VDDH.n279 8.13045
R5375 VDDH.n672 VDDH.t44 7.4369
R5376 VDDH.n704 VDDH.n5 7.11588
R5377 VDDH.n525 VDDH.n376 7.1155
R5378 VDDH.n31 VDDH.n30 6.85235
R5379 VDDH.n671 VDDH.n31 6.85235
R5380 VDDH.n692 VDDH.n691 6.85235
R5381 VDDH.n693 VDDH.n692 6.85235
R5382 VDDH.n703 VDDH 6.4005
R5383 VDDH.n97 VDDH.n96 6.13579
R5384 VDDH.n418 VDDH.n417 5.78175
R5385 VDDH.n423 VDDH.n418 5.78175
R5386 VDDH.n441 VDDH.n440 5.78175
R5387 VDDH.n442 VDDH.n441 5.78175
R5388 VDDH.n420 VDDH.n419 5.78175
R5389 VDDH.n423 VDDH.n420 5.78175
R5390 VDDH.n444 VDDH.n443 5.78175
R5391 VDDH.n443 VDDH.n442 5.78175
R5392 VDDH.n461 VDDH.n460 5.78175
R5393 VDDH.n462 VDDH.n461 5.78175
R5394 VDDH.n455 VDDH.n454 5.78175
R5395 VDDH.n454 VDDH.n453 5.78175
R5396 VDDH.n502 VDDH.n501 5.78175
R5397 VDDH.n501 VDDH.n500 5.78175
R5398 VDDH.n508 VDDH.n507 5.78175
R5399 VDDH.n509 VDDH.n508 5.78175
R5400 VDDH.n464 VDDH.n463 5.78175
R5401 VDDH.n463 VDDH.n462 5.78175
R5402 VDDH.n452 VDDH.n451 5.78175
R5403 VDDH.n453 VDDH.n452 5.78175
R5404 VDDH.n499 VDDH.n498 5.78175
R5405 VDDH.n500 VDDH.n499 5.78175
R5406 VDDH.n511 VDDH.n510 5.78175
R5407 VDDH.n510 VDDH.n509 5.78175
R5408 VDDH.n475 VDDH.n474 5.78175
R5409 VDDH.n474 VDDH.n473 5.78175
R5410 VDDH.n483 VDDH.n482 5.78175
R5411 VDDH.n484 VDDH.n483 5.78175
R5412 VDDH.n495 VDDH.n494 5.78175
R5413 VDDH.n494 VDDH.n493 5.78175
R5414 VDDH.n517 VDDH.n377 5.78175
R5415 VDDH.n518 VDDH.n517 5.78175
R5416 VDDH.n472 VDDH.n471 5.78175
R5417 VDDH.n473 VDDH.n472 5.78175
R5418 VDDH.n486 VDDH.n485 5.78175
R5419 VDDH.n485 VDDH.n484 5.78175
R5420 VDDH.n492 VDDH.n491 5.78175
R5421 VDDH.n493 VDDH.n492 5.78175
R5422 VDDH.n520 VDDH.n519 5.78175
R5423 VDDH.n519 VDDH.n518 5.78175
R5424 VDDH.n678 VDDH.n677 5.78175
R5425 VDDH.n354 VDDH.n304 5.13939
R5426 VDDH.t178 VDDH.n354 5.13939
R5427 VDDH.n352 VDDH.n313 5.13939
R5428 VDDH.n352 VDDH.t220 5.13939
R5429 VDDH.n356 VDDH.n355 5.13939
R5430 VDDH.n355 VDDH.t178 5.13939
R5431 VDDH.n351 VDDH.n350 5.13939
R5432 VDDH.t220 VDDH.n351 5.13939
R5433 VDDH.t148 VDDH.n15 4.99224
R5434 VDDH.n363 VDDH.n301 4.89462
R5435 VDDH.n697 VDDH.n696 4.89462
R5436 VDDH.n282 VDDH.n276 4.89462
R5437 VDDH.n364 VDDH.n277 4.74409
R5438 VDDH.t24 VDDH.n277 4.74409
R5439 VDDH.n342 VDDH.n341 4.40526
R5440 VDDH.n343 VDDH.n342 4.40526
R5441 VDDH.n346 VDDH.n345 4.40526
R5442 VDDH.n345 VDDH.n344 4.40526
R5443 VDDH.n297 VDDH.n296 4.40526
R5444 VDDH.n298 VDDH.n297 4.40526
R5445 VDDH.n374 VDDH.n29 4.12585
R5446 VDDH.n526 VDDH.n525 3.91654
R5447 VDDH.n547 VDDH 3.7711
R5448 VDDH VDDH.n548 3.7711
R5449 VDDH.n245 VDDH 3.7711
R5450 VDDH VDDH.n158 3.7711
R5451 VDDH.n585 VDDH 3.7711
R5452 VDDH VDDH.n586 3.7711
R5453 VDDH.n157 VDDH 3.7711
R5454 VDDH VDDH.n73 3.7711
R5455 VDDH.n636 VDDH 3.7711
R5456 VDDH VDDH.n526 3.7711
R5457 VDDH.n525 VDDH.n524 3.41321
R5458 VDDH.n688 VDDH.n687 3.38392
R5459 VDDH.n373 VDDH.n372 3.36612
R5460 VDDH.n702 VDDH.n7 3.36414
R5461 VDDH.n279 VDDH.n7 3.36414
R5462 VDDH.n433 VDDH.n432 3.13609
R5463 VDDH.n434 VDDH.n433 3.13609
R5464 VDDH.n436 VDDH.n435 3.13609
R5465 VDDH.n435 VDDH.n434 3.13609
R5466 VDDH.n375 VDDH.n373 3.1255
R5467 VDDH.n20 VDDH.n18 2.93701
R5468 VDDH.n672 VDDH.n18 2.93701
R5469 VDDH.n685 VDDH.n673 2.93701
R5470 VDDH.n673 VDDH.n672 2.93701
R5471 VDDH.n99 VDDH.t211 2.8822
R5472 VDDH.t46 VDDH.n83 2.8822
R5473 VDDH.n115 VDDH.t62 2.8822
R5474 VDDH.n622 VDDH.t30 2.8822
R5475 VDDH.n135 VDDH.t278 2.8822
R5476 VDDH.n140 VDDH.t114 2.8822
R5477 VDDH.n149 VDDH.t100 2.8822
R5478 VDDH.n172 VDDH.t10 2.8822
R5479 VDDH.n188 VDDH.t268 2.8822
R5480 VDDH.t3 VDDH.n167 2.8822
R5481 VDDH.n204 VDDH.t38 2.8822
R5482 VDDH.n571 VDDH.t205 2.8822
R5483 VDDH.n224 VDDH.t49 2.8822
R5484 VDDH.n229 VDDH.t67 2.8822
R5485 VDDH.n522 VDDH 2.73738
R5486 VDDH.n524 VDDH.n522 2.55404
R5487 VDDH.n701 VDDH.n3 2.39269
R5488 VDDH.n685 VDDH.n684 2.25932
R5489 VDDH.n524 VDDH.n523 2.23833
R5490 VDDH.n705 VDDH.n3 1.99425
R5491 VDDH.n699 VDDH.n698 1.66612
R5492 VDDH.n96 VDDH.n95 1.60272
R5493 VDDH.n344 VDDH.n343 1.563
R5494 VDDH.n679 VDDH.n28 1.48331
R5495 VDDH.n637 VDDH 1.47967
R5496 VDDH.n375 VDDH.n374 1.4624
R5497 VDDH.n706 VDDH.n705 1.3755
R5498 VDDH.n688 VDDH.n11 1.19112
R5499 VDDH.n681 VDDH.n10 1.163
R5500 VDDH.n698 VDDH.n697 1.163
R5501 VDDH.n689 VDDH.n688 1.14843
R5502 VDDH.n701 VDDH.n700 1.13331
R5503 VDDH.n679 VDDH.n11 1.08019
R5504 VDDH.n293 VDDH.n291 0.985808
R5505 VDDH.n368 VDDH.n366 0.947451
R5506 VDDH.n376 VDDH.n272 0.914875
R5507 VDDH.n294 VDDH.n285 0.873938
R5508 VDDH.n637 VDDH.n636 0.8605
R5509 VDDH.n362 VDDH.n361 0.816125
R5510 VDDH.n362 VDDH.n0 0.816125
R5511 VDDH.n365 VDDH.n275 0.753625
R5512 VDDH.n687 VDDH.n28 0.6255
R5513 VDDH.n363 VDDH.n362 0.6205
R5514 VDDH.n276 VDDH.n22 0.6205
R5515 VDDH.n636 VDDH.n73 0.61925
R5516 VDDH.n157 VDDH.n73 0.61925
R5517 VDDH.n586 VDDH.n157 0.61925
R5518 VDDH.n586 VDDH.n585 0.61925
R5519 VDDH.n585 VDDH.n158 0.61925
R5520 VDDH.n245 VDDH.n158 0.61925
R5521 VDDH.n548 VDDH.n245 0.61925
R5522 VDDH.n548 VDDH.n547 0.61925
R5523 VDDH.n700 VDDH.n699 0.61925
R5524 VDDH VDDH.n637 0.617892
R5525 VDDH.n359 VDDH.n272 0.571125
R5526 VDDH.n547 VDDH 0.56425
R5527 VDDH.n302 VDDH.n275 0.534794
R5528 VDDH.n667 VDDH.n666 0.517167
R5529 VDDH.n661 VDDH.n34 0.517167
R5530 VDDH.n64 VDDH.n63 0.517167
R5531 VDDH.n285 VDDH.n27 0.516125
R5532 VDDH.n376 VDDH.n375 0.475677
R5533 VDDH.n360 VDDH.n359 0.475145
R5534 VDDH.n699 VDDH.n10 0.40675
R5535 VDDH.n705 VDDH.n704 0.3725
R5536 VDDH.n374 VDDH.n30 0.358192
R5537 VDDH.n691 VDDH.n690 0.358192
R5538 VDDH.n680 VDDH.n679 0.3005
R5539 VDDH.n372 VDDH.n22 0.300179
R5540 VDDH.n293 VDDH.n292 0.255835
R5541 VDDH.n285 VDDH.n284 0.255835
R5542 VDDH.n366 VDDH.n273 0.255835
R5543 VDDH.n275 VDDH.n274 0.255835
R5544 VDDH.n371 VDDH.n272 0.251034
R5545 VDDH.n706 VDDH.n0 0.241125
R5546 VDDH.n365 VDDH.n364 0.238962
R5547 VDDH.n368 VDDH.n367 0.227634
R5548 VDDH.n295 VDDH.n294 0.227329
R5549 VDDH.n372 VDDH.n371 0.226462
R5550 VDDH.n36 VDDH.n35 0.218612
R5551 VDDH.n665 VDDH.n664 0.218612
R5552 VDDH.n663 VDDH.n662 0.218612
R5553 VDDH.n660 VDDH.n659 0.218612
R5554 VDDH.n690 VDDH.n22 0.214709
R5555 VDDH.n686 VDDH.n29 0.205663
R5556 VDDH VDDH.n233 0.195324
R5557 VDDH VDDH.n241 0.195324
R5558 VDDH VDDH.n546 0.195324
R5559 VDDH.n527 VDDH 0.195324
R5560 VDDH.n35 VDDH.n29 0.190551
R5561 VDDH.n27 VDDH.n26 0.185122
R5562 VDDH.n702 VDDH.n701 0.172722
R5563 VDDH.n291 VDDH.n286 0.168945
R5564 VDDH.n700 VDDH.n9 0.168674
R5565 VDDH.n3 VDDH.n2 0.168674
R5566 VDDH.n290 VDDH.n288 0.168674
R5567 VDDH.n366 VDDH.n365 0.166125
R5568 VDDH.n289 VDDH.n0 0.159794
R5569 VDDH.n291 VDDH.n290 0.153097
R5570 VDDH.n373 VDDH.n20 0.152959
R5571 VDDH.n686 VDDH.n685 0.152959
R5572 VDDH.n664 VDDH 0.145908
R5573 VDDH.n659 VDDH 0.145908
R5574 VDDH.n666 VDDH.n36 0.129327
R5575 VDDH.n662 VDDH.n661 0.129327
R5576 VDDH VDDH.n635 0.1255
R5577 VDDH.n617 VDDH 0.1255
R5578 VDDH.n602 VDDH 0.1255
R5579 VDDH VDDH.n156 0.1255
R5580 VDDH VDDH.n584 0.1255
R5581 VDDH.n566 VDDH 0.1255
R5582 VDDH VDDH.n663 0.108918
R5583 VDDH.n290 VDDH.n289 0.105208
R5584 VDDH.n370 VDDH.n369 0.105208
R5585 VDDH.n303 VDDH.n302 0.105208
R5586 VDDH.n666 VDDH.n665 0.0897857
R5587 VDDH.n661 VDDH.n660 0.0897857
R5588 VDDH.n369 VDDH.n368 0.086539
R5589 VDDH.n690 VDDH.n689 0.0865043
R5590 VDDH.n689 VDDH.n27 0.078625
R5591 VDDH.n526 VDDH 0.0555
R5592 VDDH.n106 VDDH.n105 0.047375
R5593 VDDH.n635 VDDH.n74 0.047375
R5594 VDDH.n124 VDDH.n123 0.047375
R5595 VDDH.n617 VDDH.n616 0.047375
R5596 VDDH.n611 VDDH.n130 0.047375
R5597 VDDH.n602 VDDH.n601 0.047375
R5598 VDDH.n591 VDDH.n590 0.047375
R5599 VDDH.n185 VDDH.n156 0.047375
R5600 VDDH.n195 VDDH.n194 0.047375
R5601 VDDH.n584 VDDH.n159 0.047375
R5602 VDDH.n213 VDDH.n212 0.047375
R5603 VDDH.n566 VDDH.n565 0.047375
R5604 VDDH.n560 VDDH.n219 0.047375
R5605 VDDH.n552 VDDH.n233 0.047375
R5606 VDDH.n259 VDDH.n241 0.047375
R5607 VDDH.n546 VDDH.n247 0.047375
R5608 VDDH.n527 VDDH.n266 0.047375
R5609 VDDH.n294 VDDH.n293 0.0458125
R5610 VDDH.n360 VDDH.n303 0.0386493
R5611 VDDH.n27 VDDH.n24 0.0379178
R5612 VDDH.n54 VDDH 0.0363146
R5613 VDDH VDDH.n645 0.0338567
R5614 VDDH.n95 VDDH.n90 0.0322383
R5615 VDDH.n110 VDDH.n107 0.0322383
R5616 VDDH.n631 VDDH.n79 0.0322383
R5617 VDDH.n125 VDDH.n122 0.0322383
R5618 VDDH.n615 VDDH.n128 0.0322383
R5619 VDDH.n143 VDDH.n134 0.0322383
R5620 VDDH.n600 VDDH.n146 0.0322383
R5621 VDDH.n589 VDDH.n155 0.0322383
R5622 VDDH.n184 VDDH.n179 0.0322383
R5623 VDDH.n199 VDDH.n196 0.0322383
R5624 VDDH.n580 VDDH.n164 0.0322383
R5625 VDDH.n214 VDDH.n211 0.0322383
R5626 VDDH.n564 VDDH.n217 0.0322383
R5627 VDDH.n242 VDDH.n223 0.0322383
R5628 VDDH.n551 VDDH.n240 0.0322383
R5629 VDDH.n258 VDDH.n255 0.0322383
R5630 VDDH.n269 VDDH.n250 0.0322383
R5631 VDDH.n533 VDDH.n530 0.0322383
R5632 VDDH.n61 VDDH.n50 0.0282388
R5633 VDDH.n646 VDDH.n69 0.0282388
R5634 VDDH.n638 VDDH.n71 0.0282388
R5635 VDDH VDDH.n706 0.0270625
R5636 VDDH.n64 VDDH 0.0268343
R5637 VDDH.n53 VDDH.n38 0.0257809
R5638 VDDH.n105 VDDH 0.0239375
R5639 VDDH.n123 VDDH 0.0239375
R5640 VDDH VDDH.n611 0.0239375
R5641 VDDH.n591 VDDH 0.0239375
R5642 VDDH.n194 VDDH 0.0239375
R5643 VDDH.n212 VDDH 0.0239375
R5644 VDDH VDDH.n560 0.0239375
R5645 VDDH.n656 VDDH.n37 0.023323
R5646 VDDH.n56 VDDH.n52 0.023323
R5647 VDDH.n67 VDDH.n49 0.023323
R5648 VDDH.n643 VDDH.n70 0.023323
R5649 VDDH.n549 VDDH 0.0205195
R5650 VDDH.n256 VDDH 0.0205195
R5651 VDDH VDDH.n271 0.0205195
R5652 VDDH.n532 VDDH 0.0205195
R5653 VDDH.n93 VDDH.n92 0.0200312
R5654 VDDH.n630 VDDH.n628 0.0200312
R5655 VDDH.n613 VDDH.n612 0.0200312
R5656 VDDH.n598 VDDH.n597 0.0200312
R5657 VDDH.n182 VDDH.n181 0.0200312
R5658 VDDH.n579 VDDH.n577 0.0200312
R5659 VDDH.n562 VDDH.n561 0.0200312
R5660 VDDH.n361 VDDH.n360 0.017691
R5661 VDDH VDDH.n53 0.0173539
R5662 VDDH VDDH.n61 0.0173539
R5663 VDDH.n646 VDDH 0.0173539
R5664 VDDH.n638 VDDH 0.0173539
R5665 VDDH VDDH.n658 0.0161716
R5666 VDDH.n107 VDDH.n106 0.0156367
R5667 VDDH.n109 VDDH 0.0156367
R5668 VDDH.n79 VDDH.n74 0.0156367
R5669 VDDH.n125 VDDH.n124 0.0156367
R5670 VDDH VDDH.n127 0.0156367
R5671 VDDH.n616 VDDH.n615 0.0156367
R5672 VDDH.n143 VDDH.n130 0.0156367
R5673 VDDH VDDH.n145 0.0156367
R5674 VDDH.n601 VDDH.n600 0.0156367
R5675 VDDH.n590 VDDH.n589 0.0156367
R5676 VDDH.n587 VDDH 0.0156367
R5677 VDDH.n185 VDDH.n184 0.0156367
R5678 VDDH.n196 VDDH.n195 0.0156367
R5679 VDDH.n198 VDDH 0.0156367
R5680 VDDH.n164 VDDH.n159 0.0156367
R5681 VDDH.n214 VDDH.n213 0.0156367
R5682 VDDH VDDH.n216 0.0156367
R5683 VDDH.n565 VDDH.n564 0.0156367
R5684 VDDH.n242 VDDH.n219 0.0156367
R5685 VDDH VDDH.n244 0.0156367
R5686 VDDH.n552 VDDH.n551 0.0156367
R5687 VDDH.n259 VDDH.n258 0.0156367
R5688 VDDH.n269 VDDH.n247 0.0156367
R5689 VDDH.n530 VDDH.n266 0.0156367
R5690 VDDH.n656 VDDH.n655 0.0113848
R5691 VDDH.n57 VDDH.n56 0.0113848
R5692 VDDH.n68 VDDH.n67 0.0113848
R5693 VDDH.n643 VDDH.n642 0.0113848
R5694 VDDH.n9 VDDH.n8 0.00995724
R5695 VDDH.n2 VDDH.n1 0.00995724
R5696 VDDH.n288 VDDH.n287 0.00995724
R5697 VDDH.n24 VDDH.n23 0.00995724
R5698 VDDH.n26 VDDH.n25 0.00995724
R5699 VDDH.n655 VDDH.n38 0.00892697
R5700 VDDH.n65 VDDH.n64 0.00752247
R5701 VDDH.n57 VDDH.n50 0.0064691
R5702 VDDH.n69 VDDH.n68 0.0064691
R5703 VDDH.n642 VDDH.n71 0.0064691
R5704 VDDH.n687 VDDH.n686 0.00457609
R5705 VDDH.n93 VDDH.n90 0.00391797
R5706 VDDH.n110 VDDH.n109 0.00391797
R5707 VDDH.n631 VDDH.n630 0.00391797
R5708 VDDH.n127 VDDH.n122 0.00391797
R5709 VDDH.n613 VDDH.n128 0.00391797
R5710 VDDH.n145 VDDH.n134 0.00391797
R5711 VDDH.n598 VDDH.n146 0.00391797
R5712 VDDH.n587 VDDH.n155 0.00391797
R5713 VDDH.n182 VDDH.n179 0.00391797
R5714 VDDH.n199 VDDH.n198 0.00391797
R5715 VDDH.n580 VDDH.n579 0.00391797
R5716 VDDH.n216 VDDH.n211 0.00391797
R5717 VDDH.n562 VDDH.n217 0.00391797
R5718 VDDH.n244 VDDH.n223 0.00391797
R5719 VDDH.n549 VDDH.n240 0.00391797
R5720 VDDH.n256 VDDH.n255 0.00391797
R5721 VDDH.n271 VDDH.n250 0.00391797
R5722 VDDH.n533 VDDH.n532 0.00391797
R5723 VDDH.n658 VDDH.n37 0.00295787
R5724 VDDH.n54 VDDH.n52 0.00295787
R5725 VDDH.n65 VDDH.n49 0.00295787
R5726 VDDH.n645 VDDH.n70 0.00295787
R5727 VDDH.n92 VDDH 0.000988281
R5728 VDDH.n628 VDDH 0.000988281
R5729 VDDH.n612 VDDH 0.000988281
R5730 VDDH.n597 VDDH 0.000988281
R5731 VDDH.n181 VDDH 0.000988281
R5732 VDDH.n577 VDDH 0.000988281
R5733 VDDH.n561 VDDH 0.000988281
R5734 top_segment_4_1.bb3.n2 top_segment_4_1.bb3.n1 863.124
R5735 top_segment_4_1.bb3.n1 top_segment_4_1.bb3.n0 585
R5736 top_segment_4_1.bb3 top_segment_4_1.bb3.t1 495.469
R5737 top_segment_4_1.bb3 top_segment_4_1.bb3.t0 291.983
R5738 top_segment_4_1.bb3.t0 top_segment_4_1.bb3.n25 285
R5739 top_segment_4_1.bb3.n3 top_segment_4_1.bb3.t11 217.555
R5740 top_segment_4_1.bb3.n5 top_segment_4_1.bb3.t17 217.555
R5741 top_segment_4_1.bb3.n7 top_segment_4_1.bb3.t10 216.893
R5742 top_segment_4_1.bb3.n8 top_segment_4_1.bb3.t12 216.893
R5743 top_segment_4_1.bb3.n9 top_segment_4_1.bb3.t5 216.893
R5744 top_segment_4_1.bb3.n10 top_segment_4_1.bb3.t21 216.893
R5745 top_segment_4_1.bb3.n6 top_segment_4_1.bb3.t6 216.893
R5746 top_segment_4_1.bb3.n5 top_segment_4_1.bb3.t2 216.893
R5747 top_segment_4_1.bb3.n19 top_segment_4_1.bb3.t14 213.218
R5748 top_segment_4_1.bb3.n14 top_segment_4_1.bb3.t9 213.218
R5749 top_segment_4_1.bb3.n18 top_segment_4_1.bb3.t18 212.554
R5750 top_segment_4_1.bb3.n17 top_segment_4_1.bb3.t15 212.554
R5751 top_segment_4_1.bb3.n16 top_segment_4_1.bb3.t8 212.554
R5752 top_segment_4_1.bb3.n15 top_segment_4_1.bb3.t19 212.554
R5753 top_segment_4_1.bb3.n14 top_segment_4_1.bb3.t16 212.554
R5754 top_segment_4_1.bb3.n4 top_segment_4_1.bb3.t20 212.393
R5755 top_segment_4_1.bb3.n12 top_segment_4_1.bb3.t7 212.393
R5756 top_segment_4_1.bb3.n20 top_segment_4_1.bb3.t3 208.054
R5757 top_segment_4_1.bb3.n23 top_segment_4_1.bb3.n22 152
R5758 top_segment_4_1.bb3.n1 top_segment_4_1.bb3.t1 140.738
R5759 top_segment_4_1.bb3.n22 top_segment_4_1.bb3.t4 114.031
R5760 top_segment_4_1.bb3.n22 top_segment_4_1.bb3.t13 81.5883
R5761 top_segment_4_1.bb3 top_segment_4_1.bb3.n21 29.1651
R5762 top_segment_4_1.bb3.n13 top_segment_4_1.bb3.n4 23.6838
R5763 top_segment_4_1.bb3.n21 top_segment_4_1.bb3.n13 18.9547
R5764 top_segment_4_1.bb3.n23 top_segment_4_1.bb3 16.7132
R5765 top_segment_4_1.bb3.n21 top_segment_4_1.bb3.n20 14.013
R5766 top_segment_4_1.bb3.n13 top_segment_4_1.bb3.n12 13.9942
R5767 top_segment_4_1.bb3.n24 top_segment_4_1.bb3 13.7979
R5768 top_segment_4_1.bb3 top_segment_4_1.bb3.n24 13.1884
R5769 top_segment_4_1.bb3 top_segment_4_1.bb3.n25 12.4126
R5770 top_segment_4_1.bb3.n2 top_segment_4_1.bb3 11.6369
R5771 top_segment_4_1.bb3.n0 top_segment_4_1.bb3 10.1408
R5772 top_segment_4_1.bb3.n4 top_segment_4_1.bb3.n3 4.5005
R5773 top_segment_4_1.bb3.n12 top_segment_4_1.bb3.n11 4.5005
R5774 top_segment_4_1.bb3.n20 top_segment_4_1.bb3.n19 4.5005
R5775 top_segment_4_1.bb3.n0 top_segment_4_1.bb3 2.16154
R5776 top_segment_4_1.bb3.n24 top_segment_4_1.bb3 2.16154
R5777 top_segment_4_1.bb3.n25 top_segment_4_1.bb3 1.93989
R5778 top_segment_4_1.bb3 top_segment_4_1.bb3.n23 1.16414
R5779 top_segment_4_1.bb3 top_segment_4_1.bb3.n2 0.665435
R5780 top_segment_4_1.bb3.n6 top_segment_4_1.bb3.n5 0.663962
R5781 top_segment_4_1.bb3.n11 top_segment_4_1.bb3.n6 0.663962
R5782 top_segment_4_1.bb3.n11 top_segment_4_1.bb3.n10 0.663962
R5783 top_segment_4_1.bb3.n10 top_segment_4_1.bb3.n9 0.663962
R5784 top_segment_4_1.bb3.n9 top_segment_4_1.bb3.n8 0.663962
R5785 top_segment_4_1.bb3.n8 top_segment_4_1.bb3.n7 0.663962
R5786 top_segment_4_1.bb3.n15 top_segment_4_1.bb3.n14 0.663962
R5787 top_segment_4_1.bb3.n17 top_segment_4_1.bb3.n16 0.663962
R5788 top_segment_4_1.bb3.n18 top_segment_4_1.bb3.n17 0.663962
R5789 top_segment_4_1.bb3.n19 top_segment_4_1.bb3.n18 0.663962
R5790 top_segment_4_1.bb3.n24 top_segment_4_1.bb3 0.582318
R5791 top_segment_4_1.bb3.n16 top_segment_4_1.bb3 0.541365
R5792 top_segment_4_1.bb3.n3 top_segment_4_1.bb3 0.310596
R5793 top_segment_4_1.bb3.n7 top_segment_4_1.bb3 0.293769
R5794 top_segment_4_1.bb3 top_segment_4_1.bb3.n15 0.123096
R5795 a_15714_6674.t0 a_15714_6674.n2 672.764
R5796 a_15714_6674.n0 a_15714_6674.t3 670.999
R5797 a_15714_6674.n0 a_15714_6674.t4 666.655
R5798 a_15714_6674.n2 a_15714_6674.t1 666.275
R5799 a_15714_6674.n1 a_15714_6674.t2 666.275
R5800 a_15714_6674.n2 a_15714_6674.n1 6.63383
R5801 a_15714_6674.n1 a_15714_6674.n0 2.23175
R5802 a_18769_7938.n0 a_18769_7938.t1 671.744
R5803 a_18769_7938.n0 a_18769_7938.t2 671.292
R5804 a_18769_7938.t0 a_18769_7938.n0 665.34
R5805 top_segment_2_0.rseg_2_v3_0.v42.t0 top_segment_2_0.rseg_2_v3_0.v42.n0 240.321
R5806 top_segment_2_0.rseg_2_v3_0.v42.n0 top_segment_2_0.rseg_2_v3_0.v42.t2 10.7966
R5807 top_segment_2_0.rseg_2_v3_0.v42.n0 top_segment_2_0.rseg_2_v3_0.v42.t1 10.6741
R5808 top_segment_2_0.rseg_2_v3_0.v41.t0 top_segment_2_0.rseg_2_v3_0.v41.n0 240.44
R5809 top_segment_2_0.rseg_2_v3_0.v41.n0 top_segment_2_0.rseg_2_v3_0.v41.t1 10.7488
R5810 top_segment_2_0.rseg_2_v3_0.v41.n0 top_segment_2_0.rseg_2_v3_0.v41.t2 10.6292
R5811 top_segment_2_0.DEC2[2].n0 top_segment_2_0.DEC2[2].t0 334.788
R5812 top_segment_2_0.DEC2[2].n11 top_segment_2_0.DEC2[2].t6 213.218
R5813 top_segment_2_0.DEC2[2].n16 top_segment_2_0.DEC2[2].t8 213.218
R5814 top_segment_2_0.DEC2[2].n5 top_segment_2_0.DEC2[2].t22 213.218
R5815 top_segment_2_0.DEC2[2] top_segment_2_0.DEC2[2].t3 212.887
R5816 top_segment_2_0.DEC2[2].n11 top_segment_2_0.DEC2[2].t17 212.554
R5817 top_segment_2_0.DEC2[2].n12 top_segment_2_0.DEC2[2].t4 212.554
R5818 top_segment_2_0.DEC2[2].n13 top_segment_2_0.DEC2[2].t23 212.554
R5819 top_segment_2_0.DEC2[2].n14 top_segment_2_0.DEC2[2].t19 212.554
R5820 top_segment_2_0.DEC2[2].n15 top_segment_2_0.DEC2[2].t14 212.554
R5821 top_segment_2_0.DEC2[2].n10 top_segment_2_0.DEC2[2].t20 212.554
R5822 top_segment_2_0.DEC2[2].n9 top_segment_2_0.DEC2[2].t5 212.554
R5823 top_segment_2_0.DEC2[2].n8 top_segment_2_0.DEC2[2].t11 212.554
R5824 top_segment_2_0.DEC2[2].n7 top_segment_2_0.DEC2[2].t21 212.554
R5825 top_segment_2_0.DEC2[2].n6 top_segment_2_0.DEC2[2].t18 212.554
R5826 top_segment_2_0.DEC2[2].n5 top_segment_2_0.DEC2[2].t13 212.554
R5827 top_segment_2_0.DEC2[2].n4 top_segment_2_0.DEC2[2].t9 208.054
R5828 top_segment_2_0.DEC2[2].n18 top_segment_2_0.DEC2[2].t7 208.054
R5829 top_segment_2_0.DEC2[2].n17 top_segment_2_0.DEC2[2].t10 208.054
R5830 top_segment_2_0.DEC2[2].n22 top_segment_2_0.DEC2[2].n21 152
R5831 top_segment_2_0.DEC2[2].n2 top_segment_2_0.DEC2[2].t2 126.27
R5832 top_segment_2_0.DEC2[2].n2 top_segment_2_0.DEC2[2].t15 125.558
R5833 top_segment_2_0.DEC2[2].n1 top_segment_2_0.DEC2[2].t24 121.127
R5834 top_segment_2_0.DEC2[2].n21 top_segment_2_0.DEC2[2].t12 114.031
R5835 top_segment_2_0.DEC2[2].n0 top_segment_2_0.DEC2[2].t1 87.8063
R5836 top_segment_2_0.DEC2[2].n21 top_segment_2_0.DEC2[2].t16 81.5883
R5837 top_segment_2_0.DEC2[2].n20 top_segment_2_0.DEC2[2].n4 39.4293
R5838 top_segment_2_0.DEC2[2] top_segment_2_0.DEC2[2].n20 28.2979
R5839 top_segment_2_0.DEC2[2].n23 top_segment_2_0.DEC2[2] 15.1345
R5840 top_segment_2_0.DEC2[2].n20 top_segment_2_0.DEC2[2] 13.0029
R5841 top_segment_2_0.DEC2[2] top_segment_2_0.DEC2[2].n22 11.4706
R5842 top_segment_2_0.DEC2[2].n3 top_segment_2_0.DEC2[2].n2 5.73592
R5843 top_segment_2_0.DEC2[2] top_segment_2_0.DEC2[2].n3 5.388
R5844 top_segment_2_0.DEC2[2].n4 top_segment_2_0.DEC2[2] 4.83223
R5845 top_segment_2_0.DEC2[2].n17 top_segment_2_0.DEC2[2].n16 4.5005
R5846 top_segment_2_0.DEC2[2].n19 top_segment_2_0.DEC2[2].n18 4.5005
R5847 top_segment_2_0.DEC2[2].n22 top_segment_2_0.DEC2[2] 4.48881
R5848 top_segment_2_0.DEC2[2].n18 top_segment_2_0.DEC2[2].n17 2.59281
R5849 top_segment_2_0.DEC2[2] top_segment_2_0.DEC2[2].n23 1.02758
R5850 top_segment_2_0.DEC2[2].n23 top_segment_2_0.DEC2[2] 0.7755
R5851 top_segment_2_0.DEC2[2].n16 top_segment_2_0.DEC2[2].n15 0.663962
R5852 top_segment_2_0.DEC2[2].n15 top_segment_2_0.DEC2[2].n14 0.663962
R5853 top_segment_2_0.DEC2[2].n14 top_segment_2_0.DEC2[2].n13 0.663962
R5854 top_segment_2_0.DEC2[2].n13 top_segment_2_0.DEC2[2].n12 0.663962
R5855 top_segment_2_0.DEC2[2].n12 top_segment_2_0.DEC2[2].n11 0.663962
R5856 top_segment_2_0.DEC2[2].n6 top_segment_2_0.DEC2[2].n5 0.663962
R5857 top_segment_2_0.DEC2[2].n7 top_segment_2_0.DEC2[2].n6 0.663962
R5858 top_segment_2_0.DEC2[2].n8 top_segment_2_0.DEC2[2].n7 0.663962
R5859 top_segment_2_0.DEC2[2].n9 top_segment_2_0.DEC2[2].n8 0.663962
R5860 top_segment_2_0.DEC2[2].n10 top_segment_2_0.DEC2[2].n9 0.663962
R5861 top_segment_2_0.DEC2[2].n19 top_segment_2_0.DEC2[2].n10 0.663962
R5862 top_segment_2_0.DEC2[2].n1 top_segment_2_0.DEC2[2].n0 0.322615
R5863 top_segment_2_0.DEC2[2] top_segment_2_0.DEC2[2].n19 0.291365
R5864 top_segment_2_0.DEC2[2].n3 top_segment_2_0.DEC2[2].n1 0.177583
R5865 a_41529_17118.t0 a_41529_17118.t1 65.941
R5866 a_41787_17118.t0 a_41787_17118.t1 65.941
R5867 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t5 231.017
R5868 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t6 230.155
R5869 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t11 229.369
R5870 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t12 229.369
R5871 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t17 229.369
R5872 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t9 229.369
R5873 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t13 228.649
R5874 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n22 203.923
R5875 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t16 158.716
R5876 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n14 157.927
R5877 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t7 157.856
R5878 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t14 157.07
R5879 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t15 157.07
R5880 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t10 157.07
R5881 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t4 157.07
R5882 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t8 156.35
R5883 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n2 156.268
R5884 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n5 153.423
R5885 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n15 152
R5886 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n12 152
R5887 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n9 152
R5888 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n3 152
R5889 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n0 101.49
R5890 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 53.8309
R5891 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n19 43.993
R5892 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t0 26.5955
R5893 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t1 26.5955
R5894 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t2 24.9236
R5895 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t3 24.9236
R5896 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n10 18.4368
R5897 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n4 16.4183
R5898 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n6 14.4998
R5899 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n16 13.1513
R5900 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 13.0565
R5901 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n13 11.3143
R5902 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 10.7525
R5903 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n17 9.3005
R5904 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 7.11161
R5905 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 6.6565
R5906 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n18 6.60324
R5907 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 5.92643
R5908 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 5.92643
R5909 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n21 5.04292
R5910 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 4.5042
R5911 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n20 4.3525
R5912 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n1 2.5605
R5913 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 2.3045
R5914 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 1.93989
R5915 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 1.43334
R5916 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n8 1.13136
R5917 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n7 1.10597
R5918 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n11 0.699719
R5919 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.529797
R5920 a_41714_2150.t0 a_41714_2150.t1 49.8467
R5921 top_segment_2_0.rseg_2_v3_0.v4.n0 top_segment_2_0.rseg_2_v3_0.v4.t1 239.142
R5922 top_segment_2_0.rseg_2_v3_0.v4.t0 top_segment_2_0.rseg_2_v3_0.v4.n0 10.5871
R5923 top_segment_2_0.rseg_2_v3_0.v4.n0 top_segment_2_0.rseg_2_v3_0.v4.t2 10.5739
R5924 top_segment_2_0.rseg_2_v3_0.v5.n0 top_segment_2_0.rseg_2_v3_0.v5.t2 242.369
R5925 top_segment_2_0.rseg_2_v3_0.v5.t0 top_segment_2_0.rseg_2_v3_0.v5.n0 10.5394
R5926 top_segment_2_0.rseg_2_v3_0.v5.n0 top_segment_2_0.rseg_2_v3_0.v5.t1 10.5285
R5927 top_segment_2_0.DEC2[0].n0 top_segment_2_0.DEC2[0].t0 334.771
R5928 top_segment_2_0.DEC2[0].n12 top_segment_2_0.DEC2[0].t10 213.218
R5929 top_segment_2_0.DEC2[0].n8 top_segment_2_0.DEC2[0].t23 213.218
R5930 top_segment_2_0.DEC2[0].n5 top_segment_2_0.DEC2[0].t21 213.218
R5931 top_segment_2_0.DEC2[0] top_segment_2_0.DEC2[0].t18 212.895
R5932 top_segment_2_0.DEC2[0].n18 top_segment_2_0.DEC2[0].t5 212.554
R5933 top_segment_2_0.DEC2[0].n17 top_segment_2_0.DEC2[0].t2 212.554
R5934 top_segment_2_0.DEC2[0].n16 top_segment_2_0.DEC2[0].t12 212.554
R5935 top_segment_2_0.DEC2[0].n15 top_segment_2_0.DEC2[0].t22 212.554
R5936 top_segment_2_0.DEC2[0].n14 top_segment_2_0.DEC2[0].t16 212.554
R5937 top_segment_2_0.DEC2[0].n13 top_segment_2_0.DEC2[0].t13 212.554
R5938 top_segment_2_0.DEC2[0].n12 top_segment_2_0.DEC2[0].t17 212.554
R5939 top_segment_2_0.DEC2[0].n8 top_segment_2_0.DEC2[0].t8 212.554
R5940 top_segment_2_0.DEC2[0].n9 top_segment_2_0.DEC2[0].t4 212.554
R5941 top_segment_2_0.DEC2[0].n10 top_segment_2_0.DEC2[0].t24 212.554
R5942 top_segment_2_0.DEC2[0].n7 top_segment_2_0.DEC2[0].t9 212.554
R5943 top_segment_2_0.DEC2[0].n6 top_segment_2_0.DEC2[0].t19 212.554
R5944 top_segment_2_0.DEC2[0].n5 top_segment_2_0.DEC2[0].t14 212.554
R5945 top_segment_2_0.DEC2[0].n4 top_segment_2_0.DEC2[0].t6 208.054
R5946 top_segment_2_0.DEC2[0].n22 top_segment_2_0.DEC2[0].n21 152
R5947 top_segment_2_0.DEC2[0].n1 top_segment_2_0.DEC2[0].t15 126.278
R5948 top_segment_2_0.DEC2[0].n1 top_segment_2_0.DEC2[0].t7 125.566
R5949 top_segment_2_0.DEC2[0].n2 top_segment_2_0.DEC2[0].t20 125.566
R5950 top_segment_2_0.DEC2[0].n21 top_segment_2_0.DEC2[0].t11 114.031
R5951 top_segment_2_0.DEC2[0].n0 top_segment_2_0.DEC2[0].t1 87.8568
R5952 top_segment_2_0.DEC2[0].n21 top_segment_2_0.DEC2[0].t3 81.5883
R5953 top_segment_2_0.DEC2[0] top_segment_2_0.DEC2[0].n20 43.6567
R5954 top_segment_2_0.DEC2[0].n20 top_segment_2_0.DEC2[0].n4 20.963
R5955 top_segment_2_0.DEC2[0].n20 top_segment_2_0.DEC2[0].n19 19.2422
R5956 top_segment_2_0.DEC2[0].n23 top_segment_2_0.DEC2[0] 15.6308
R5957 top_segment_2_0.DEC2[0] top_segment_2_0.DEC2[0].n22 11.4706
R5958 top_segment_2_0.DEC2[0].n19 top_segment_2_0.DEC2[0] 7.31717
R5959 top_segment_2_0.DEC2[0].n19 top_segment_2_0.DEC2[0].n11 7.0755
R5960 top_segment_2_0.DEC2[0] top_segment_2_0.DEC2[0].n3 5.04008
R5961 top_segment_2_0.DEC2[0].n4 top_segment_2_0.DEC2[0] 4.82262
R5962 top_segment_2_0.DEC2[0].n3 top_segment_2_0.DEC2[0].n2 4.68383
R5963 top_segment_2_0.DEC2[0].n22 top_segment_2_0.DEC2[0] 4.48881
R5964 top_segment_2_0.DEC2[0] top_segment_2_0.DEC2[0].n23 1.01508
R5965 top_segment_2_0.DEC2[0].n3 top_segment_2_0.DEC2[0].n0 0.876942
R5966 top_segment_2_0.DEC2[0].n23 top_segment_2_0.DEC2[0] 0.7755
R5967 top_segment_2_0.DEC2[0].n2 top_segment_2_0.DEC2[0].n1 0.713
R5968 top_segment_2_0.DEC2[0].n13 top_segment_2_0.DEC2[0].n12 0.663962
R5969 top_segment_2_0.DEC2[0].n14 top_segment_2_0.DEC2[0].n13 0.663962
R5970 top_segment_2_0.DEC2[0].n15 top_segment_2_0.DEC2[0].n14 0.663962
R5971 top_segment_2_0.DEC2[0].n16 top_segment_2_0.DEC2[0].n15 0.663962
R5972 top_segment_2_0.DEC2[0].n17 top_segment_2_0.DEC2[0].n16 0.663962
R5973 top_segment_2_0.DEC2[0].n18 top_segment_2_0.DEC2[0].n17 0.663962
R5974 top_segment_2_0.DEC2[0].n10 top_segment_2_0.DEC2[0].n9 0.663962
R5975 top_segment_2_0.DEC2[0].n9 top_segment_2_0.DEC2[0].n8 0.663962
R5976 top_segment_2_0.DEC2[0].n6 top_segment_2_0.DEC2[0].n5 0.663962
R5977 top_segment_2_0.DEC2[0].n7 top_segment_2_0.DEC2[0].n6 0.663962
R5978 top_segment_2_0.DEC2[0].n11 top_segment_2_0.DEC2[0].n10 0.312199
R5979 top_segment_2_0.DEC2[0].n11 top_segment_2_0.DEC2[0].n7 0.312199
R5980 top_segment_2_0.DEC2[0] top_segment_2_0.DEC2[0].n18 0.254667
R5981 a_28603_6674.n2 a_28603_6674.t4 246.061
R5982 a_28603_6674.n0 a_28603_6674.t2 240.989
R5983 a_28603_6674.n0 a_28603_6674.t1 240.81
R5984 a_28603_6674.n1 a_28603_6674.t3 238.775
R5985 a_28603_6674.t0 a_28603_6674.n2 238.775
R5986 a_28603_6674.n2 a_28603_6674.n1 6.788
R5987 a_28603_6674.n1 a_28603_6674.n0 4.54842
R5988 top_segment_1_0.rseg_1_v3_1.v9 top_segment_1_0.rseg_1_v3_1.v9.t1 249.345
R5989 top_segment_1_0.rseg_1_v3_1.v9.n0 top_segment_1_0.rseg_1_v3_1.v9.t2 10.5773
R5990 top_segment_1_0.rseg_1_v3_1.v9.n0 top_segment_1_0.rseg_1_v3_1.v9.t0 10.5739
R5991 top_segment_1_0.rseg_1_v3_1.v9 top_segment_1_0.rseg_1_v3_1.v9.n0 4.18158
R5992 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t1 673.212
R5993 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t0 10.7613
R5994 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t2 10.7113
R5995 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.n0 2.72292
R5996 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t2 673.572
R5997 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t1 10.7178
R5998 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.t0 10.6903
R5999 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54.n0 3.41701
R6000 top_segment_2_0.DEC0[0].n17 top_segment_2_0.DEC0[0].t1 334.771
R6001 top_segment_2_0.DEC0[0].n5 top_segment_2_0.DEC0[0].t2 213.218
R6002 top_segment_2_0.DEC0[0].n5 top_segment_2_0.DEC0[0].t9 212.554
R6003 top_segment_2_0.DEC0[0].n6 top_segment_2_0.DEC0[0].t18 212.554
R6004 top_segment_2_0.DEC0[0].n7 top_segment_2_0.DEC0[0].t3 212.554
R6005 top_segment_2_0.DEC0[0].n8 top_segment_2_0.DEC0[0].t11 212.554
R6006 top_segment_2_0.DEC0[0].n9 top_segment_2_0.DEC0[0].t10 212.554
R6007 top_segment_2_0.DEC0[0].n10 top_segment_2_0.DEC0[0].t13 212.554
R6008 top_segment_2_0.DEC0[0].n11 top_segment_2_0.DEC0[0].t5 212.554
R6009 top_segment_2_0.DEC0[0].n12 top_segment_2_0.DEC0[0].t12 212.554
R6010 top_segment_2_0.DEC0[0].n13 top_segment_2_0.DEC0[0].t19 212.554
R6011 top_segment_2_0.DEC0[0].n14 top_segment_2_0.DEC0[0].t7 212.554
R6012 top_segment_2_0.DEC0[0].n4 top_segment_2_0.DEC0[0].t4 212.554
R6013 top_segment_2_0.DEC0[0].n3 top_segment_2_0.DEC0[0].t15 212.554
R6014 top_segment_2_0.DEC0[0].n2 top_segment_2_0.DEC0[0].t20 212.554
R6015 top_segment_2_0.DEC0[0].n1 top_segment_2_0.DEC0[0].t8 212.554
R6016 top_segment_2_0.DEC0[0].n0 top_segment_2_0.DEC0[0].t16 212.554
R6017 top_segment_2_0.DEC0[0].n16 top_segment_2_0.DEC0[0].t17 208.054
R6018 top_segment_2_0.DEC0[0].n18 top_segment_2_0.DEC0[0].t14 126.278
R6019 top_segment_2_0.DEC0[0].n18 top_segment_2_0.DEC0[0].t21 125.566
R6020 top_segment_2_0.DEC0[0].n19 top_segment_2_0.DEC0[0].t6 125.566
R6021 top_segment_2_0.DEC0[0].n17 top_segment_2_0.DEC0[0].t0 87.8568
R6022 top_segment_2_0.DEC0[0] top_segment_2_0.DEC0[0].n16 62.8505
R6023 top_segment_2_0.DEC0[0] top_segment_2_0.DEC0[0].n20 5.04008
R6024 top_segment_2_0.DEC0[0].n20 top_segment_2_0.DEC0[0].n19 4.68383
R6025 top_segment_2_0.DEC0[0].n16 top_segment_2_0.DEC0[0].n15 4.5005
R6026 top_segment_2_0.DEC0[0].n20 top_segment_2_0.DEC0[0].n17 0.876942
R6027 top_segment_2_0.DEC0[0].n19 top_segment_2_0.DEC0[0].n18 0.713
R6028 top_segment_2_0.DEC0[0].n1 top_segment_2_0.DEC0[0].n0 0.663962
R6029 top_segment_2_0.DEC0[0].n2 top_segment_2_0.DEC0[0].n1 0.663962
R6030 top_segment_2_0.DEC0[0].n3 top_segment_2_0.DEC0[0].n2 0.663962
R6031 top_segment_2_0.DEC0[0].n4 top_segment_2_0.DEC0[0].n3 0.663962
R6032 top_segment_2_0.DEC0[0].n15 top_segment_2_0.DEC0[0].n4 0.663962
R6033 top_segment_2_0.DEC0[0].n15 top_segment_2_0.DEC0[0].n14 0.663962
R6034 top_segment_2_0.DEC0[0].n14 top_segment_2_0.DEC0[0].n13 0.663962
R6035 top_segment_2_0.DEC0[0].n13 top_segment_2_0.DEC0[0].n12 0.663962
R6036 top_segment_2_0.DEC0[0].n12 top_segment_2_0.DEC0[0].n11 0.663962
R6037 top_segment_2_0.DEC0[0].n11 top_segment_2_0.DEC0[0].n10 0.663962
R6038 top_segment_2_0.DEC0[0].n10 top_segment_2_0.DEC0[0].n9 0.663962
R6039 top_segment_2_0.DEC0[0].n9 top_segment_2_0.DEC0[0].n8 0.663962
R6040 top_segment_2_0.DEC0[0].n8 top_segment_2_0.DEC0[0].n7 0.663962
R6041 top_segment_2_0.DEC0[0].n7 top_segment_2_0.DEC0[0].n6 0.663962
R6042 top_segment_2_0.DEC0[0].n6 top_segment_2_0.DEC0[0].n5 0.663962
R6043 top_segment_2_0.DEC0[0].n0 top_segment_2_0.DEC0[0] 0.209635
R6044 a_19094_19162.t0 a_19094_19162.n1 250.803
R6045 a_19094_19162.n0 a_19094_19162.t2 248.238
R6046 a_19094_19162.n1 a_19094_19162.t3 240.714
R6047 a_19094_19162.n0 a_19094_19162.t1 239.833
R6048 a_19094_19162.n1 a_19094_19162.n0 2.56508
R6049 top_segment_2_0.rseg_2_v3_0.v10.n0 top_segment_2_0.rseg_2_v3_0.v10.t2 239.999
R6050 top_segment_2_0.rseg_2_v3_0.v10.t0 top_segment_2_0.rseg_2_v3_0.v10.n0 10.5782
R6051 top_segment_2_0.rseg_2_v3_0.v10.n0 top_segment_2_0.rseg_2_v3_0.v10.t1 10.5739
R6052 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t4 761.467
R6053 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 203.923
R6054 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 101.49
R6055 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t2 26.5955
R6056 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t3 26.5955
R6057 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t0 24.9236
R6058 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t1 24.9236
R6059 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 13.0565
R6060 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 10.7525
R6061 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y 6.6565
R6062 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y 5.04292
R6063 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y 4.3525
R6064 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y 2.5605
R6065 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 1.93989
R6066 a_42781_13270.t0 a_42781_13270.t1 114.052
R6067 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t1 227.856
R6068 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n2 152.333
R6069 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t2 140.382
R6070 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t3 114.031
R6071 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t0 83.3993
R6072 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.t4 81.5883
R6073 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n3 14.4422
R6074 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n1 7.56882
R6075 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n0 5.08175
R6076 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R6077 a_42271_12320.t0 a_42271_12320.t1 55.3905
R6078 a_42245_11724.t0 a_42245_11724.n0 228.04
R6079 a_42245_11724.n0 a_42245_11724.t2 145.648
R6080 a_42245_11724.n0 a_42245_11724.t1 83.2159
R6081 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[4] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t3 753.758
R6082 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t5 230.576
R6083 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t0 216.44
R6084 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t4 158.275
R6085 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 153.661
R6086 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 152
R6087 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 28.99
R6088 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t2 24.9236
R6089 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t1 24.9236
R6090 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[4] 18.1258
R6091 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 11.7913
R6092 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 10.7516
R6093 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 10.238
R6094 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.A 6.66717
R6095 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[4] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[4] 0.7505
R6096 a_42781_9310.t0 a_42781_9310.t1 114.052
R6097 top_segment_2_0.DEC2[3].n0 top_segment_2_0.DEC2[3].t1 334.822
R6098 top_segment_2_0.DEC2[3].n11 top_segment_2_0.DEC2[3].t7 213.218
R6099 top_segment_2_0.DEC2[3].n16 top_segment_2_0.DEC2[3].t14 213.218
R6100 top_segment_2_0.DEC2[3].n5 top_segment_2_0.DEC2[3].t13 213.218
R6101 top_segment_2_0.DEC2[3] top_segment_2_0.DEC2[3].t11 212.864
R6102 top_segment_2_0.DEC2[3].n11 top_segment_2_0.DEC2[3].t20 212.554
R6103 top_segment_2_0.DEC2[3].n12 top_segment_2_0.DEC2[3].t3 212.554
R6104 top_segment_2_0.DEC2[3].n13 top_segment_2_0.DEC2[3].t24 212.554
R6105 top_segment_2_0.DEC2[3].n14 top_segment_2_0.DEC2[3].t21 212.554
R6106 top_segment_2_0.DEC2[3].n15 top_segment_2_0.DEC2[3].t4 212.554
R6107 top_segment_2_0.DEC2[3].n10 top_segment_2_0.DEC2[3].t23 212.554
R6108 top_segment_2_0.DEC2[3].n9 top_segment_2_0.DEC2[3].t19 212.554
R6109 top_segment_2_0.DEC2[3].n8 top_segment_2_0.DEC2[3].t18 212.554
R6110 top_segment_2_0.DEC2[3].n7 top_segment_2_0.DEC2[3].t15 212.554
R6111 top_segment_2_0.DEC2[3].n6 top_segment_2_0.DEC2[3].t12 212.554
R6112 top_segment_2_0.DEC2[3].n5 top_segment_2_0.DEC2[3].t10 212.554
R6113 top_segment_2_0.DEC2[3].n4 top_segment_2_0.DEC2[3].t22 208.054
R6114 top_segment_2_0.DEC2[3].n18 top_segment_2_0.DEC2[3].t2 208.054
R6115 top_segment_2_0.DEC2[3].n17 top_segment_2_0.DEC2[3].t17 208.054
R6116 top_segment_2_0.DEC2[3].n22 top_segment_2_0.DEC2[3].n21 152
R6117 top_segment_2_0.DEC2[3].n1 top_segment_2_0.DEC2[3].t8 126.27
R6118 top_segment_2_0.DEC2[3].n2 top_segment_2_0.DEC2[3].t9 125.558
R6119 top_segment_2_0.DEC2[3].n1 top_segment_2_0.DEC2[3].t6 125.558
R6120 top_segment_2_0.DEC2[3].n21 top_segment_2_0.DEC2[3].t16 114.031
R6121 top_segment_2_0.DEC2[3].n0 top_segment_2_0.DEC2[3].t0 87.8063
R6122 top_segment_2_0.DEC2[3].n21 top_segment_2_0.DEC2[3].t5 81.5883
R6123 top_segment_2_0.DEC2[3].n20 top_segment_2_0.DEC2[3].n4 47.4151
R6124 top_segment_2_0.DEC2[3] top_segment_2_0.DEC2[3].n20 21.8672
R6125 top_segment_2_0.DEC2[3].n23 top_segment_2_0.DEC2[3] 13.9702
R6126 top_segment_2_0.DEC2[3].n20 top_segment_2_0.DEC2[3] 12.6356
R6127 top_segment_2_0.DEC2[3] top_segment_2_0.DEC2[3].n22 11.4706
R6128 top_segment_2_0.DEC2[3].n3 top_segment_2_0.DEC2[3].n2 5.73592
R6129 top_segment_2_0.DEC2[3] top_segment_2_0.DEC2[3].n3 5.66196
R6130 top_segment_2_0.DEC2[3].n4 top_segment_2_0.DEC2[3] 4.85387
R6131 top_segment_2_0.DEC2[3].n17 top_segment_2_0.DEC2[3].n16 4.5005
R6132 top_segment_2_0.DEC2[3].n19 top_segment_2_0.DEC2[3].n18 4.5005
R6133 top_segment_2_0.DEC2[3].n22 top_segment_2_0.DEC2[3] 4.48881
R6134 top_segment_2_0.DEC2[3].n18 top_segment_2_0.DEC2[3].n17 2.588
R6135 top_segment_2_0.DEC2[3] top_segment_2_0.DEC2[3].n23 1.02238
R6136 top_segment_2_0.DEC2[3].n23 top_segment_2_0.DEC2[3] 0.7755
R6137 top_segment_2_0.DEC2[3].n2 top_segment_2_0.DEC2[3].n1 0.713
R6138 top_segment_2_0.DEC2[3].n16 top_segment_2_0.DEC2[3].n15 0.663962
R6139 top_segment_2_0.DEC2[3].n15 top_segment_2_0.DEC2[3].n14 0.663962
R6140 top_segment_2_0.DEC2[3].n14 top_segment_2_0.DEC2[3].n13 0.663962
R6141 top_segment_2_0.DEC2[3].n13 top_segment_2_0.DEC2[3].n12 0.663962
R6142 top_segment_2_0.DEC2[3].n12 top_segment_2_0.DEC2[3].n11 0.663962
R6143 top_segment_2_0.DEC2[3].n6 top_segment_2_0.DEC2[3].n5 0.663962
R6144 top_segment_2_0.DEC2[3].n7 top_segment_2_0.DEC2[3].n6 0.663962
R6145 top_segment_2_0.DEC2[3].n8 top_segment_2_0.DEC2[3].n7 0.663962
R6146 top_segment_2_0.DEC2[3].n9 top_segment_2_0.DEC2[3].n8 0.663962
R6147 top_segment_2_0.DEC2[3].n10 top_segment_2_0.DEC2[3].n9 0.663962
R6148 top_segment_2_0.DEC2[3].n19 top_segment_2_0.DEC2[3].n10 0.663962
R6149 top_segment_2_0.DEC2[3] top_segment_2_0.DEC2[3].n19 0.311626
R6150 top_segment_2_0.DEC2[3].n3 top_segment_2_0.DEC2[3].n0 0.197295
R6151 a_28327_6674.n2 a_28327_6674.t3 245.879
R6152 a_28327_6674.n0 a_28327_6674.t1 241.619
R6153 a_28327_6674.n0 a_28327_6674.t4 240.234
R6154 a_28327_6674.n1 a_28327_6674.t2 238.593
R6155 a_28327_6674.t0 a_28327_6674.n2 238.593
R6156 a_28327_6674.n2 a_28327_6674.n1 6.788
R6157 a_28327_6674.n1 a_28327_6674.n0 4.94008
R6158 top_segment_1_0.rseg_1_v3_1.v56 top_segment_1_0.rseg_1_v3_1.v56.t1 249.738
R6159 top_segment_1_0.rseg_1_v3_1.v56.n0 top_segment_1_0.rseg_1_v3_1.v56.t2 13.4579
R6160 top_segment_1_0.rseg_1_v3_1.v56.n0 top_segment_1_0.rseg_1_v3_1.v56.t0 10.7857
R6161 top_segment_1_0.rseg_1_v3_1.v56 top_segment_1_0.rseg_1_v3_1.v56.n0 4.72836
R6162 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n6 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t9 142.488
R6163 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n5 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t10 142.488
R6164 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t12 142.488
R6165 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t6 142.488
R6166 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n6 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t13 141.704
R6167 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n5 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t11 141.704
R6168 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t8 141.704
R6169 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t7 141.704
R6170 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n8 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t2 139.454
R6171 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t0 139.454
R6172 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n12 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t4 135.305
R6173 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n10 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t1 135.246
R6174 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t3 135.246
R6175 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t5 135.244
R6176 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n12 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n11 12.38
R6177 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n11 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n0 5.038
R6178 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n11 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n10 4.5005
R6179 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n8 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n7 2.2505
R6180 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n3 2.2505
R6181 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n9 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n4 0.842167
R6182 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n9 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n8 0.842167
R6183 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n7 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n5 0.783833
R6184 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n7 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n6 0.783833
R6185 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n1 0.783833
R6186 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n2 0.783833
R6187 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n9 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n0 0.26925
R6188 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n10 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n9 0.26925
R6189 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n12 0.063
R6190 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t0 157.346
R6191 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t2 142.179
R6192 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t3 140.314
R6193 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t1 140.065
R6194 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n0 7.42011
R6195 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n2 0.063
R6196 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n1 0.0171667
R6197 a_26167_5238.n2 a_26167_5238.t3 247.553
R6198 a_26167_5238.n0 a_26167_5238.t4 245.569
R6199 a_26167_5238.n1 a_26167_5238.t2 244.964
R6200 a_26167_5238.n0 a_26167_5238.t1 238.899
R6201 a_26167_5238.t0 a_26167_5238.n2 238.899
R6202 a_26167_5238.n1 a_26167_5238.n0 5.463
R6203 a_26167_5238.n2 a_26167_5238.n1 1.55883
R6204 a_32181_7938.n0 a_32181_7938.t2 244.725
R6205 a_32181_7938.n0 a_32181_7938.t1 242.994
R6206 a_32181_7938.t0 a_32181_7938.n0 239.673
R6207 top_segment_1_0.rseg_1_v3_1.v39 top_segment_1_0.rseg_1_v3_1.v39.t2 248.075
R6208 top_segment_1_0.rseg_1_v3_1.v39.n0 top_segment_1_0.rseg_1_v3_1.v39.t0 10.575
R6209 top_segment_1_0.rseg_1_v3_1.v39.n0 top_segment_1_0.rseg_1_v3_1.v39.t1 10.5739
R6210 top_segment_1_0.rseg_1_v3_1.v39 top_segment_1_0.rseg_1_v3_1.v39.n0 4.2135
R6211 top_segment_1_0.rseg_1_v3_1.v38 top_segment_1_0.rseg_1_v3_1.v38.t2 246.885
R6212 top_segment_1_0.rseg_1_v3_1.v38.n0 top_segment_1_0.rseg_1_v3_1.v38.t0 10.5306
R6213 top_segment_1_0.rseg_1_v3_1.v38.n0 top_segment_1_0.rseg_1_v3_1.v38.t1 10.5285
R6214 top_segment_1_0.rseg_1_v3_1.v38 top_segment_1_0.rseg_1_v3_1.v38.n0 3.53633
R6215 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t12 739.633
R6216 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t11 229.369
R6217 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t7 229.369
R6218 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t6 212.081
R6219 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t5 212.081
R6220 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 203.923
R6221 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 186.001
R6222 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t4 157.07
R6223 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t8 157.07
R6224 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 152.712
R6225 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 152.475
R6226 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t10 139.78
R6227 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t9 139.78
R6228 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 101.49
R6229 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 61.346
R6230 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t2 26.5955
R6231 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t3 26.5955
R6232 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t0 24.9236
R6233 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t1 24.9236
R6234 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 15.8609
R6235 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[0] 13.7651
R6236 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 13.5685
R6237 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 10.7525
R6238 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 10.2234
R6239 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 9.77342
R6240 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 9.64425
R6241 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 9.30224
R6242 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y 6.6565
R6243 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.B 5.45235
R6244 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.B 5.21532
R6245 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y 5.04292
R6246 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 4.91925
R6247 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y 3.8405
R6248 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.A 3.0725
R6249 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y 2.5605
R6250 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 1.93989
R6251 a_43570_17828.t0 a_43570_17828.t1 49.8467
R6252 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t19 241.536
R6253 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t11 241.536
R6254 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t14 230.155
R6255 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t6 230.155
R6256 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t5 229.369
R6257 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t4 228.649
R6258 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t8 212.081
R6259 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t18 212.081
R6260 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n21 203.922
R6261 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n3 186.001
R6262 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t12 169.237
R6263 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t7 169.237
R6264 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n5 157.927
R6265 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t17 157.856
R6266 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t15 157.856
R6267 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t9 157.07
R6268 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t16 156.35
R6269 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n11 154.934
R6270 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n13 154.744
R6271 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n15 154.744
R6272 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n8 153.338
R6273 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n6 152
R6274 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t13 139.78
R6275 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t10 139.78
R6276 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n0 101.49
R6277 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n2 61.346
R6278 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t3 26.5955
R6279 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t0 26.5955
R6280 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t1 24.9236
R6281 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t2 24.9236
R6282 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 24.013
R6283 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 21.1432
R6284 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 19.8144
R6285 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n7 19.6746
R6286 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n16 18.2347
R6287 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n9 18.2231
R6288 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 17.3957
R6289 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 13.5685
R6290 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n17 12.788
R6291 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 10.7525
R6292 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n18 9.64425
R6293 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n4 9.30224
R6294 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 6.6565
R6295 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n20 5.04292
R6296 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n19 3.8405
R6297 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 3.0725
R6298 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 3.05722
R6299 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n1 2.5605
R6300 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n14 2.37941
R6301 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 2.13383
R6302 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 1.93989
R6303 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n12 1.08448
R6304 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n10 1.05323
R6305 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.186047
R6306 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n1 267.599
R6307 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t6 229.369
R6308 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n0 202.094
R6309 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t5 157.07
R6310 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n3 152
R6311 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t4 132.982
R6312 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n5 61.3652
R6313 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t3 32.5055
R6314 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t2 32.5055
R6315 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t1 26.5955
R6316 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.t0 26.5955
R6317 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n4 19.8407
R6318 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 5.92643
R6319 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n6 4.04261
R6320 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B.n2 1.12991
R6321 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[3] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t5 748.038
R6322 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 237.577
R6323 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t4 230.576
R6324 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t3 158.275
R6325 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 152.8
R6326 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t1 139.514
R6327 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t0 26.5955
R6328 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t2 26.5955
R6329 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y 16.1887
R6330 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 10.0771
R6331 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 9.63258
R6332 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 9.41227
R6333 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y 6.98232
R6334 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_0.A 5.86717
R6335 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[3] 5.74157
R6336 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y 2.23542
R6337 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[3] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[3] 0.830857
R6338 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 0.508436
R6339 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 0.291409
R6340 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[3] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t2 756.356
R6341 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t0 235.56
R6342 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_0.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t1 152.889
R6343 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[3] 14.6392
R6344 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_0.Y 2.22659
R6345 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_0.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 1.55202
R6346 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[3] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[3] 0.826393
R6347 top_segment_3_0.bb[6].n2 top_segment_3_0.bb[6].n1 863.124
R6348 top_segment_3_0.bb[6].n1 top_segment_3_0.bb[6].n0 585
R6349 top_segment_3_0.bb[6] top_segment_3_0.bb[6].t0 495.469
R6350 top_segment_3_0.bb[6].n4 top_segment_3_0.bb[6].t6 217.555
R6351 top_segment_3_0.bb[6].n11 top_segment_3_0.bb[6].t9 216.893
R6352 top_segment_3_0.bb[6].n4 top_segment_3_0.bb[6].t11 216.893
R6353 top_segment_3_0.bb[6].n5 top_segment_3_0.bb[6].t5 216.893
R6354 top_segment_3_0.bb[6].n6 top_segment_3_0.bb[6].t10 216.893
R6355 top_segment_3_0.bb[6].n7 top_segment_3_0.bb[6].t12 216.893
R6356 top_segment_3_0.bb[6].n8 top_segment_3_0.bb[6].t8 216.893
R6357 top_segment_3_0.bb[6].n9 top_segment_3_0.bb[6].t2 216.893
R6358 top_segment_3_0.bb[6].n10 top_segment_3_0.bb[6].t4 216.893
R6359 top_segment_3_0.bb[6].n14 top_segment_3_0.bb[6].n13 152
R6360 top_segment_3_0.bb[6].n3 top_segment_3_0.bb[6].t1 141.189
R6361 top_segment_3_0.bb[6].n1 top_segment_3_0.bb[6].t0 140.738
R6362 top_segment_3_0.bb[6].n13 top_segment_3_0.bb[6].t3 114.031
R6363 top_segment_3_0.bb[6].n13 top_segment_3_0.bb[6].t7 81.5883
R6364 top_segment_3_0.bb[6] top_segment_3_0.bb[6].n12 73.9371
R6365 top_segment_3_0.bb[6].n14 top_segment_3_0.bb[6] 16.7132
R6366 top_segment_3_0.bb[6].n15 top_segment_3_0.bb[6] 13.7979
R6367 top_segment_3_0.bb[6].n15 top_segment_3_0.bb[6] 13.1884
R6368 top_segment_3_0.bb[6].n2 top_segment_3_0.bb[6] 11.6369
R6369 top_segment_3_0.bb[6].n0 top_segment_3_0.bb[6] 10.1408
R6370 top_segment_3_0.bb[6] top_segment_3_0.bb[6].n3 7.94225
R6371 top_segment_3_0.bb[6].n3 top_segment_3_0.bb[6] 6.14988
R6372 top_segment_3_0.bb[6].n15 top_segment_3_0.bb[6] 2.16154
R6373 top_segment_3_0.bb[6].n0 top_segment_3_0.bb[6] 2.16154
R6374 top_segment_3_0.bb[6] top_segment_3_0.bb[6].n14 1.16414
R6375 top_segment_3_0.bb[6] top_segment_3_0.bb[6].n2 0.665435
R6376 top_segment_3_0.bb[6].n10 top_segment_3_0.bb[6].n9 0.663962
R6377 top_segment_3_0.bb[6].n9 top_segment_3_0.bb[6].n8 0.663962
R6378 top_segment_3_0.bb[6].n8 top_segment_3_0.bb[6].n7 0.663962
R6379 top_segment_3_0.bb[6].n7 top_segment_3_0.bb[6].n6 0.663962
R6380 top_segment_3_0.bb[6].n6 top_segment_3_0.bb[6].n5 0.663962
R6381 top_segment_3_0.bb[6].n5 top_segment_3_0.bb[6].n4 0.663962
R6382 top_segment_3_0.bb[6].n11 top_segment_3_0.bb[6].n10 0.658467
R6383 top_segment_3_0.bb[6] top_segment_3_0.bb[6].n15 0.582318
R6384 top_segment_3_0.bb[6].n12 top_segment_3_0.bb[6] 0.155033
R6385 top_segment_3_0.bb[6].n12 top_segment_3_0.bb[6].n11 0.0138929
R6386 top_segment_3_0.rseg_3_v3_0.v2.t0 top_segment_3_0.rseg_3_v3_0.v2.n0 675.611
R6387 top_segment_3_0.rseg_3_v3_0.v2.n0 top_segment_3_0.rseg_3_v3_0.v2.t2 10.8307
R6388 top_segment_3_0.rseg_3_v3_0.v2.n0 top_segment_3_0.rseg_3_v3_0.v2.t1 10.5739
R6389 a_15143_17684.n0 a_15143_17684.t1 671.159
R6390 a_15143_17684.n0 a_15143_17684.t2 666.597
R6391 a_15143_17684.t0 a_15143_17684.n0 665.672
R6392 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t2 672.309
R6393 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t1 10.8249
R6394 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.t0 10.5739
R6395 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51.n0 1.38332
R6396 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t2 673.491
R6397 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t0 10.7482
R6398 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.t1 10.6526
R6399 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50.n0 0.679794
R6400 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t9 241.536
R6401 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t4 241.536
R6402 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t16 230.363
R6403 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t17 230.155
R6404 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t6 230.155
R6405 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t10 229.369
R6406 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t8 229.369
R6407 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n0 203.923
R6408 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n7 181.496
R6409 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t5 169.237
R6410 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t15 169.237
R6411 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n5 159.37
R6412 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t12 158.064
R6413 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n17 157.927
R6414 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t14 157.856
R6415 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t13 157.856
R6416 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t7 157.07
R6417 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t11 157.07
R6418 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n11 156.655
R6419 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n2 153.529
R6420 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n18 152
R6421 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n14 152
R6422 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n23 101.49
R6423 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n21 44.3335
R6424 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n6 40.9264
R6425 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n12 29.3297
R6426 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t1 26.5955
R6427 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t2 26.5955
R6428 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t3 24.9236
R6429 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t0 24.9236
R6430 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n15 18.1923
R6431 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n20 16.335
R6432 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n3 16.0286
R6433 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 13.1418
R6434 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n22 13.0565
R6435 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n1 10.7525
R6436 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n8 9.3005
R6437 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n19 7.9365
R6438 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 6.6565
R6439 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n9 6.5302
R6440 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 5.04292
R6441 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 4.3525
R6442 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 3.49141
R6443 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.86617
R6444 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.5605
R6445 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.5605
R6446 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.3045
R6447 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.10199
R6448 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.03686
R6449 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n24 1.93989
R6450 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n10 1.39698
R6451 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n16 1.06105
R6452 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n13 0.988781
R6453 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n4 0.852062
R6454 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.338391
R6455 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 593.165
R6456 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 237.577
R6457 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 140.53
R6458 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 26.5955
R6459 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 26.5955
R6460 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 16.5652
R6461 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 9.03579
R6462 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 1.72748
R6463 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t0 227.856
R6464 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n2 152.333
R6465 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t3 140.382
R6466 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t4 114.031
R6467 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t1 83.3993
R6468 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.t2 81.5883
R6469 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n3 14.4422
R6470 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n1 7.56882
R6471 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n0 5.08175
R6472 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R6473 top_segment_3_0.bb[4].n2 top_segment_3_0.bb[4].n1 863.124
R6474 top_segment_3_0.bb[4].n1 top_segment_3_0.bb[4].n0 585
R6475 top_segment_3_0.bb[4] top_segment_3_0.bb[4].t1 495.469
R6476 top_segment_3_0.bb[4] top_segment_3_0.bb[4].t0 291.983
R6477 top_segment_3_0.bb[4].t0 top_segment_3_0.bb[4].n9 285
R6478 top_segment_3_0.bb[4].n4 top_segment_3_0.bb[4].t4 217.555
R6479 top_segment_3_0.bb[4].n3 top_segment_3_0.bb[4].t2 216.893
R6480 top_segment_3_0.bb[4].n5 top_segment_3_0.bb[4].t6 212.393
R6481 top_segment_3_0.bb[4].n7 top_segment_3_0.bb[4].n6 152
R6482 top_segment_3_0.bb[4].n1 top_segment_3_0.bb[4].t1 140.738
R6483 top_segment_3_0.bb[4].n6 top_segment_3_0.bb[4].t3 114.031
R6484 top_segment_3_0.bb[4].n6 top_segment_3_0.bb[4].t5 81.5883
R6485 top_segment_3_0.bb[4] top_segment_3_0.bb[4].n5 76.1359
R6486 top_segment_3_0.bb[4].n7 top_segment_3_0.bb[4] 16.7132
R6487 top_segment_3_0.bb[4].n8 top_segment_3_0.bb[4] 13.7979
R6488 top_segment_3_0.bb[4] top_segment_3_0.bb[4].n8 13.1884
R6489 top_segment_3_0.bb[4] top_segment_3_0.bb[4].n9 12.4126
R6490 top_segment_3_0.bb[4].n2 top_segment_3_0.bb[4] 11.6369
R6491 top_segment_3_0.bb[4].n0 top_segment_3_0.bb[4] 10.1408
R6492 top_segment_3_0.bb[4].n5 top_segment_3_0.bb[4].n4 4.5005
R6493 top_segment_3_0.bb[4].n0 top_segment_3_0.bb[4] 2.16154
R6494 top_segment_3_0.bb[4].n8 top_segment_3_0.bb[4] 2.16154
R6495 top_segment_3_0.bb[4].n9 top_segment_3_0.bb[4] 1.93989
R6496 top_segment_3_0.bb[4] top_segment_3_0.bb[4].n7 1.16414
R6497 top_segment_3_0.bb[4] top_segment_3_0.bb[4].n2 0.665435
R6498 top_segment_3_0.bb[4].n4 top_segment_3_0.bb[4].n3 0.663962
R6499 top_segment_3_0.bb[4].n8 top_segment_3_0.bb[4] 0.582318
R6500 top_segment_3_0.bb[4].n3 top_segment_3_0.bb[4] 0.272135
R6501 top_segment_4_1.bb2.n2 top_segment_4_1.bb2.n1 863.124
R6502 top_segment_4_1.bb2.n1 top_segment_4_1.bb2.n0 585
R6503 top_segment_4_1.bb2 top_segment_4_1.bb2.t1 495.469
R6504 top_segment_4_1.bb2 top_segment_4_1.bb2.t0 291.983
R6505 top_segment_4_1.bb2.t0 top_segment_4_1.bb2.n14 285
R6506 top_segment_4_1.bb2.n3 top_segment_4_1.bb2.t4 217.555
R6507 top_segment_4_1.bb2.n4 top_segment_4_1.bb2.t3 216.893
R6508 top_segment_4_1.bb2.n3 top_segment_4_1.bb2.t5 216.893
R6509 top_segment_4_1.bb2.n8 top_segment_4_1.bb2.t2 213.218
R6510 top_segment_4_1.bb2.n7 top_segment_4_1.bb2.t9 213.218
R6511 top_segment_4_1.bb2.n7 top_segment_4_1.bb2.t11 212.554
R6512 top_segment_4_1.bb2.n6 top_segment_4_1.bb2.t8 212.393
R6513 top_segment_4_1.bb2.n9 top_segment_4_1.bb2.t7 208.054
R6514 top_segment_4_1.bb2.n12 top_segment_4_1.bb2.n11 152
R6515 top_segment_4_1.bb2.n1 top_segment_4_1.bb2.t1 140.738
R6516 top_segment_4_1.bb2.n11 top_segment_4_1.bb2.t10 114.031
R6517 top_segment_4_1.bb2.n11 top_segment_4_1.bb2.t6 81.5883
R6518 top_segment_4_1.bb2.n10 top_segment_4_1.bb2.n6 40.4505
R6519 top_segment_4_1.bb2 top_segment_4_1.bb2.n10 22.0693
R6520 top_segment_4_1.bb2.n12 top_segment_4_1.bb2 16.7132
R6521 top_segment_4_1.bb2.n13 top_segment_4_1.bb2 13.7979
R6522 top_segment_4_1.bb2 top_segment_4_1.bb2.n13 13.1884
R6523 top_segment_4_1.bb2 top_segment_4_1.bb2.n14 12.4126
R6524 top_segment_4_1.bb2.n2 top_segment_4_1.bb2 11.6369
R6525 top_segment_4_1.bb2.n10 top_segment_4_1.bb2.n9 11.3942
R6526 top_segment_4_1.bb2.n0 top_segment_4_1.bb2 10.1408
R6527 top_segment_4_1.bb2.n6 top_segment_4_1.bb2.n5 4.5005
R6528 top_segment_4_1.bb2.n9 top_segment_4_1.bb2.n8 4.5005
R6529 top_segment_4_1.bb2.n0 top_segment_4_1.bb2 2.16154
R6530 top_segment_4_1.bb2.n13 top_segment_4_1.bb2 2.16154
R6531 top_segment_4_1.bb2.n14 top_segment_4_1.bb2 1.93989
R6532 top_segment_4_1.bb2 top_segment_4_1.bb2.n12 1.16414
R6533 top_segment_4_1.bb2 top_segment_4_1.bb2.n2 0.665435
R6534 top_segment_4_1.bb2.n5 top_segment_4_1.bb2.n3 0.663962
R6535 top_segment_4_1.bb2.n5 top_segment_4_1.bb2.n4 0.663962
R6536 top_segment_4_1.bb2.n13 top_segment_4_1.bb2 0.582318
R6537 top_segment_4_1.bb2 top_segment_4_1.bb2.n7 0.445212
R6538 top_segment_4_1.bb2.n4 top_segment_4_1.bb2 0.28175
R6539 top_segment_4_1.bb2.n8 top_segment_4_1.bb2 0.21925
R6540 a_31905_7938.n0 a_31905_7938.t2 244.542
R6541 a_31905_7938.t0 a_31905_7938.n0 242.81
R6542 a_31905_7938.n0 a_31905_7938.t1 239.857
R6543 a_34580_9019.n0 a_34580_9019.t1 241.075
R6544 a_34580_9019.t0 a_34580_9019.n0 239.35
R6545 a_34580_9019.n0 a_34580_9019.t2 238.716
R6546 top_segment_1_0.rseg_1_v3_1.v47.n0 top_segment_1_0.rseg_1_v3_1.v47.t1 240.469
R6547 top_segment_1_0.rseg_1_v3_1.v47.t0 top_segment_1_0.rseg_1_v3_1.v47.n0 10.6713
R6548 top_segment_1_0.rseg_1_v3_1.v47.n0 top_segment_1_0.rseg_1_v3_1.v47.t2 10.5739
R6549 top_segment_1_0.rseg_1_v3_1.v46 top_segment_1_0.rseg_1_v3_1.v46.t2 249.239
R6550 top_segment_1_0.rseg_1_v3_1.v46.n0 top_segment_1_0.rseg_1_v3_1.v46.t1 10.6247
R6551 top_segment_1_0.rseg_1_v3_1.v46.n0 top_segment_1_0.rseg_1_v3_1.v46.t0 10.5295
R6552 top_segment_1_0.rseg_1_v3_1.v46 top_segment_1_0.rseg_1_v3_1.v46.n0 0.872789
R6553 top_segment_4_1.DEC2.n2 top_segment_4_1.DEC2.n1 863.124
R6554 top_segment_4_1.DEC2.n1 top_segment_4_1.DEC2.n0 585
R6555 top_segment_4_1.DEC2 top_segment_4_1.DEC2.t1 495.469
R6556 top_segment_4_1.DEC2.t0 top_segment_4_1.DEC2 291.983
R6557 top_segment_4_1.DEC2.n19 top_segment_4_1.DEC2.t0 285
R6558 top_segment_4_1.DEC2.n9 top_segment_4_1.DEC2.t8 217.555
R6559 top_segment_4_1.DEC2.n14 top_segment_4_1.DEC2.t17 217.555
R6560 top_segment_4_1.DEC2.n3 top_segment_4_1.DEC2.t10 217.555
R6561 top_segment_4_1.DEC2.n9 top_segment_4_1.DEC2.t12 216.893
R6562 top_segment_4_1.DEC2.n10 top_segment_4_1.DEC2.t11 216.893
R6563 top_segment_4_1.DEC2.n11 top_segment_4_1.DEC2.t9 216.893
R6564 top_segment_4_1.DEC2.n12 top_segment_4_1.DEC2.t2 216.893
R6565 top_segment_4_1.DEC2.n13 top_segment_4_1.DEC2.t3 216.893
R6566 top_segment_4_1.DEC2.n8 top_segment_4_1.DEC2.t13 216.893
R6567 top_segment_4_1.DEC2.n7 top_segment_4_1.DEC2.t5 216.893
R6568 top_segment_4_1.DEC2.n6 top_segment_4_1.DEC2.t16 216.893
R6569 top_segment_4_1.DEC2.n5 top_segment_4_1.DEC2.t14 216.893
R6570 top_segment_4_1.DEC2.n4 top_segment_4_1.DEC2.t6 216.893
R6571 top_segment_4_1.DEC2.n3 top_segment_4_1.DEC2.t4 216.893
R6572 top_segment_4_1.DEC2.n16 top_segment_4_1.DEC2.t15 212.393
R6573 top_segment_4_1.DEC2.n15 top_segment_4_1.DEC2.t7 212.393
R6574 top_segment_4_1.DEC2.n1 top_segment_4_1.DEC2.t1 140.738
R6575 top_segment_4_1.DEC2 top_segment_4_1.DEC2.n17 71.8985
R6576 top_segment_4_1.DEC2.n18 top_segment_4_1.DEC2 14.7588
R6577 top_segment_4_1.DEC2.n19 top_segment_4_1.DEC2 12.4126
R6578 top_segment_4_1.DEC2.n2 top_segment_4_1.DEC2 11.6369
R6579 top_segment_4_1.DEC2.n0 top_segment_4_1.DEC2 10.1408
R6580 top_segment_4_1.DEC2.n18 top_segment_4_1.DEC2 7.75808
R6581 top_segment_4_1.DEC2 top_segment_4_1.DEC2.n18 6.59444
R6582 top_segment_4_1.DEC2.n15 top_segment_4_1.DEC2.n14 4.5005
R6583 top_segment_4_1.DEC2.n17 top_segment_4_1.DEC2.n16 4.5005
R6584 top_segment_4_1.DEC2.n0 top_segment_4_1.DEC2 2.16154
R6585 top_segment_4_1.DEC2 top_segment_4_1.DEC2.n19 1.93989
R6586 top_segment_4_1.DEC2 top_segment_4_1.DEC2.n15 1.89425
R6587 top_segment_4_1.DEC2 top_segment_4_1.DEC2.n2 0.665435
R6588 top_segment_4_1.DEC2.n14 top_segment_4_1.DEC2.n13 0.663962
R6589 top_segment_4_1.DEC2.n13 top_segment_4_1.DEC2.n12 0.663962
R6590 top_segment_4_1.DEC2.n12 top_segment_4_1.DEC2.n11 0.663962
R6591 top_segment_4_1.DEC2.n11 top_segment_4_1.DEC2.n10 0.663962
R6592 top_segment_4_1.DEC2.n10 top_segment_4_1.DEC2.n9 0.663962
R6593 top_segment_4_1.DEC2.n4 top_segment_4_1.DEC2.n3 0.663962
R6594 top_segment_4_1.DEC2.n5 top_segment_4_1.DEC2.n4 0.663962
R6595 top_segment_4_1.DEC2.n6 top_segment_4_1.DEC2.n5 0.663962
R6596 top_segment_4_1.DEC2.n7 top_segment_4_1.DEC2.n6 0.663962
R6597 top_segment_4_1.DEC2.n8 top_segment_4_1.DEC2.n7 0.663962
R6598 top_segment_4_1.DEC2.n17 top_segment_4_1.DEC2.n8 0.663962
R6599 top_segment_4_1.DEC2.n16 top_segment_4_1.DEC2 0.65675
R6600 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t0 672.795
R6601 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t1 10.7151
R6602 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.t2 10.6674
R6603 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36.n0 2.05222
R6604 a_13588_5238.n0 a_13588_5238.t3 672.827
R6605 a_13588_5238.n1 a_13588_5238.t1 672.455
R6606 a_13588_5238.t0 a_13588_5238.n2 671.236
R6607 a_13588_5238.n1 a_13588_5238.t4 666.034
R6608 a_13588_5238.n0 a_13588_5238.t2 666.034
R6609 a_13588_5238.n2 a_13588_5238.n1 5.78175
R6610 a_13588_5238.n2 a_13588_5238.n0 0.779667
R6611 top_segment_4_1.b2.n2 top_segment_4_1.b2.n1 863.124
R6612 top_segment_4_1.b2.n1 top_segment_4_1.b2.n0 585
R6613 top_segment_4_1.b2 top_segment_4_1.b2.t1 495.469
R6614 top_segment_4_1.b2.t0 top_segment_4_1.b2 291.983
R6615 top_segment_4_1.b2.n12 top_segment_4_1.b2.t0 285
R6616 top_segment_4_1.b2.n5 top_segment_4_1.b2.t4 217.555
R6617 top_segment_4_1.b2.n4 top_segment_4_1.b2.t9 216.893
R6618 top_segment_4_1.b2.n3 top_segment_4_1.b2.t8 216.893
R6619 top_segment_4_1.b2.n8 top_segment_4_1.b2.t2 213.218
R6620 top_segment_4_1.b2.n7 top_segment_4_1.b2.t3 213.218
R6621 top_segment_4_1.b2.n7 top_segment_4_1.b2.t5 212.554
R6622 top_segment_4_1.b2.n6 top_segment_4_1.b2.t7 212.393
R6623 top_segment_4_1.b2.n9 top_segment_4_1.b2.t6 208.054
R6624 top_segment_4_1.b2.n1 top_segment_4_1.b2.t1 140.738
R6625 top_segment_4_1.b2.n10 top_segment_4_1.b2.n6 45.4047
R6626 top_segment_4_1.b2 top_segment_4_1.b2.n10 19.6734
R6627 top_segment_4_1.b2.n11 top_segment_4_1.b2 14.3755
R6628 top_segment_4_1.b2.n12 top_segment_4_1.b2 12.4126
R6629 top_segment_4_1.b2.n2 top_segment_4_1.b2 11.6369
R6630 top_segment_4_1.b2.n10 top_segment_4_1.b2.n9 11.5776
R6631 top_segment_4_1.b2.n0 top_segment_4_1.b2 10.1408
R6632 top_segment_4_1.b2.n11 top_segment_4_1.b2 8.53383
R6633 top_segment_4_1.b2 top_segment_4_1.b2.n11 5.81868
R6634 top_segment_4_1.b2.n6 top_segment_4_1.b2.n5 4.5005
R6635 top_segment_4_1.b2.n9 top_segment_4_1.b2.n8 4.5005
R6636 top_segment_4_1.b2.n0 top_segment_4_1.b2 2.16154
R6637 top_segment_4_1.b2 top_segment_4_1.b2.n12 1.93989
R6638 top_segment_4_1.b2 top_segment_4_1.b2.n2 0.665435
R6639 top_segment_4_1.b2.n4 top_segment_4_1.b2.n3 0.663962
R6640 top_segment_4_1.b2.n5 top_segment_4_1.b2.n4 0.663962
R6641 top_segment_4_1.b2.n8 top_segment_4_1.b2 0.380308
R6642 top_segment_4_1.b2 top_segment_4_1.b2.n7 0.284154
R6643 top_segment_4_1.b2.n3 top_segment_4_1.b2 0.180788
R6644 a_32851_7938.n0 a_32851_7938.t2 245.95
R6645 a_32851_7938.t0 a_32851_7938.n0 243.918
R6646 a_32851_7938.n0 a_32851_7938.t1 239.124
R6647 VL2.n0 VL2.t2 240.29
R6648 VL2.n2 VL2.t3 239.082
R6649 VL2.n1 VL2.t1 239.082
R6650 VL2.n0 VL2.t0 239.082
R6651 VL2.n1 VL2.n0 1.20883
R6652 VL2 VL2.n1 0.94425
R6653 VL2 VL2.n2 0.265083
R6654 VL2.n2 VL2 0.063
R6655 a_21596_17121.n0 a_21596_17121.t3 242.181
R6656 a_21596_17121.n3 a_21596_17121.t5 240.082
R6657 a_21596_17121.t0 a_21596_17121.n3 239.415
R6658 a_21596_17121.n2 a_21596_17121.t2 239.248
R6659 a_21596_17121.n1 a_21596_17121.t1 239.248
R6660 a_21596_17121.n0 a_21596_17121.t4 239.248
R6661 a_21596_17121.n3 a_21596_17121.n2 3.40883
R6662 a_21596_17121.n1 a_21596_17121.n0 2.93383
R6663 a_21596_17121.n2 a_21596_17121.n1 2.93383
R6664 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t4 232.293
R6665 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t5 222.117
R6666 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t15 139.66
R6667 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t0 139.454
R6668 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t2 139.454
R6669 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n25 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t12 139.206
R6670 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t9 139.206
R6671 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t6 139.206
R6672 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t26 139.206
R6673 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t21 139.206
R6674 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t18 139.206
R6675 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t14 139.206
R6676 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t13 139.206
R6677 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t10 139.206
R6678 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t7 139.206
R6679 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t27 139.206
R6680 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t23 139.206
R6681 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t20 139.206
R6682 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t22 139.206
R6683 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t19 139.206
R6684 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t16 139.206
R6685 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t8 139.206
R6686 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t11 139.206
R6687 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t25 139.206
R6688 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t28 139.206
R6689 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t17 139.206
R6690 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t1 135.197
R6691 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t3 134.625
R6692 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t24 17.157
R6693 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n27 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n26 13.2737
R6694 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n27 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n4 6.81925
R6695 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n2 4.5005
R6696 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n27 4.44425
R6697 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n3 1.10467
R6698 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R6699 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n23 0.804667
R6700 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R6701 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n21 0.804667
R6702 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R6703 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n19 0.804667
R6704 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R6705 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n17 0.804667
R6706 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R6707 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n15 0.804667
R6708 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R6709 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n13 0.804667
R6710 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R6711 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n11 0.804667
R6712 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R6713 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n9 0.804667
R6714 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R6715 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n7 0.804667
R6716 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.804667
R6717 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n5 0.804667
R6718 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n0 0.701587
R6719 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n26 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n25 0.660917
R6720 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n1 0.51454
R6721 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n25 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n24 0.454667
R6722 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n22 0.454667
R6723 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n20 0.454667
R6724 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n18 0.454667
R6725 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n16 0.454667
R6726 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n14 0.454667
R6727 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n12 0.454667
R6728 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n10 0.454667
R6729 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n8 0.454667
R6730 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n6 0.454667
R6731 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n26 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.01925
R6732 a_42271_15290.t0 a_42271_15290.t1 55.3905
R6733 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t3 221.851
R6734 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t1 221.851
R6735 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t5 140.625
R6736 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t4 140.244
R6737 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t7 113.648
R6738 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t6 113.648
R6739 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t0 108.365
R6740 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.t2 108.365
R6741 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.D1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n5 12.9957
R6742 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n5 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n4 1.44557
R6743 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n3 0.557293
R6744 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n1 0.557293
R6745 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n5 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n2 0.266714
R6746 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.D1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D1.n0 0.063
R6747 a_35435_18538.n1 a_35435_18538.t0 239.831
R6748 a_35435_18538.t1 a_35435_18538.n1 226.853
R6749 a_35435_18538.n0 a_35435_18538.t3 223.633
R6750 a_35435_18538.n0 a_35435_18538.t2 221.851
R6751 a_35435_18538.n1 a_35435_18538.n0 5.73071
R6752 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t17 739.082
R6753 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t15 241.536
R6754 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t4 230.155
R6755 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t13 230.155
R6756 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t6 230.155
R6757 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t14 230.155
R6758 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t9 230.155
R6759 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t11 230.155
R6760 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n26 203.922
R6761 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 181.496
R6762 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t10 169.237
R6763 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t7 157.856
R6764 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t18 157.856
R6765 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t16 157.856
R6766 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t8 157.856
R6767 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t5 157.856
R6768 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t12 157.856
R6769 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 154.867
R6770 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 153.911
R6771 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 153.338
R6772 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 152
R6773 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 152
R6774 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 152
R6775 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 101.49
R6776 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n26 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t0 26.5955
R6777 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n26 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t3 26.5955
R6778 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 25.9222
R6779 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t1 24.9236
R6780 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t2 24.9236
R6781 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 21.542
R6782 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 21.248
R6783 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 19.5688
R6784 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 19.3054
R6785 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 18.6011
R6786 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 18.542
R6787 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y 13.0565
R6788 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[0] 12.2693
R6789 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 12.2559
R6790 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 11.1817
R6791 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 11.0199
R6792 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y 10.7525
R6793 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y 6.6565
R6794 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 5.10675
R6795 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 5.04292
R6796 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 4.3525
R6797 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x2.A 3.05722
R6798 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x1.B 2.5605
R6799 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 2.5605
R6800 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.A 2.48408
R6801 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.A 2.10199
R6802 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.A 2.10199
R6803 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x2.A 2.10199
R6804 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y 1.93989
R6805 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x3.A 1.52886
R6806 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 1.40284
R6807 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 1.23683
R6808 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 0.926281
R6809 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 0.842297
R6810 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[6] 0.119641
R6811 a_18217_7938.t0 a_18217_7938.n0 671.409
R6812 a_18217_7938.n0 a_18217_7938.t2 670.924
R6813 a_18217_7938.n0 a_18217_7938.t1 665.707
R6814 a_19479_9019.n0 a_19479_9019.t2 667.659
R6815 a_19479_9019.n0 a_19479_9019.t1 665.933
R6816 a_19479_9019.t0 a_19479_9019.n0 665.299
R6817 top_segment_1_0.rseg_1_v3_1.v49.n0 top_segment_1_0.rseg_1_v3_1.v49.t1 236.649
R6818 top_segment_1_0.rseg_1_v3_1.v49.n0 top_segment_1_0.rseg_1_v3_1.v49.t2 10.6713
R6819 top_segment_1_0.rseg_1_v3_1.v49.t0 top_segment_1_0.rseg_1_v3_1.v49.n0 10.5739
R6820 top_segment_1_0.rseg_1_v3_1.v50 top_segment_1_0.rseg_1_v3_1.v50.t1 246.716
R6821 top_segment_1_0.rseg_1_v3_1.v50.n0 top_segment_1_0.rseg_1_v3_1.v50.t0 10.5306
R6822 top_segment_1_0.rseg_1_v3_1.v50.n0 top_segment_1_0.rseg_1_v3_1.v50.t2 10.5285
R6823 top_segment_1_0.rseg_1_v3_1.v50 top_segment_1_0.rseg_1_v3_1.v50.n0 0.886534
R6824 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t0 157.49
R6825 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t2 142.079
R6826 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t1 140.304
R6827 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t3 139.327
R6828 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n0 7.54544
R6829 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n1 0.063
R6830 top_segment_4_1.b3.n2 top_segment_4_1.b3.n1 863.124
R6831 top_segment_4_1.b3.n1 top_segment_4_1.b3.n0 585
R6832 top_segment_4_1.b3 top_segment_4_1.b3.t1 495.469
R6833 top_segment_4_1.b3.t0 top_segment_4_1.b3 291.983
R6834 top_segment_4_1.b3.n23 top_segment_4_1.b3.t0 285
R6835 top_segment_4_1.b3.n11 top_segment_4_1.b3.t15 217.555
R6836 top_segment_4_1.b3.n9 top_segment_4_1.b3.t16 217.555
R6837 top_segment_4_1.b3.n8 top_segment_4_1.b3.t6 216.893
R6838 top_segment_4_1.b3.n7 top_segment_4_1.b3.t4 216.893
R6839 top_segment_4_1.b3.n6 top_segment_4_1.b3.t11 216.893
R6840 top_segment_4_1.b3.n5 top_segment_4_1.b3.t7 216.893
R6841 top_segment_4_1.b3.n4 top_segment_4_1.b3.t18 216.893
R6842 top_segment_4_1.b3.n3 top_segment_4_1.b3.t3 216.893
R6843 top_segment_4_1.b3.n14 top_segment_4_1.b3.t19 213.218
R6844 top_segment_4_1.b3 top_segment_4_1.b3.t14 212.77
R6845 top_segment_4_1.b3.n18 top_segment_4_1.b3.t17 212.554
R6846 top_segment_4_1.b3.n17 top_segment_4_1.b3.t8 212.554
R6847 top_segment_4_1.b3.n16 top_segment_4_1.b3.t5 212.554
R6848 top_segment_4_1.b3.n15 top_segment_4_1.b3.t13 212.554
R6849 top_segment_4_1.b3.n14 top_segment_4_1.b3.t9 212.554
R6850 top_segment_4_1.b3.n12 top_segment_4_1.b3.t2 212.393
R6851 top_segment_4_1.b3.n10 top_segment_4_1.b3.t10 212.393
R6852 top_segment_4_1.b3.n20 top_segment_4_1.b3.t12 208.054
R6853 top_segment_4_1.b3.n1 top_segment_4_1.b3.t1 140.738
R6854 top_segment_4_1.b3.n21 top_segment_4_1.b3.n13 39.9172
R6855 top_segment_4_1.b3 top_segment_4_1.b3.n21 18.2588
R6856 top_segment_4_1.b3.n13 top_segment_4_1.b3.n10 15.6484
R6857 top_segment_4_1.b3.n13 top_segment_4_1.b3.n12 14.6859
R6858 top_segment_4_1.b3.n22 top_segment_4_1.b3 14.3755
R6859 top_segment_4_1.b3.n21 top_segment_4_1.b3.n20 14.1963
R6860 top_segment_4_1.b3.n23 top_segment_4_1.b3 12.4126
R6861 top_segment_4_1.b3.n2 top_segment_4_1.b3 11.6369
R6862 top_segment_4_1.b3.n0 top_segment_4_1.b3 10.1408
R6863 top_segment_4_1.b3.n22 top_segment_4_1.b3 8.53383
R6864 top_segment_4_1.b3 top_segment_4_1.b3.n22 5.81868
R6865 top_segment_4_1.b3.n12 top_segment_4_1.b3.n11 4.5005
R6866 top_segment_4_1.b3.n10 top_segment_4_1.b3.n9 4.5005
R6867 top_segment_4_1.b3.n20 top_segment_4_1.b3.n19 4.5005
R6868 top_segment_4_1.b3.n0 top_segment_4_1.b3 2.16154
R6869 top_segment_4_1.b3 top_segment_4_1.b3.n23 1.93989
R6870 top_segment_4_1.b3 top_segment_4_1.b3.n2 0.665435
R6871 top_segment_4_1.b3.n4 top_segment_4_1.b3.n3 0.663962
R6872 top_segment_4_1.b3.n5 top_segment_4_1.b3.n4 0.663962
R6873 top_segment_4_1.b3.n6 top_segment_4_1.b3.n5 0.663962
R6874 top_segment_4_1.b3.n7 top_segment_4_1.b3.n6 0.663962
R6875 top_segment_4_1.b3.n8 top_segment_4_1.b3.n7 0.663962
R6876 top_segment_4_1.b3.n9 top_segment_4_1.b3.n8 0.663962
R6877 top_segment_4_1.b3.n15 top_segment_4_1.b3.n14 0.663962
R6878 top_segment_4_1.b3.n16 top_segment_4_1.b3.n15 0.663962
R6879 top_segment_4_1.b3.n17 top_segment_4_1.b3.n16 0.663962
R6880 top_segment_4_1.b3.n19 top_segment_4_1.b3.n17 0.663962
R6881 top_segment_4_1.b3.n19 top_segment_4_1.b3.n18 0.663962
R6882 top_segment_4_1.b3.n18 top_segment_4_1.b3 0.447615
R6883 top_segment_4_1.b3.n11 top_segment_4_1.b3 0.322615
R6884 top_segment_4_1.b3.n3 top_segment_4_1.b3 0.226462
R6885 a_16555_17684.t0 a_16555_17684.n1 667.399
R6886 a_16555_17684.n0 a_16555_17684.t2 666.116
R6887 a_16555_17684.n1 a_16555_17684.t3 665.615
R6888 a_16555_17684.n0 a_16555_17684.t1 665.484
R6889 a_16555_17684.n1 a_16555_17684.n0 1.39217
R6890 VH3 VH3.t0 666.581
R6891 VH3.n0 VH3.t1 665.433
R6892 VH3.n0 VH3 0.063
R6893 VH3 VH3.n0 0.0588333
R6894 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 593.158
R6895 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 231.554
R6896 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 140.53
R6897 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 26.5955
R6898 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 26.5955
R6899 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 16.5652
R6900 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 9.03579
R6901 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 6.02403
R6902 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 1.72748
R6903 a_42609_17081.t0 a_42609_17081.t1 129.28
R6904 a_19922_19162.n0 a_19922_19162.t2 251.903
R6905 a_19922_19162.t0 a_19922_19162.n1 248.659
R6906 a_19922_19162.n0 a_19922_19162.t3 241.815
R6907 a_19922_19162.n1 a_19922_19162.t1 238.732
R6908 a_19922_19162.n1 a_19922_19162.n0 3.24425
R6909 top_segment_2_0.rseg_2_v3_0.v16.n0 top_segment_2_0.rseg_2_v3_0.v16.t3 237.774
R6910 top_segment_2_0.rseg_2_v3_0.v16.n1 top_segment_2_0.rseg_2_v3_0.v16.t1 237.685
R6911 top_segment_2_0.rseg_2_v3_0.v16.n0 top_segment_2_0.rseg_2_v3_0.v16.t2 10.6569
R6912 top_segment_2_0.rseg_2_v3_0.v16.t0 top_segment_2_0.rseg_2_v3_0.v16.n1 10.6569
R6913 top_segment_2_0.rseg_2_v3_0.v16.n1 top_segment_2_0.rseg_2_v3_0.v16.n0 3.39554
R6914 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t5 221.851
R6915 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t3 221.851
R6916 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t0 140.061
R6917 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t1 139.566
R6918 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t17 120.969
R6919 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t10 120.969
R6920 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t13 120.969
R6921 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t15 120.969
R6922 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t14 120.969
R6923 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t6 120.969
R6924 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t16 120.969
R6925 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t8 120.969
R6926 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t7 120.969
R6927 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t12 120.969
R6928 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t9 120.969
R6929 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t11 120.969
R6930 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t4 108.365
R6931 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t2 108.365
R6932 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n0 15.3463
R6933 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n15 13.5257
R6934 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n19 8.1267
R6935 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n16 5.84703
R6936 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n1 4.95104
R6937 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n18 4.79425
R6938 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n20 1.21717
R6939 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n3 0.713
R6940 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n4 0.713
R6941 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n5 0.713
R6942 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n13 0.713
R6943 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n12 0.713
R6944 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n11 0.713
R6945 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n9 0.713
R6946 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n8 0.713
R6947 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n7 0.713
R6948 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n10 0.690083
R6949 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.598417
R6950 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n0 0.557293
R6951 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n17 0.546515
R6952 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.523417
R6953 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n14 0.167167
R6954 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n6 0.140083
R6955 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.140083
R6956 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.140083
R6957 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.08175
R6958 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n21 0.063
R6959 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.0525833
R6960 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n2 0.0143889
R6961 a_35957_18086.t1 a_35957_18086.n1 229.328
R6962 a_35957_18086.n1 a_35957_18086.t0 226.986
R6963 a_35957_18086.n0 a_35957_18086.t3 127.692
R6964 a_35957_18086.n1 a_35957_18086.n0 12.484
R6965 a_35957_18086.n0 a_35957_18086.t2 10.584
R6966 a_33679_7938.n0 a_33679_7938.t2 246.316
R6967 a_33679_7938.n0 a_33679_7938.t1 244.469
R6968 a_33679_7938.t0 a_33679_7938.n0 238.573
R6969 a_33724_9019.n0 a_33724_9019.t1 243.633
R6970 a_33724_9019.t0 a_33724_9019.n0 241.625
R6971 a_33724_9019.n0 a_33724_9019.t2 239.267
R6972 a_29155_6674.n2 a_29155_6674.t3 246.429
R6973 a_29155_6674.n0 a_29155_6674.t4 241.959
R6974 a_29155_6674.n0 a_29155_6674.t1 239.822
R6975 a_29155_6674.n1 a_29155_6674.t2 239.143
R6976 a_29155_6674.t0 a_29155_6674.n2 239.143
R6977 a_29155_6674.n2 a_29155_6674.n1 6.788
R6978 a_29155_6674.n1 a_29155_6674.n0 3.76508
R6979 top_segment_1_0.rseg_1_v3_1.v27 top_segment_1_0.rseg_1_v3_1.v27.t0 248.95
R6980 top_segment_1_0.rseg_1_v3_1.v27.n0 top_segment_1_0.rseg_1_v3_1.v27.t2 10.6701
R6981 top_segment_1_0.rseg_1_v3_1.v27.n0 top_segment_1_0.rseg_1_v3_1.v27.t1 10.5739
R6982 top_segment_1_0.rseg_1_v3_1.v27 top_segment_1_0.rseg_1_v3_1.v27.n0 2.76539
R6983 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t3 274.793
R6984 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t0 268.077
R6985 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t0 263.695
R6986 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t4 232.214
R6987 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n1 205.28
R6988 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t5 159.915
R6989 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n3 152.207
R6990 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n2 54.4975
R6991 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n0 36.5181
R6992 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t2 26.5955
R6993 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.t1 26.5955
R6994 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n4 20.6093
R6995 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n5 12.9887
R6996 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 4.54244
R6997 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t2 675.533
R6998 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t0 10.7601
R6999 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.t1 10.7161
R7000 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27.n0 2.73056
R7001 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t2 676.553
R7002 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t1 10.7798
R7003 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t0 10.6302
R7004 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.n0 3.43637
R7005 a_42245_14694.t0 a_42245_14694.n0 228.04
R7006 a_42245_14694.n0 a_42245_14694.t2 145.648
R7007 a_42245_14694.n0 a_42245_14694.t1 83.2159
R7008 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t1 227.856
R7009 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n2 152.333
R7010 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t3 140.382
R7011 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t4 114.031
R7012 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t0 83.3993
R7013 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.t2 81.5883
R7014 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n3 14.4422
R7015 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n1 7.56882
R7016 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n0 5.08175
R7017 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R7018 a_42271_14854.t0 a_42271_14854.t1 55.3905
R7019 a_19045_7938.t0 a_19045_7938.n0 671.928
R7020 a_19045_7938.n0 a_19045_7938.t2 671.475
R7021 a_19045_7938.n0 a_19045_7938.t1 665.158
R7022 a_18623_9019.t0 a_18623_9019.n0 670.216
R7023 a_18623_9019.n0 a_18623_9019.t2 668.208
R7024 a_18623_9019.n0 a_18623_9019.t1 665.85
R7025 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 593.165
R7026 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 237.577
R7027 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 140.53
R7028 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 26.5955
R7029 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 26.5955
R7030 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 16.5652
R7031 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 9.03579
R7032 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 1.72748
R7033 top_segment_4_1.DEC0.n2 top_segment_4_1.DEC0.n1 863.124
R7034 top_segment_4_1.DEC0.n1 top_segment_4_1.DEC0.n0 585
R7035 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y top_segment_4_1.DEC0.t1 495.469
R7036 top_segment_4_1.DEC0.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 291.983
R7037 top_segment_4_1.DEC0.n20 top_segment_4_1.DEC0.t0 285
R7038 top_segment_4_1.DEC0.n6 top_segment_4_1.DEC0.t17 217.555
R7039 top_segment_4_1.DEC0.n3 top_segment_4_1.DEC0.t5 217.555
R7040 top_segment_4_1.DEC0.n10 top_segment_4_1.DEC0.t6 216.893
R7041 top_segment_4_1.DEC0.n11 top_segment_4_1.DEC0.t12 216.893
R7042 top_segment_4_1.DEC0.n12 top_segment_4_1.DEC0.t10 216.893
R7043 top_segment_4_1.DEC0.n13 top_segment_4_1.DEC0.t7 216.893
R7044 top_segment_4_1.DEC0.n14 top_segment_4_1.DEC0.t13 216.893
R7045 top_segment_4_1.DEC0.n15 top_segment_4_1.DEC0.t3 216.893
R7046 top_segment_4_1.DEC0.n16 top_segment_4_1.DEC0.t2 216.893
R7047 top_segment_4_1.DEC0.n17 top_segment_4_1.DEC0.t4 216.893
R7048 top_segment_4_1.DEC0.n6 top_segment_4_1.DEC0.t16 216.893
R7049 top_segment_4_1.DEC0.n7 top_segment_4_1.DEC0.t8 216.893
R7050 top_segment_4_1.DEC0.n8 top_segment_4_1.DEC0.t14 216.893
R7051 top_segment_4_1.DEC0.n5 top_segment_4_1.DEC0.t11 216.893
R7052 top_segment_4_1.DEC0.n4 top_segment_4_1.DEC0.t9 216.893
R7053 top_segment_4_1.DEC0.n3 top_segment_4_1.DEC0.t15 216.893
R7054 top_segment_4_1.DEC0.n1 top_segment_4_1.DEC0.t1 140.738
R7055 top_segment_4_1.DEC0.n18 top_segment_4_1.DEC0.n17 101.117
R7056 top_segment_4_1.DEC0.n19 top_segment_4_1.DEC0.n18 13.9797
R7057 top_segment_4_1.DEC0.n10 top_segment_4_1.DEC0.n9 12.8332
R7058 top_segment_4_1.DEC0.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 12.4126
R7059 top_segment_4_1.DEC0.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 11.6369
R7060 top_segment_4_1.DEC0.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 10.1408
R7061 top_segment_4_1.DEC0.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 8.14595
R7062 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y top_segment_4_1.DEC0.n19 6.20656
R7063 top_segment_4_1.DEC0.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y 2.16154
R7064 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y top_segment_4_1.DEC0.n20 1.93989
R7065 top_segment_4_1.DEC0.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec2b[0] 0.7755
R7066 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y top_segment_4_1.DEC0.n2 0.665435
R7067 top_segment_4_1.DEC0.n8 top_segment_4_1.DEC0.n7 0.663962
R7068 top_segment_4_1.DEC0.n7 top_segment_4_1.DEC0.n6 0.663962
R7069 top_segment_4_1.DEC0.n4 top_segment_4_1.DEC0.n3 0.663962
R7070 top_segment_4_1.DEC0.n5 top_segment_4_1.DEC0.n4 0.663962
R7071 top_segment_4_1.DEC0.n17 top_segment_4_1.DEC0.n16 0.663962
R7072 top_segment_4_1.DEC0.n16 top_segment_4_1.DEC0.n15 0.663962
R7073 top_segment_4_1.DEC0.n15 top_segment_4_1.DEC0.n14 0.663962
R7074 top_segment_4_1.DEC0.n14 top_segment_4_1.DEC0.n13 0.663962
R7075 top_segment_4_1.DEC0.n13 top_segment_4_1.DEC0.n12 0.663962
R7076 top_segment_4_1.DEC0.n12 top_segment_4_1.DEC0.n11 0.663962
R7077 top_segment_4_1.DEC0.n11 top_segment_4_1.DEC0.n10 0.663962
R7078 top_segment_4_1.DEC0.n9 top_segment_4_1.DEC0.n8 0.320692
R7079 top_segment_4_1.DEC0.n9 top_segment_4_1.DEC0.n5 0.320692
R7080 a_41271_17118.t0 a_41271_17118.t1 65.941
R7081 top_segment_4_1.b1.n2 top_segment_4_1.b1.n1 863.124
R7082 top_segment_4_1.b1.n1 top_segment_4_1.b1.n0 585
R7083 top_segment_4_1.b1 top_segment_4_1.b1.t0 495.469
R7084 top_segment_4_1.b1.n4 top_segment_4_1.b1.t4 217.555
R7085 top_segment_4_1.b1 top_segment_4_1.b1.t2 212.911
R7086 top_segment_4_1.b1.n5 top_segment_4_1.b1.t5 212.393
R7087 top_segment_4_1.b1.n6 top_segment_4_1.b1.t3 208.054
R7088 top_segment_4_1.b1.n3 top_segment_4_1.b1.t1 141.189
R7089 top_segment_4_1.b1.n1 top_segment_4_1.b1.t0 140.738
R7090 top_segment_4_1.b1.n7 top_segment_4_1.b1.n5 41.4463
R7091 top_segment_4_1.b1 top_segment_4_1.b1.n7 26.7318
R7092 top_segment_4_1.b1.n8 top_segment_4_1.b1 14.3755
R7093 top_segment_4_1.b1.n2 top_segment_4_1.b1 11.6369
R7094 top_segment_4_1.b1.n7 top_segment_4_1.b1.n6 11.2109
R7095 top_segment_4_1.b1.n0 top_segment_4_1.b1 10.1408
R7096 top_segment_4_1.b1 top_segment_4_1.b1.n8 8.53383
R7097 top_segment_4_1.b1 top_segment_4_1.b1.n3 7.94225
R7098 top_segment_4_1.b1.n3 top_segment_4_1.b1 6.14988
R7099 top_segment_4_1.b1.n8 top_segment_4_1.b1 5.81868
R7100 top_segment_4_1.b1.n6 top_segment_4_1.b1 4.80819
R7101 top_segment_4_1.b1.n5 top_segment_4_1.b1.n4 4.5005
R7102 top_segment_4_1.b1.n0 top_segment_4_1.b1 2.16154
R7103 top_segment_4_1.b1 top_segment_4_1.b1.n2 0.665435
R7104 top_segment_4_1.b1.n4 top_segment_4_1.b1 0.214442
R7105 a_33420_9019.t0 a_33420_9019.n0 240.13
R7106 a_33420_9019.n0 a_33420_9019.t1 239.512
R7107 a_33420_9019.n0 a_33420_9019.t2 238.921
R7108 a_34000_9019.n0 a_34000_9019.t1 242.075
R7109 a_34000_9019.t0 a_34000_9019.n0 241.441
R7110 a_34000_9019.n0 a_34000_9019.t2 239.083
R7111 top_segment_1_0.rseg_1_v3_1.v10 top_segment_1_0.rseg_1_v3_1.v10.t1 250.332
R7112 top_segment_1_0.rseg_1_v3_1.v10.n0 top_segment_1_0.rseg_1_v3_1.v10.t0 10.5317
R7113 top_segment_1_0.rseg_1_v3_1.v10.n0 top_segment_1_0.rseg_1_v3_1.v10.t2 10.5285
R7114 top_segment_1_0.rseg_1_v3_1.v10 top_segment_1_0.rseg_1_v3_1.v10.n0 3.51046
R7115 top_segment_4_1.DEC1.n2 top_segment_4_1.DEC1.n1 863.124
R7116 top_segment_4_1.DEC1.n1 top_segment_4_1.DEC1.n0 585
R7117 top_segment_4_1.DEC1 top_segment_4_1.DEC1.t1 495.469
R7118 top_segment_4_1.DEC1.t0 top_segment_4_1.DEC1 291.983
R7119 top_segment_4_1.DEC1.n20 top_segment_4_1.DEC1.t0 285
R7120 top_segment_4_1.DEC1.n9 top_segment_4_1.DEC1.t9 217.555
R7121 top_segment_4_1.DEC1.n14 top_segment_4_1.DEC1.t2 217.555
R7122 top_segment_4_1.DEC1.n3 top_segment_4_1.DEC1.t11 217.555
R7123 top_segment_4_1.DEC1.n9 top_segment_4_1.DEC1.t7 216.893
R7124 top_segment_4_1.DEC1.n10 top_segment_4_1.DEC1.t6 216.893
R7125 top_segment_4_1.DEC1.n11 top_segment_4_1.DEC1.t10 216.893
R7126 top_segment_4_1.DEC1.n12 top_segment_4_1.DEC1.t8 216.893
R7127 top_segment_4_1.DEC1.n13 top_segment_4_1.DEC1.t17 216.893
R7128 top_segment_4_1.DEC1.n8 top_segment_4_1.DEC1.t15 216.893
R7129 top_segment_4_1.DEC1.n7 top_segment_4_1.DEC1.t13 216.893
R7130 top_segment_4_1.DEC1.n6 top_segment_4_1.DEC1.t12 216.893
R7131 top_segment_4_1.DEC1.n5 top_segment_4_1.DEC1.t16 216.893
R7132 top_segment_4_1.DEC1.n4 top_segment_4_1.DEC1.t14 216.893
R7133 top_segment_4_1.DEC1.n3 top_segment_4_1.DEC1.t5 216.893
R7134 top_segment_4_1.DEC1.n16 top_segment_4_1.DEC1.t3 212.393
R7135 top_segment_4_1.DEC1.n15 top_segment_4_1.DEC1.t4 212.393
R7136 top_segment_4_1.DEC1.n1 top_segment_4_1.DEC1.t1 140.738
R7137 top_segment_4_1.DEC1.n18 top_segment_4_1.DEC1.n17 109.279
R7138 top_segment_4_1.DEC1.n19 top_segment_4_1.DEC1.n18 13.9817
R7139 top_segment_4_1.DEC1.n20 top_segment_4_1.DEC1 12.4126
R7140 top_segment_4_1.DEC1.n2 top_segment_4_1.DEC1 11.6369
R7141 top_segment_4_1.DEC1.n0 top_segment_4_1.DEC1 10.1408
R7142 top_segment_4_1.DEC1.n19 top_segment_4_1.DEC1 7.56414
R7143 top_segment_4_1.DEC1 top_segment_4_1.DEC1.n19 6.78838
R7144 top_segment_4_1.DEC1.n15 top_segment_4_1.DEC1.n14 4.5005
R7145 top_segment_4_1.DEC1.n17 top_segment_4_1.DEC1.n16 4.5005
R7146 top_segment_4_1.DEC1.n0 top_segment_4_1.DEC1 2.16154
R7147 top_segment_4_1.DEC1 top_segment_4_1.DEC1.n20 1.93989
R7148 top_segment_4_1.DEC1 top_segment_4_1.DEC1.n15 1.88512
R7149 top_segment_4_1.DEC1.n18 top_segment_4_1.DEC1 0.7755
R7150 top_segment_4_1.DEC1.n16 top_segment_4_1.DEC1 0.6755
R7151 top_segment_4_1.DEC1 top_segment_4_1.DEC1.n2 0.665435
R7152 top_segment_4_1.DEC1.n14 top_segment_4_1.DEC1.n13 0.663962
R7153 top_segment_4_1.DEC1.n13 top_segment_4_1.DEC1.n12 0.663962
R7154 top_segment_4_1.DEC1.n12 top_segment_4_1.DEC1.n11 0.663962
R7155 top_segment_4_1.DEC1.n11 top_segment_4_1.DEC1.n10 0.663962
R7156 top_segment_4_1.DEC1.n10 top_segment_4_1.DEC1.n9 0.663962
R7157 top_segment_4_1.DEC1.n4 top_segment_4_1.DEC1.n3 0.663962
R7158 top_segment_4_1.DEC1.n5 top_segment_4_1.DEC1.n4 0.663962
R7159 top_segment_4_1.DEC1.n6 top_segment_4_1.DEC1.n5 0.663962
R7160 top_segment_4_1.DEC1.n7 top_segment_4_1.DEC1.n6 0.663962
R7161 top_segment_4_1.DEC1.n8 top_segment_4_1.DEC1.n7 0.663962
R7162 top_segment_4_1.DEC1.n17 top_segment_4_1.DEC1.n8 0.663962
R7163 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t1 674.658
R7164 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t2 10.7661
R7165 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t0 10.7361
R7166 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.n0 4.09773
R7167 a_14416_5238.n0 a_14416_5238.t1 673.378
R7168 a_14416_5238.n1 a_14416_5238.t4 673.005
R7169 a_14416_5238.t0 a_14416_5238.n2 669.523
R7170 a_14416_5238.n1 a_14416_5238.t3 666.583
R7171 a_14416_5238.n0 a_14416_5238.t2 666.583
R7172 a_14416_5238.n2 a_14416_5238.n1 4.60675
R7173 a_14416_5238.n2 a_14416_5238.n0 1.95467
R7174 top_segment_3_0.bb[5].n2 top_segment_3_0.bb[5].n1 863.124
R7175 top_segment_3_0.bb[5].n1 top_segment_3_0.bb[5].n0 585
R7176 top_segment_3_0.bb[5] top_segment_3_0.bb[5].t1 495.469
R7177 top_segment_3_0.bb[5] top_segment_3_0.bb[5].t0 291.983
R7178 top_segment_3_0.bb[5].t0 top_segment_3_0.bb[5].n11 285
R7179 top_segment_3_0.bb[5].n4 top_segment_3_0.bb[5].t5 217.555
R7180 top_segment_3_0.bb[5].n4 top_segment_3_0.bb[5].t6 216.893
R7181 top_segment_3_0.bb[5].n5 top_segment_3_0.bb[5].t4 216.893
R7182 top_segment_3_0.bb[5].n3 top_segment_3_0.bb[5].t3 216.893
R7183 top_segment_3_0.bb[5].n7 top_segment_3_0.bb[5].t8 212.393
R7184 top_segment_3_0.bb[5].n9 top_segment_3_0.bb[5].n8 152
R7185 top_segment_3_0.bb[5].n1 top_segment_3_0.bb[5].t1 140.738
R7186 top_segment_3_0.bb[5].n8 top_segment_3_0.bb[5].t7 114.031
R7187 top_segment_3_0.bb[5] top_segment_3_0.bb[5].n7 93.4484
R7188 top_segment_3_0.bb[5].n8 top_segment_3_0.bb[5].t2 81.5883
R7189 top_segment_3_0.bb[5].n9 top_segment_3_0.bb[5] 16.7132
R7190 top_segment_3_0.bb[5].n10 top_segment_3_0.bb[5] 13.7979
R7191 top_segment_3_0.bb[5] top_segment_3_0.bb[5].n10 13.1884
R7192 top_segment_3_0.bb[5] top_segment_3_0.bb[5].n11 12.4126
R7193 top_segment_3_0.bb[5].n2 top_segment_3_0.bb[5] 11.6369
R7194 top_segment_3_0.bb[5].n0 top_segment_3_0.bb[5] 10.1408
R7195 top_segment_3_0.bb[5].n7 top_segment_3_0.bb[5].n6 4.5005
R7196 top_segment_3_0.bb[5].n0 top_segment_3_0.bb[5] 2.16154
R7197 top_segment_3_0.bb[5].n10 top_segment_3_0.bb[5] 2.16154
R7198 top_segment_3_0.bb[5].n11 top_segment_3_0.bb[5] 1.93989
R7199 top_segment_3_0.bb[5] top_segment_3_0.bb[5].n9 1.16414
R7200 top_segment_3_0.bb[5] top_segment_3_0.bb[5].n2 0.665435
R7201 top_segment_3_0.bb[5].n6 top_segment_3_0.bb[5].n3 0.663962
R7202 top_segment_3_0.bb[5].n6 top_segment_3_0.bb[5].n5 0.663962
R7203 top_segment_3_0.bb[5].n5 top_segment_3_0.bb[5].n4 0.663962
R7204 top_segment_3_0.bb[5].n10 top_segment_3_0.bb[5] 0.582318
R7205 top_segment_3_0.bb[5].n3 top_segment_3_0.bb[5] 0.202423
R7206 top_segment_1_0.rseg_1_v3_1.v35 top_segment_1_0.rseg_1_v3_1.v35.t2 245.728
R7207 top_segment_1_0.rseg_1_v3_1.v35.n0 top_segment_1_0.rseg_1_v3_1.v35.t0 10.5752
R7208 top_segment_1_0.rseg_1_v3_1.v35.n0 top_segment_1_0.rseg_1_v3_1.v35.t1 10.5739
R7209 top_segment_1_0.rseg_1_v3_1.v35 top_segment_1_0.rseg_1_v3_1.v35.n0 1.55257
R7210 top_segment_1_0.rseg_1_v3_1.v36 top_segment_1_0.rseg_1_v3_1.v36.t2 246.268
R7211 top_segment_1_0.rseg_1_v3_1.v36.n0 top_segment_1_0.rseg_1_v3_1.v36.t0 10.5306
R7212 top_segment_1_0.rseg_1_v3_1.v36.n0 top_segment_1_0.rseg_1_v3_1.v36.t1 10.5285
R7213 top_segment_1_0.rseg_1_v3_1.v36 top_segment_1_0.rseg_1_v3_1.v36.n0 2.15701
R7214 top_segment_1_0.rseg_1_v3_1.v18 top_segment_1_0.rseg_1_v3_1.v18.t0 247.037
R7215 top_segment_1_0.rseg_1_v3_1.v18.n0 top_segment_1_0.rseg_1_v3_1.v18.t1 10.5307
R7216 top_segment_1_0.rseg_1_v3_1.v18.n0 top_segment_1_0.rseg_1_v3_1.v18.t2 10.5285
R7217 top_segment_1_0.rseg_1_v3_1.v18 top_segment_1_0.rseg_1_v3_1.v18.n0 0.885467
R7218 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t0 230.517
R7219 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t4 229.369
R7220 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t2 229.369
R7221 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t1 157.62
R7222 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t5 157.07
R7223 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t3 157.07
R7224 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n0 152.712
R7225 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n2 152.475
R7226 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 24.2121
R7227 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n5 23.559
R7228 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 11.6875
R7229 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n1 10.2234
R7230 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n3 9.77342
R7231 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 7.23528
R7232 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 5.45235
R7233 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 5.21532
R7234 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n7 5.04292
R7235 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n6 4.73093
R7236 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n4 4.6005
R7237 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.31925
R7238 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 593.158
R7239 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 231.554
R7240 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 140.53
R7241 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 26.5955
R7242 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 26.5955
R7243 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 16.5652
R7244 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 9.03579
R7245 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 6.02403
R7246 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 1.72748
R7247 a_13900_6674.n1 a_13900_6674.t2 671.663
R7248 a_13900_6674.n0 a_13900_6674.t4 668.203
R7249 a_13900_6674.n0 a_13900_6674.t3 667.22
R7250 a_13900_6674.n1 a_13900_6674.t1 665.176
R7251 a_13900_6674.t0 a_13900_6674.n2 665.176
R7252 a_13900_6674.n2 a_13900_6674.n1 6.63383
R7253 a_13900_6674.n2 a_13900_6674.n0 4.91092
R7254 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t0 676.321
R7255 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t1 13.4699
R7256 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t2 10.7776
R7257 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.n0 4.72836
R7258 a_42781_14260.t0 a_42781_14260.t1 114.052
R7259 a_42245_13704.n0 a_42245_13704.t1 228.04
R7260 a_42245_13704.n0 a_42245_13704.t2 145.648
R7261 a_42245_13704.t0 a_42245_13704.n0 83.2159
R7262 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t0 675.929
R7263 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t2 10.8219
R7264 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t1 10.6741
R7265 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.n0 4.11026
R7266 top_segment_2_0.rseg_2_v3_0.v6.n0 top_segment_2_0.rseg_2_v3_0.v6.t1 240.188
R7267 top_segment_2_0.rseg_2_v3_0.v6.n0 top_segment_2_0.rseg_2_v3_0.v6.t2 10.5827
R7268 top_segment_2_0.rseg_2_v3_0.v6.t0 top_segment_2_0.rseg_2_v3_0.v6.n0 10.5739
R7269 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t9 230.363
R7270 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t11 230.155
R7271 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t12 229.369
R7272 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t10 212.081
R7273 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t4 212.081
R7274 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n17 203.922
R7275 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n3 186.001
R7276 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t5 158.064
R7277 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t6 157.856
R7278 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t8 157.07
R7279 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n8 155.058
R7280 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n11 154.91
R7281 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n5 152
R7282 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t7 139.78
R7283 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t13 139.78
R7284 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n0 101.49
R7285 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n2 61.346
R7286 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n9 33.2524
R7287 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n13 29.6212
R7288 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t3 26.5955
R7289 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t0 26.5955
R7290 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t1 24.9236
R7291 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t2 24.9236
R7292 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n6 20.0252
R7293 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n12 18.1725
R7294 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 13.5685
R7295 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 10.7525
R7296 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n14 9.64425
R7297 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n4 9.30224
R7298 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 6.6565
R7299 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 5.92643
R7300 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n16 5.04292
R7301 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n15 3.8405
R7302 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 3.78232
R7303 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 3.0725
R7304 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n1 2.5605
R7305 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n7 2.17042
R7306 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 1.93989
R7307 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n10 1.93214
R7308 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 1.33781
R7309 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.490734
R7310 top_segment_3_0.b[4].n2 top_segment_3_0.b[4].n1 863.124
R7311 top_segment_3_0.b[4].n1 top_segment_3_0.b[4].n0 585
R7312 top_segment_3_0.b[4] top_segment_3_0.b[4].t1 495.469
R7313 top_segment_3_0.b[4].t0 top_segment_3_0.b[4] 291.983
R7314 top_segment_3_0.b[4].n7 top_segment_3_0.b[4].t0 285
R7315 top_segment_3_0.b[4].n4 top_segment_3_0.b[4].t3 217.555
R7316 top_segment_3_0.b[4].n3 top_segment_3_0.b[4].t2 216.893
R7317 top_segment_3_0.b[4].n5 top_segment_3_0.b[4].t4 212.393
R7318 top_segment_3_0.b[4].n1 top_segment_3_0.b[4].t1 140.738
R7319 top_segment_3_0.b[4] top_segment_3_0.b[4].n5 77.7359
R7320 top_segment_3_0.b[4].n6 top_segment_3_0.b[4] 14.3755
R7321 top_segment_3_0.b[4].n7 top_segment_3_0.b[4] 12.4126
R7322 top_segment_3_0.b[4].n2 top_segment_3_0.b[4] 11.6369
R7323 top_segment_3_0.b[4].n0 top_segment_3_0.b[4] 10.1408
R7324 top_segment_3_0.b[4].n6 top_segment_3_0.b[4] 8.53383
R7325 top_segment_3_0.b[4] top_segment_3_0.b[4].n6 5.81868
R7326 top_segment_3_0.b[4].n5 top_segment_3_0.b[4].n4 4.5005
R7327 top_segment_3_0.b[4].n0 top_segment_3_0.b[4] 2.16154
R7328 top_segment_3_0.b[4] top_segment_3_0.b[4].n7 1.93989
R7329 top_segment_3_0.b[4] top_segment_3_0.b[4].n2 0.665435
R7330 top_segment_3_0.b[4].n4 top_segment_3_0.b[4].n3 0.663962
R7331 top_segment_3_0.b[4].n3 top_segment_3_0.b[4] 0.317808
R7332 a_13613_17684.n1 a_13613_17684.t2 669.294
R7333 a_13613_17684.n0 a_13613_17684.t3 666.299
R7334 a_13613_17684.n0 a_13613_17684.t1 665.667
R7335 a_13613_17684.t0 a_13613_17684.n1 665.664
R7336 a_13613_17684.n1 a_13613_17684.n0 2.7505
R7337 a_16831_17684.n0 a_16831_17684.t1 672.731
R7338 a_16831_17684.t0 a_16831_17684.n0 671.336
R7339 a_16831_17684.n0 a_16831_17684.t2 660.739
R7340 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t6 739.816
R7341 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t5 230.155
R7342 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t8 230.155
R7343 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 203.922
R7344 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t7 157.856
R7345 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t4 157.856
R7346 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 152
R7347 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 152
R7348 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 101.49
R7349 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t1 26.5955
R7350 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t0 26.5955
R7351 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 25.1816
R7352 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t3 24.9236
R7353 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t2 24.9236
R7354 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[0] 14.1609
R7355 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y 13.0565
R7356 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 12.2559
R7357 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 11.0199
R7358 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y 10.7525
R7359 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y 6.6565
R7360 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 5.10675
R7361 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 5.04292
R7362 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 4.3525
R7363 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 2.5605
R7364 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.A 2.10199
R7365 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.A 2.10199
R7366 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y 1.93989
R7367 a_43570_18104.t0 a_43570_18104.t1 49.8467
R7368 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 593.154
R7369 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 231.554
R7370 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 140.53
R7371 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 26.5955
R7372 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 26.5955
R7373 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 16.5652
R7374 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 9.03579
R7375 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 6.02403
R7376 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 1.72748
R7377 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t1 675.77
R7378 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t2 10.7383
R7379 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.t0 10.6512
R7380 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14.n0 0.682179
R7381 top_segment_1_0.rseg_1_v3_1.v25 top_segment_1_0.rseg_1_v3_1.v25.t0 249.345
R7382 top_segment_1_0.rseg_1_v3_1.v25.n0 top_segment_1_0.rseg_1_v3_1.v25.t1 10.6701
R7383 top_segment_1_0.rseg_1_v3_1.v25.n0 top_segment_1_0.rseg_1_v3_1.v25.t2 10.5739
R7384 top_segment_1_0.rseg_1_v3_1.v25 top_segment_1_0.rseg_1_v3_1.v25.n0 4.15498
R7385 top_segment_1_0.rseg_1_v3_1.v26 top_segment_1_0.rseg_1_v3_1.v26.t0 250.066
R7386 top_segment_1_0.rseg_1_v3_1.v26.n0 top_segment_1_0.rseg_1_v3_1.v26.t1 10.5296
R7387 top_segment_1_0.rseg_1_v3_1.v26.n0 top_segment_1_0.rseg_1_v3_1.v26.t2 10.5285
R7388 top_segment_1_0.rseg_1_v3_1.v26 top_segment_1_0.rseg_1_v3_1.v26.n0 3.52631
R7389 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t10 231.017
R7390 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t4 230.155
R7391 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t11 230.155
R7392 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t13 229.369
R7393 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t14 229.369
R7394 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t6 229.369
R7395 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t5 229.369
R7396 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n24 203.922
R7397 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t7 158.716
R7398 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n2 157.927
R7399 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t8 157.856
R7400 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t12 157.856
R7401 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t16 157.07
R7402 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t9 157.07
R7403 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t15 157.07
R7404 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t17 157.07
R7405 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n6 152.475
R7406 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n12 152.475
R7407 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n18 152.238
R7408 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n3 152
R7409 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n15 152
R7410 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n9 152
R7411 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n0 101.49
R7412 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t0 26.5955
R7413 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t1 26.5955
R7414 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 25.0963
R7415 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t3 24.9236
R7416 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t2 24.9236
R7417 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n20 23.8264
R7418 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n21 21.9086
R7419 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n16 19.8154
R7420 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n10 18.9229
R7421 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n7 17.1938
R7422 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n13 16.9661
R7423 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n19 15.7596
R7424 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n5 14.4113
R7425 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 13.0565
R7426 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n4 12.5635
R7427 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 10.7525
R7428 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 7.11161
R7429 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 6.6565
R7430 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 5.68939
R7431 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 5.45235
R7432 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 5.45235
R7433 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n23 5.04292
R7434 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n22 4.3525
R7435 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n1 2.5605
R7436 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 2.47068
R7437 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 2.13383
R7438 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 2.10199
R7439 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 1.93989
R7440 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n17 1.38917
R7441 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n8 1.30714
R7442 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n14 0.920422
R7443 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n11 0.900891
R7444 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.229016
R7445 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 593.396
R7446 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 231.554
R7447 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 140.53
R7448 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 26.5955
R7449 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 26.5955
R7450 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 16.5652
R7451 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 9.03579
R7452 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 6.02403
R7453 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 1.72748
R7454 DIN7.n1 DIN7.t1 212.081
R7455 DIN7.n0 DIN7.t0 212.081
R7456 DIN7.n2 DIN7.n1 183.185
R7457 DIN7.n1 DIN7.t3 139.78
R7458 DIN7.n0 DIN7.t2 139.78
R7459 DIN7.n1 DIN7.n0 61.346
R7460 DIN7 DIN7.n2 14.2776
R7461 DIN7.n2 DIN7 5.8885
R7462 top_segment_2_0.DEC0[2].n16 top_segment_2_0.DEC0[2].t1 334.788
R7463 top_segment_2_0.DEC0[2].n7 top_segment_2_0.DEC0[2].t4 213.218
R7464 top_segment_2_0.DEC0[2].n0 top_segment_2_0.DEC0[2].t2 213.218
R7465 top_segment_2_0.DEC0[2].n7 top_segment_2_0.DEC0[2].t20 212.554
R7466 top_segment_2_0.DEC0[2].n8 top_segment_2_0.DEC0[2].t5 212.554
R7467 top_segment_2_0.DEC0[2].n9 top_segment_2_0.DEC0[2].t8 212.554
R7468 top_segment_2_0.DEC0[2].n10 top_segment_2_0.DEC0[2].t6 212.554
R7469 top_segment_2_0.DEC0[2].n11 top_segment_2_0.DEC0[2].t15 212.554
R7470 top_segment_2_0.DEC0[2].n12 top_segment_2_0.DEC0[2].t10 212.554
R7471 top_segment_2_0.DEC0[2].n13 top_segment_2_0.DEC0[2].t9 212.554
R7472 top_segment_2_0.DEC0[2].n14 top_segment_2_0.DEC0[2].t16 212.554
R7473 top_segment_2_0.DEC0[2].n6 top_segment_2_0.DEC0[2].t12 212.554
R7474 top_segment_2_0.DEC0[2].n5 top_segment_2_0.DEC0[2].t17 212.554
R7475 top_segment_2_0.DEC0[2].n4 top_segment_2_0.DEC0[2].t21 212.554
R7476 top_segment_2_0.DEC0[2].n3 top_segment_2_0.DEC0[2].t13 212.554
R7477 top_segment_2_0.DEC0[2].n2 top_segment_2_0.DEC0[2].t19 212.554
R7478 top_segment_2_0.DEC0[2].n1 top_segment_2_0.DEC0[2].t11 212.554
R7479 top_segment_2_0.DEC0[2].n0 top_segment_2_0.DEC0[2].t14 212.554
R7480 top_segment_2_0.DEC0[2].n18 top_segment_2_0.DEC0[2].t7 126.27
R7481 top_segment_2_0.DEC0[2].n18 top_segment_2_0.DEC0[2].t3 125.558
R7482 top_segment_2_0.DEC0[2].n17 top_segment_2_0.DEC0[2].t18 121.127
R7483 top_segment_2_0.DEC0[2].n16 top_segment_2_0.DEC0[2].t0 87.8063
R7484 top_segment_2_0.DEC0[2] top_segment_2_0.DEC0[2].n15 81.7495
R7485 top_segment_2_0.DEC0[2].n19 top_segment_2_0.DEC0[2].n18 5.73592
R7486 top_segment_2_0.DEC0[2] top_segment_2_0.DEC0[2].n19 5.388
R7487 top_segment_2_0.DEC0[2].n14 top_segment_2_0.DEC0[2].n13 0.663962
R7488 top_segment_2_0.DEC0[2].n13 top_segment_2_0.DEC0[2].n12 0.663962
R7489 top_segment_2_0.DEC0[2].n12 top_segment_2_0.DEC0[2].n11 0.663962
R7490 top_segment_2_0.DEC0[2].n11 top_segment_2_0.DEC0[2].n10 0.663962
R7491 top_segment_2_0.DEC0[2].n10 top_segment_2_0.DEC0[2].n9 0.663962
R7492 top_segment_2_0.DEC0[2].n9 top_segment_2_0.DEC0[2].n8 0.663962
R7493 top_segment_2_0.DEC0[2].n8 top_segment_2_0.DEC0[2].n7 0.663962
R7494 top_segment_2_0.DEC0[2].n1 top_segment_2_0.DEC0[2].n0 0.663962
R7495 top_segment_2_0.DEC0[2].n2 top_segment_2_0.DEC0[2].n1 0.663962
R7496 top_segment_2_0.DEC0[2].n4 top_segment_2_0.DEC0[2].n3 0.663962
R7497 top_segment_2_0.DEC0[2].n5 top_segment_2_0.DEC0[2].n4 0.663962
R7498 top_segment_2_0.DEC0[2].n6 top_segment_2_0.DEC0[2].n5 0.663962
R7499 top_segment_2_0.DEC0[2].n15 top_segment_2_0.DEC0[2].n6 0.518014
R7500 top_segment_2_0.DEC0[2] top_segment_2_0.DEC0[2].n2 0.442808
R7501 top_segment_2_0.DEC0[2].n17 top_segment_2_0.DEC0[2].n16 0.322615
R7502 top_segment_2_0.DEC0[2].n3 top_segment_2_0.DEC0[2] 0.221654
R7503 top_segment_2_0.DEC0[2].n19 top_segment_2_0.DEC0[2].n17 0.177583
R7504 top_segment_2_0.DEC0[2].n15 top_segment_2_0.DEC0[2].n14 0.133398
R7505 a_23510_19162.n0 a_23510_19162.t1 250.252
R7506 a_23510_19162.n1 a_23510_19162.t2 245.975
R7507 a_23510_19162.t0 a_23510_19162.n1 240.382
R7508 a_23510_19162.n0 a_23510_19162.t3 240.165
R7509 a_23510_19162.n1 a_23510_19162.n0 4.27758
R7510 top_segment_2_0.rseg_2_v3_0.v39.n0 top_segment_2_0.rseg_2_v3_0.v39.t2 240.298
R7511 top_segment_2_0.rseg_2_v3_0.v39.n0 top_segment_2_0.rseg_2_v3_0.v39.t1 10.7108
R7512 top_segment_2_0.rseg_2_v3_0.v39.t0 top_segment_2_0.rseg_2_v3_0.v39.n0 10.687
R7513 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t0 274.793
R7514 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t4 230.576
R7515 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t6 230.155
R7516 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t8 229.369
R7517 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n9 205.28
R7518 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t5 158.275
R7519 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n0 157.927
R7520 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t7 157.856
R7521 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t9 157.07
R7522 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n5 153.067
R7523 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n1 152
R7524 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t1 133.124
R7525 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n10 67.4857
R7526 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n8 36.3299
R7527 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t2 26.5955
R7528 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t3 26.5955
R7529 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n4 24.8988
R7530 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n3 13.8092
R7531 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n2 12.5635
R7532 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n7 10.6878
R7533 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n6 9.3005
R7534 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 7.11161
R7535 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 5.67507
R7536 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 5.6005
R7537 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 2.13383
R7538 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.602583
R7539 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t4 230.155
R7540 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t2 229.369
R7541 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t0 221.538
R7542 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n0 157.927
R7543 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t5 157.856
R7544 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t3 157.07
R7545 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t1 152.889
R7546 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n1 152
R7547 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n3 24.6696
R7548 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n2 19.6746
R7549 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 17.3671
R7550 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n4 14.023
R7551 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 13.8127
R7552 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 2.22659
R7553 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 2.13383
R7554 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n5 1.55202
R7555 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.602583
R7556 top_segment_4_1.DEC3.n2 top_segment_4_1.DEC3.n1 863.124
R7557 top_segment_4_1.DEC3.n1 top_segment_4_1.DEC3.n0 585
R7558 top_segment_4_1.DEC3 top_segment_4_1.DEC3.t1 495.469
R7559 top_segment_4_1.DEC3.t0 top_segment_4_1.DEC3 291.983
R7560 top_segment_4_1.DEC3.n19 top_segment_4_1.DEC3.t0 285
R7561 top_segment_4_1.DEC3.n13 top_segment_4_1.DEC3.t8 217.555
R7562 top_segment_4_1.DEC3.n10 top_segment_4_1.DEC3.t15 217.555
R7563 top_segment_4_1.DEC3.n3 top_segment_4_1.DEC3.t9 217.555
R7564 top_segment_4_1.DEC3.n13 top_segment_4_1.DEC3.t11 216.893
R7565 top_segment_4_1.DEC3.n14 top_segment_4_1.DEC3.t5 216.893
R7566 top_segment_4_1.DEC3.n15 top_segment_4_1.DEC3.t3 216.893
R7567 top_segment_4_1.DEC3.n12 top_segment_4_1.DEC3.t7 216.893
R7568 top_segment_4_1.DEC3.n11 top_segment_4_1.DEC3.t6 216.893
R7569 top_segment_4_1.DEC3.n10 top_segment_4_1.DEC3.t4 216.893
R7570 top_segment_4_1.DEC3.n9 top_segment_4_1.DEC3.t2 216.893
R7571 top_segment_4_1.DEC3.n8 top_segment_4_1.DEC3.t17 216.893
R7572 top_segment_4_1.DEC3.n7 top_segment_4_1.DEC3.t16 216.893
R7573 top_segment_4_1.DEC3.n6 top_segment_4_1.DEC3.t13 216.893
R7574 top_segment_4_1.DEC3.n5 top_segment_4_1.DEC3.t12 216.893
R7575 top_segment_4_1.DEC3.n4 top_segment_4_1.DEC3.t10 216.893
R7576 top_segment_4_1.DEC3.n3 top_segment_4_1.DEC3.t14 216.893
R7577 top_segment_4_1.DEC3.n1 top_segment_4_1.DEC3.t1 140.738
R7578 top_segment_4_1.DEC3 top_segment_4_1.DEC3.n17 65.2685
R7579 top_segment_4_1.DEC3.n18 top_segment_4_1.DEC3 14.7463
R7580 top_segment_4_1.DEC3.n19 top_segment_4_1.DEC3 12.4126
R7581 top_segment_4_1.DEC3.n2 top_segment_4_1.DEC3 11.6369
R7582 top_segment_4_1.DEC3.n0 top_segment_4_1.DEC3 10.1408
R7583 top_segment_4_1.DEC3.n18 top_segment_4_1.DEC3 7.75808
R7584 top_segment_4_1.DEC3 top_segment_4_1.DEC3.n18 6.59444
R7585 top_segment_4_1.DEC3 top_segment_4_1.DEC3.n16 6.48592
R7586 top_segment_4_1.DEC3.n17 top_segment_4_1.DEC3 6.37342
R7587 top_segment_4_1.DEC3.n0 top_segment_4_1.DEC3 2.16154
R7588 top_segment_4_1.DEC3 top_segment_4_1.DEC3.n19 1.93989
R7589 top_segment_4_1.DEC3 top_segment_4_1.DEC3.n2 0.665435
R7590 top_segment_4_1.DEC3.n15 top_segment_4_1.DEC3.n14 0.663962
R7591 top_segment_4_1.DEC3.n14 top_segment_4_1.DEC3.n13 0.663962
R7592 top_segment_4_1.DEC3.n11 top_segment_4_1.DEC3.n10 0.663962
R7593 top_segment_4_1.DEC3.n12 top_segment_4_1.DEC3.n11 0.663962
R7594 top_segment_4_1.DEC3.n4 top_segment_4_1.DEC3.n3 0.663962
R7595 top_segment_4_1.DEC3.n5 top_segment_4_1.DEC3.n4 0.663962
R7596 top_segment_4_1.DEC3.n6 top_segment_4_1.DEC3.n5 0.663962
R7597 top_segment_4_1.DEC3.n7 top_segment_4_1.DEC3.n6 0.663962
R7598 top_segment_4_1.DEC3.n8 top_segment_4_1.DEC3.n7 0.663962
R7599 top_segment_4_1.DEC3.n9 top_segment_4_1.DEC3.n8 0.663962
R7600 top_segment_4_1.DEC3.n16 top_segment_4_1.DEC3.n15 0.320692
R7601 top_segment_4_1.DEC3.n16 top_segment_4_1.DEC3.n12 0.320692
R7602 top_segment_4_1.DEC3.n17 top_segment_4_1.DEC3.n9 0.274859
R7603 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t2 676.321
R7604 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t0 13.5978
R7605 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t1 10.7628
R7606 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.n0 4.72836
R7607 top_segment_1_0.rseg_1_v3_1.v33.n0 top_segment_1_0.rseg_1_v3_1.v33.t2 236.65
R7608 top_segment_1_0.rseg_1_v3_1.v33.n0 top_segment_1_0.rseg_1_v3_1.v33.t1 10.6732
R7609 top_segment_1_0.rseg_1_v3_1.v33.t0 top_segment_1_0.rseg_1_v3_1.v33.n0 10.5739
R7610 top_segment_1_0.rseg_1_v3_1.v34 top_segment_1_0.rseg_1_v3_1.v34.t2 246.804
R7611 top_segment_1_0.rseg_1_v3_1.v34.n0 top_segment_1_0.rseg_1_v3_1.v34.t1 10.6247
R7612 top_segment_1_0.rseg_1_v3_1.v34.n0 top_segment_1_0.rseg_1_v3_1.v34.t0 10.5295
R7613 top_segment_1_0.rseg_1_v3_1.v34 top_segment_1_0.rseg_1_v3_1.v34.n0 0.86158
R7614 top_segment_2_0.rseg_2_v3_0.v12.n0 top_segment_2_0.rseg_2_v3_0.v12.t1 239.088
R7615 top_segment_2_0.rseg_2_v3_0.v12.n0 top_segment_2_0.rseg_2_v3_0.v12.t2 10.5771
R7616 top_segment_2_0.rseg_2_v3_0.v12.t0 top_segment_2_0.rseg_2_v3_0.v12.n0 10.5739
R7617 top_segment_2_0.rseg_2_v3_0.v13.n0 top_segment_2_0.rseg_2_v3_0.v13.t1 238.671
R7618 top_segment_2_0.rseg_2_v3_0.v13.t0 top_segment_2_0.rseg_2_v3_0.v13.n0 10.5319
R7619 top_segment_2_0.rseg_2_v3_0.v13.n0 top_segment_2_0.rseg_2_v3_0.v13.t2 10.5285
R7620 top_segment_2_0.DEC1[3].n4 top_segment_2_0.DEC1[3].t0 334.822
R7621 top_segment_2_0.DEC1[3].n1 top_segment_2_0.DEC1[3].t8 213.218
R7622 top_segment_2_0.DEC1[3].n0 top_segment_2_0.DEC1[3].t5 213.218
R7623 top_segment_2_0.DEC1[3].n1 top_segment_2_0.DEC1[3].t4 212.554
R7624 top_segment_2_0.DEC1[3].n0 top_segment_2_0.DEC1[3].t3 212.554
R7625 top_segment_2_0.DEC1[3].n3 top_segment_2_0.DEC1[3].t7 208.054
R7626 top_segment_2_0.DEC1[3].n5 top_segment_2_0.DEC1[3].t2 126.27
R7627 top_segment_2_0.DEC1[3].n6 top_segment_2_0.DEC1[3].t9 125.558
R7628 top_segment_2_0.DEC1[3].n5 top_segment_2_0.DEC1[3].t6 125.558
R7629 top_segment_2_0.DEC1[3].n4 top_segment_2_0.DEC1[3].t1 87.8063
R7630 top_segment_2_0.DEC1[3] top_segment_2_0.DEC1[3].n3 63.3651
R7631 top_segment_2_0.DEC1[3].n7 top_segment_2_0.DEC1[3].n6 5.73592
R7632 top_segment_2_0.DEC1[3] top_segment_2_0.DEC1[3].n7 5.66196
R7633 top_segment_2_0.DEC1[3].n3 top_segment_2_0.DEC1[3].n2 4.5005
R7634 top_segment_2_0.DEC1[3].n6 top_segment_2_0.DEC1[3].n5 0.713
R7635 top_segment_2_0.DEC1[3].n2 top_segment_2_0.DEC1[3].n1 0.663962
R7636 top_segment_2_0.DEC1[3].n2 top_segment_2_0.DEC1[3] 0.457231
R7637 top_segment_2_0.DEC1[3] top_segment_2_0.DEC1[3].n0 0.207231
R7638 top_segment_2_0.DEC1[3].n7 top_segment_2_0.DEC1[3].n4 0.197295
R7639 a_41787_18542.t0 a_41787_18542.t1 65.941
R7640 top_segment_2_0.DEC1[0].n4 top_segment_2_0.DEC1[0].t1 334.771
R7641 top_segment_2_0.DEC1[0].n1 top_segment_2_0.DEC1[0].t8 213.218
R7642 top_segment_2_0.DEC1[0].n0 top_segment_2_0.DEC1[0].t6 213.218
R7643 top_segment_2_0.DEC1[0].n1 top_segment_2_0.DEC1[0].t5 212.554
R7644 top_segment_2_0.DEC1[0].n0 top_segment_2_0.DEC1[0].t3 212.554
R7645 top_segment_2_0.DEC1[0].n3 top_segment_2_0.DEC1[0].t9 208.054
R7646 top_segment_2_0.DEC1[0].n5 top_segment_2_0.DEC1[0].t2 126.278
R7647 top_segment_2_0.DEC1[0].n5 top_segment_2_0.DEC1[0].t7 125.566
R7648 top_segment_2_0.DEC1[0].n6 top_segment_2_0.DEC1[0].t4 125.566
R7649 top_segment_2_0.DEC1[0].n4 top_segment_2_0.DEC1[0].t0 87.8568
R7650 top_segment_2_0.DEC1[0] top_segment_2_0.DEC1[0].n3 65.2609
R7651 top_segment_2_0.DEC1[0] top_segment_2_0.DEC1[0].n7 5.04008
R7652 top_segment_2_0.DEC1[0].n7 top_segment_2_0.DEC1[0].n6 4.68383
R7653 top_segment_2_0.DEC1[0].n3 top_segment_2_0.DEC1[0].n2 4.5005
R7654 top_segment_2_0.DEC1[0].n7 top_segment_2_0.DEC1[0].n4 0.876942
R7655 top_segment_2_0.DEC1[0].n6 top_segment_2_0.DEC1[0].n5 0.713
R7656 top_segment_2_0.DEC1[0].n2 top_segment_2_0.DEC1[0].n1 0.663962
R7657 top_segment_2_0.DEC1[0] top_segment_2_0.DEC1[0].n0 0.363481
R7658 top_segment_2_0.DEC1[0].n2 top_segment_2_0.DEC1[0] 0.300981
R7659 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n2 270.841
R7660 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t1 258.846
R7661 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t4 241.536
R7662 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n5 224.775
R7663 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t3 169.237
R7664 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n0 152
R7665 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n1 31.0273
R7666 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t0 26.5955
R7667 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.t2 26.5955
R7668 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 3.92583
R7669 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n4 3.76521
R7670 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n3 3.03935
R7671 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 2.30266
R7672 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 1.19762
R7673 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.921363
R7674 top_segment_3_0.rseg_3_v3_0.v4.n0 top_segment_3_0.rseg_3_v3_0.v4.t1 677.225
R7675 top_segment_3_0.rseg_3_v3_0.v4.t0 top_segment_3_0.rseg_3_v3_0.v4.n0 10.7534
R7676 top_segment_3_0.rseg_3_v3_0.v4.n0 top_segment_3_0.rseg_3_v3_0.v4.t2 10.7113
R7677 top_segment_3_0.rseg_3_v3_0.v5.n0 top_segment_3_0.rseg_3_v3_0.v5.t1 677.378
R7678 top_segment_3_0.rseg_3_v3_0.v5.n0 top_segment_3_0.rseg_3_v3_0.v5.t2 10.7234
R7679 top_segment_3_0.rseg_3_v3_0.v5.t0 top_segment_3_0.rseg_3_v3_0.v5.n0 10.6693
R7680 a_26443_5238.n2 a_26443_5238.t3 247.736
R7681 a_26443_5238.n0 a_26443_5238.t4 245.752
R7682 a_26443_5238.n1 a_26443_5238.t2 245.172
R7683 a_26443_5238.n0 a_26443_5238.t1 239.083
R7684 a_26443_5238.t0 a_26443_5238.n2 239.083
R7685 a_26443_5238.n1 a_26443_5238.n0 5.85467
R7686 a_26443_5238.n2 a_26443_5238.n1 1.16717
R7687 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 593.396
R7688 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 231.554
R7689 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 140.53
R7690 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 26.5955
R7691 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 26.5955
R7692 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 16.5652
R7693 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 9.03579
R7694 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 6.02403
R7695 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 1.72748
R7696 a_42609_20641.t0 a_42609_20641.t1 129.28
R7697 a_42271_11884.t0 a_42271_11884.t1 55.3905
R7698 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t6 230.155
R7699 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t5 230.155
R7700 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t7 229.369
R7701 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t12 212.081
R7702 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t11 212.081
R7703 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n0 203.923
R7704 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n3 186.001
R7705 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n8 157.927
R7706 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t13 157.856
R7707 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t10 157.856
R7708 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t4 157.07
R7709 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n5 153.338
R7710 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n9 152
R7711 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t9 139.78
R7712 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t8 139.78
R7713 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n15 101.49
R7714 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n2 61.346
R7715 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n11 31.3499
R7716 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n12 29.8627
R7717 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t1 26.5955
R7718 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t3 26.5955
R7719 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t0 24.9236
R7720 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t2 24.9236
R7721 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n6 17.8391
R7722 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n14 13.5685
R7723 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 11.0938
R7724 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n1 10.7525
R7725 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n10 9.9845
R7726 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n13 9.64425
R7727 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n4 9.30224
R7728 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 6.6565
R7729 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 5.04292
R7730 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 3.8405
R7731 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 3.0725
R7732 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 3.05722
R7733 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 2.5605
R7734 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 2.3045
R7735 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n7 2.24073
R7736 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n16 1.93989
R7737 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.600109
R7738 a_42802_2702.t0 a_42802_2702.t1 49.8467
R7739 top_segment_1_0.rseg_1_v3_1.v2 top_segment_1_0.rseg_1_v3_1.v2.t2 248.405
R7740 top_segment_1_0.rseg_1_v3_1.v2.n0 top_segment_1_0.rseg_1_v3_1.v2.t1 10.5394
R7741 top_segment_1_0.rseg_1_v3_1.v2.n0 top_segment_1_0.rseg_1_v3_1.v2.t0 10.5295
R7742 top_segment_1_0.rseg_1_v3_1.v2 top_segment_1_0.rseg_1_v3_1.v2.n0 0.791214
R7743 top_segment_2_0.rseg_2_v3_0.v44.n0 top_segment_2_0.rseg_2_v3_0.v44.t2 239.357
R7744 top_segment_2_0.rseg_2_v3_0.v44.t0 top_segment_2_0.rseg_2_v3_0.v44.n0 10.7707
R7745 top_segment_2_0.rseg_2_v3_0.v44.n0 top_segment_2_0.rseg_2_v3_0.v44.t1 10.7309
R7746 top_segment_2_0.rseg_2_v3_0.v43.n0 top_segment_2_0.rseg_2_v3_0.v43.t2 239.483
R7747 top_segment_2_0.rseg_2_v3_0.v43.t0 top_segment_2_0.rseg_2_v3_0.v43.n0 10.7266
R7748 top_segment_2_0.rseg_2_v3_0.v43.n0 top_segment_2_0.rseg_2_v3_0.v43.t1 10.6898
R7749 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t1 673.212
R7750 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t2 10.7601
R7751 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t0 10.7161
R7752 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.n0 2.72817
R7753 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t1 673.34
R7754 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t0 10.7217
R7755 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.t2 10.6931
R7756 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22.n0 3.42321
R7757 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n7 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t6 142.488
R7758 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t9 142.488
R7759 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t11 142.488
R7760 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n7 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t10 141.704
R7761 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t13 141.704
R7762 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t12 141.704
R7763 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n6 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t8 141.704
R7764 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n5 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t7 141.704
R7765 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t4 139.454
R7766 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n9 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t2 139.454
R7767 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t1 135.329
R7768 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n11 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t3 135.231
R7769 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n11 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t5 135.231
R7770 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t0 134.444
R7771 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n5 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n4 6.41092
R7772 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.D0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n11 4.563
R7773 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n3 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n2 2.2505
R7774 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n9 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n8 2.2505
R7775 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n10 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n3 0.829667
R7776 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n10 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n9 0.829667
R7777 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n0 0.783833
R7778 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n1 0.783833
R7779 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n6 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n5 0.783833
R7780 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n8 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n6 0.783833
R7781 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n8 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n7 0.783833
R7782 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n11 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n10 0.224458
R7783 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t3 221.851
R7784 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t5 221.851
R7785 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t1 140.244
R7786 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t0 140.056
R7787 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t14 122.656
R7788 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t18 122.656
R7789 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t9 122.656
R7790 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t17 122.656
R7791 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t13 122.656
R7792 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t15 122.656
R7793 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t7 122.656
R7794 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t11 122.656
R7795 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t16 122.656
R7796 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t10 122.656
R7797 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t12 122.656
R7798 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t6 122.656
R7799 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t2 108.365
R7800 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t4 108.365
R7801 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n17 14.4346
R7802 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t8 13.3032
R7803 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n18 12.8291
R7804 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n2 11.1702
R7805 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n20 4.63108
R7806 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n0 3.9493
R7807 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n19 3.4105
R7808 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n21 2.67342
R7809 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n4 2.26409
R7810 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n1 2.25675
R7811 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n5 0.742167
R7812 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n6 0.742167
R7813 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n7 0.742167
R7814 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n15 0.742167
R7815 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n14 0.742167
R7816 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n13 0.742167
R7817 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n11 0.742167
R7818 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n10 0.742167
R7819 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n9 0.742167
R7820 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n16 0.652583
R7821 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n12 0.652583
R7822 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n1 0.546515
R7823 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n3 0.527402
R7824 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.504667
R7825 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.0900833
R7826 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.0900833
R7827 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.0650833
R7828 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n22 0.063
R7829 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.0498421
R7830 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n8 0.0255
R7831 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t2 158.145
R7832 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t1 142.477
R7833 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t0 140.496
R7834 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t3 140.082
R7835 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n0 7.35744
R7836 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n1 0.0463333
R7837 top_segment_1_0.rseg_1_v3_1.v53 top_segment_1_0.rseg_1_v3_1.v53.t2 246.63
R7838 top_segment_1_0.rseg_1_v3_1.v53.n0 top_segment_1_0.rseg_1_v3_1.v53.t0 10.6701
R7839 top_segment_1_0.rseg_1_v3_1.v53.n0 top_segment_1_0.rseg_1_v3_1.v53.t1 10.5739
R7840 top_segment_1_0.rseg_1_v3_1.v53 top_segment_1_0.rseg_1_v3_1.v53.n0 2.77493
R7841 a_27429_5238.n2 a_27429_5238.t3 248.286
R7842 a_27429_5238.n0 a_27429_5238.t4 246.303
R7843 a_27429_5238.n1 a_27429_5238.t2 244.629
R7844 a_27429_5238.n0 a_27429_5238.t1 239.633
R7845 a_27429_5238.t0 a_27429_5238.n2 239.633
R7846 a_27429_5238.n2 a_27429_5238.n1 5.93592
R7847 a_27429_5238.n1 a_27429_5238.n0 1.08592
R7848 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t1 227.856
R7849 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R7850 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t3 140.163
R7851 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t4 114.031
R7852 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t0 83.3993
R7853 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.t2 81.5883
R7854 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R7855 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R7856 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R7857 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R7858 a_42781_5984.t0 a_42781_5984.t1 114.052
R7859 top_segment_2_0.rseg_2_v3_0.v26.t0 top_segment_2_0.rseg_2_v3_0.v26.n0 239.869
R7860 top_segment_2_0.rseg_2_v3_0.v26.n0 top_segment_2_0.rseg_2_v3_0.v26.t1 10.8275
R7861 top_segment_2_0.rseg_2_v3_0.v26.n0 top_segment_2_0.rseg_2_v3_0.v26.t2 10.677
R7862 top_segment_2_0.rseg_2_v3_0.v25.n0 top_segment_2_0.rseg_2_v3_0.v25.t2 240.24
R7863 top_segment_2_0.rseg_2_v3_0.v25.t0 top_segment_2_0.rseg_2_v3_0.v25.n0 10.7836
R7864 top_segment_2_0.rseg_2_v3_0.v25.n0 top_segment_2_0.rseg_2_v3_0.v25.t1 10.6292
R7865 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 593.154
R7866 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 231.554
R7867 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 140.53
R7868 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 26.5955
R7869 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 26.5955
R7870 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 16.5652
R7871 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 9.03579
R7872 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 6.02403
R7873 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 1.72748
R7874 a_42609_19573.t0 a_42609_19573.t1 129.28
R7875 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t0 672.956
R7876 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t2 10.716
R7877 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.t1 10.6712
R7878 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52.n0 2.0484
R7879 top_segment_2_0.rseg_2_v3_0.v8.n0 top_segment_2_0.rseg_2_v3_0.v8.t1 240.773
R7880 top_segment_2_0.rseg_2_v3_0.v8.n0 top_segment_2_0.rseg_2_v3_0.v8.t2 13.9942
R7881 top_segment_2_0.rseg_2_v3_0.v8.t0 top_segment_2_0.rseg_2_v3_0.v8.n0 11.0596
R7882 top_segment_2_0.rseg_2_v3_0.v7.n0 top_segment_2_0.rseg_2_v3_0.v7.t1 243.41
R7883 top_segment_2_0.rseg_2_v3_0.v7.t0 top_segment_2_0.rseg_2_v3_0.v7.n0 10.5372
R7884 top_segment_2_0.rseg_2_v3_0.v7.n0 top_segment_2_0.rseg_2_v3_0.v7.t2 10.5285
R7885 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t4 228.463
R7886 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n5 224.775
R7887 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t3 157.07
R7888 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n2 152
R7889 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t2 132.067
R7890 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n3 30.3559
R7891 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t1 26.5955
R7892 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.t0 26.5955
R7893 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 4.20621
R7894 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n0 4.15748
R7895 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n1 2.25932
R7896 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n4 1.50638
R7897 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 1.17559
R7898 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A 0.921363
R7899 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t1 227.856
R7900 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n2 152.333
R7901 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t2 140.382
R7902 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t3 114.031
R7903 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t0 83.3993
R7904 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.t4 81.5883
R7905 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n3 14.4422
R7906 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n1 7.56882
R7907 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n0 5.08175
R7908 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R7909 a_42271_16280.t0 a_42271_16280.t1 55.3905
R7910 a_42245_15684.n0 a_42245_15684.t1 228.04
R7911 a_42245_15684.n0 a_42245_15684.t2 145.648
R7912 a_42245_15684.t0 a_42245_15684.n0 83.2159
R7913 a_43890_3526.t0 a_43890_3526.t1 49.8467
R7914 a_43890_3610.t0 a_43890_3610.t1 60.9236
R7915 top_segment_1_0.rseg_1_v3_1.v31.t0 top_segment_1_0.rseg_1_v3_1.v31.n0 240.469
R7916 top_segment_1_0.rseg_1_v3_1.v31.n0 top_segment_1_0.rseg_1_v3_1.v31.t1 10.6701
R7917 top_segment_1_0.rseg_1_v3_1.v31.n0 top_segment_1_0.rseg_1_v3_1.v31.t2 10.5739
R7918 top_segment_1_0.rseg_1_v3_1.v32.n0 top_segment_1_0.rseg_1_v3_1.v32.t1 241.547
R7919 top_segment_1_0.rseg_1_v3_1.v32.t0 top_segment_1_0.rseg_1_v3_1.v32.n0 12.1531
R7920 top_segment_1_0.rseg_1_v3_1.v32.n0 top_segment_1_0.rseg_1_v3_1.v32.t2 12.0758
R7921 top_segment_3_0.rseg_3_v3_0.v12.t0 top_segment_3_0.rseg_3_v3_0.v12.n0 679.261
R7922 top_segment_3_0.rseg_3_v3_0.v12.n0 top_segment_3_0.rseg_3_v3_0.v12.t1 10.7728
R7923 top_segment_3_0.rseg_3_v3_0.v12.n0 top_segment_3_0.rseg_3_v3_0.v12.t2 10.7357
R7924 top_segment_3_0.rseg_3_v3_0.v13.n0 top_segment_3_0.rseg_3_v3_0.v13.t2 676.942
R7925 top_segment_3_0.rseg_3_v3_0.v13.t0 top_segment_3_0.rseg_3_v3_0.v13.n0 10.7308
R7926 top_segment_3_0.rseg_3_v3_0.v13.n0 top_segment_3_0.rseg_3_v3_0.v13.t1 10.6636
R7927 a_17823_7938.n0 a_17823_7938.t1 670.519
R7928 a_17823_7938.n0 a_17823_7938.t2 670.183
R7929 a_17823_7938.t0 a_17823_7938.n0 666.073
R7930 a_14452_6674.n0 a_14452_6674.t3 672.03
R7931 a_14452_6674.t0 a_14452_6674.n2 668.37
R7932 a_14452_6674.n2 a_14452_6674.t4 666.942
R7933 a_14452_6674.n0 a_14452_6674.t2 665.543
R7934 a_14452_6674.n1 a_14452_6674.t1 665.543
R7935 a_14452_6674.n1 a_14452_6674.n0 6.63383
R7936 a_14452_6674.n2 a_14452_6674.n1 4.12758
R7937 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t1 673.212
R7938 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t0 10.7577
R7939 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t2 10.7161
R7940 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.n0 2.72817
R7941 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t2 673.412
R7942 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t0 10.7213
R7943 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.t1 10.6898
R7944 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38.n0 3.42178
R7945 top_segment_2_0.rseg_2_v3_0.v2.n0 top_segment_2_0.rseg_2_v3_0.v2.t2 238.046
R7946 top_segment_2_0.rseg_2_v3_0.v2.t0 top_segment_2_0.rseg_2_v3_0.v2.n0 10.7009
R7947 top_segment_2_0.rseg_2_v3_0.v2.n0 top_segment_2_0.rseg_2_v3_0.v2.t1 10.5739
R7948 top_segment_2_0.rseg_2_v3_0.v1.n0 top_segment_2_0.rseg_2_v3_0.v1.t1 240.27
R7949 top_segment_2_0.rseg_2_v3_0.v1.t0 top_segment_2_0.rseg_2_v3_0.v1.n0 10.6702
R7950 top_segment_2_0.rseg_2_v3_0.v1.n0 top_segment_2_0.rseg_2_v3_0.v1.t2 10.5285
R7951 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t3 593.154
R7952 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 231.554
R7953 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t1 140.53
R7954 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t0 26.5955
R7955 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.t2 26.5955
R7956 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 16.5652
R7957 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 9.03579
R7958 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n1 6.02403
R7959 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 1.72748
R7960 a_42609_20997.t0 a_42609_20997.t1 129.28
R7961 a_13154_5238.n0 a_13154_5238.t1 672.644
R7962 a_13154_5238.n1 a_13154_5238.t4 672.27
R7963 a_13154_5238.t0 a_13154_5238.n2 671.963
R7964 a_13154_5238.n1 a_13154_5238.t3 665.85
R7965 a_13154_5238.n0 a_13154_5238.t2 665.85
R7966 a_13154_5238.n2 a_13154_5238.n0 5.78175
R7967 a_13154_5238.n2 a_13154_5238.n1 0.779667
R7968 a_18099_7938.n0 a_18099_7938.t1 670.775
R7969 a_18099_7938.n0 a_18099_7938.t2 670.366
R7970 a_18099_7938.t0 a_18099_7938.n0 665.89
R7971 a_41938_2230.t0 a_41938_2230.t1 49.8467
R7972 a_41938_2314.t0 a_41938_2314.t1 60.9236
R7973 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 272.038
R7974 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t2 258.846
R7975 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t4 228.463
R7976 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n5 224.775
R7977 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t3 157.07
R7978 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n0 153.28
R7979 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t1 26.5955
R7980 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.t0 26.5955
R7981 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n1 21.3673
R7982 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n4 3.76521
R7983 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n3 3.03935
R7984 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 2.92621
R7985 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n2 1.56597
R7986 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A 0.921363
R7987 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A.n2 0.737191
R7988 a_28879_6674.n2 a_28879_6674.t3 246.244
R7989 a_28879_6674.n0 a_28879_6674.t4 241.385
R7990 a_28879_6674.n0 a_28879_6674.t1 240.358
R7991 a_28879_6674.n1 a_28879_6674.t2 238.959
R7992 a_28879_6674.t0 a_28879_6674.n2 238.959
R7993 a_28879_6674.n2 a_28879_6674.n1 6.788
R7994 a_28879_6674.n1 a_28879_6674.n0 4.15675
R7995 top_segment_1_0.rseg_1_v3_1.v42 top_segment_1_0.rseg_1_v3_1.v42.t2 249.947
R7996 top_segment_1_0.rseg_1_v3_1.v42.n0 top_segment_1_0.rseg_1_v3_1.v42.t1 10.5296
R7997 top_segment_1_0.rseg_1_v3_1.v42.n0 top_segment_1_0.rseg_1_v3_1.v42.t0 10.5295
R7998 top_segment_1_0.rseg_1_v3_1.v42 top_segment_1_0.rseg_1_v3_1.v42.n0 3.5287
R7999 a_15438_6674.n0 a_15438_6674.t3 672.581
R8000 a_15438_6674.t0 a_15438_6674.n2 670.423
R8001 a_15438_6674.n2 a_15438_6674.t4 666.391
R8002 a_15438_6674.n0 a_15438_6674.t2 666.092
R8003 a_15438_6674.n1 a_15438_6674.t1 666.092
R8004 a_15438_6674.n1 a_15438_6674.n0 6.63383
R8005 a_15438_6674.n2 a_15438_6674.n1 2.62342
R8006 a_18493_7938.t0 a_18493_7938.n0 671.561
R8007 a_18493_7938.n0 a_18493_7938.t2 671.109
R8008 a_18493_7938.n0 a_18493_7938.t1 665.524
R8009 top_segment_1_0.rseg_1_v3_1.v21 top_segment_1_0.rseg_1_v3_1.v21.t0 246.63
R8010 top_segment_1_0.rseg_1_v3_1.v21.n0 top_segment_1_0.rseg_1_v3_1.v21.t1 10.6701
R8011 top_segment_1_0.rseg_1_v3_1.v21.n0 top_segment_1_0.rseg_1_v3_1.v21.t2 10.5739
R8012 top_segment_1_0.rseg_1_v3_1.v21 top_segment_1_0.rseg_1_v3_1.v21.n0 2.78018
R8013 top_segment_2_0.rseg_2_v3_0.v22.n0 top_segment_2_0.rseg_2_v3_0.v22.t1 240.143
R8014 top_segment_2_0.rseg_2_v3_0.v22.t0 top_segment_2_0.rseg_2_v3_0.v22.n0 10.575
R8015 top_segment_2_0.rseg_2_v3_0.v22.n0 top_segment_2_0.rseg_2_v3_0.v22.t2 10.5739
R8016 top_segment_2_0.rseg_2_v3_0.v23.n0 top_segment_2_0.rseg_2_v3_0.v23.t2 240.311
R8017 top_segment_2_0.rseg_2_v3_0.v23.n0 top_segment_2_0.rseg_2_v3_0.v23.t1 10.6058
R8018 top_segment_2_0.rseg_2_v3_0.v23.t0 top_segment_2_0.rseg_2_v3_0.v23.n0 10.6
R8019 a_41529_17802.t0 a_41529_17802.t1 65.941
R8020 a_41787_17802.t0 a_41787_17802.t1 65.941
R8021 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n0 267.599
R8022 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t5 230.155
R8023 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n3 196.889
R8024 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t6 157.856
R8025 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n1 152
R8026 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t1 132.982
R8027 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n5 62.4946
R8028 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t0 32.5055
R8029 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t2 32.5055
R8030 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n2 30.2423
R8031 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t3 26.5955
R8032 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.t4 26.5955
R8033 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n4 5.2056
R8034 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n6 4.04261
R8035 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A 2.3045
R8036 top_segment_2_0.rseg_2_v3_0.v40.n0 top_segment_2_0.rseg_2_v3_0.v40.t2 240.804
R8037 top_segment_2_0.rseg_2_v3_0.v40.t0 top_segment_2_0.rseg_2_v3_0.v40.n0 13.9904
R8038 top_segment_2_0.rseg_2_v3_0.v40.n0 top_segment_2_0.rseg_2_v3_0.v40.t1 10.8053
R8039 top_segment_2_0.rseg_2_v3_0.v36.n0 top_segment_2_0.rseg_2_v3_0.v36.t2 238.819
R8040 top_segment_2_0.rseg_2_v3_0.v36.t0 top_segment_2_0.rseg_2_v3_0.v36.n0 10.758
R8041 top_segment_2_0.rseg_2_v3_0.v36.n0 top_segment_2_0.rseg_2_v3_0.v36.t1 10.7137
R8042 top_segment_2_0.rseg_2_v3_0.v35.n0 top_segment_2_0.rseg_2_v3_0.v35.t2 238.345
R8043 top_segment_2_0.rseg_2_v3_0.v35.n0 top_segment_2_0.rseg_2_v3_0.v35.t1 10.7398
R8044 top_segment_2_0.rseg_2_v3_0.v35.t0 top_segment_2_0.rseg_2_v3_0.v35.n0 10.6498
R8045 top_segment_1_0.rseg_1_v3_1.v8 top_segment_1_0.rseg_1_v3_1.v8.t1 249.738
R8046 top_segment_1_0.rseg_1_v3_1.v8.n0 top_segment_1_0.rseg_1_v3_1.v8.t0 13.5854
R8047 top_segment_1_0.rseg_1_v3_1.v8.n0 top_segment_1_0.rseg_1_v3_1.v8.t2 10.8954
R8048 top_segment_1_0.rseg_1_v3_1.v8 top_segment_1_0.rseg_1_v3_1.v8.n0 4.7255
R8049 DIN6.n1 DIN6.t1 212.081
R8050 DIN6.n0 DIN6.t0 212.081
R8051 DIN6.n2 DIN6.n1 183.185
R8052 DIN6.n1 DIN6.t3 139.78
R8053 DIN6.n0 DIN6.t2 139.78
R8054 DIN6.n1 DIN6.n0 61.346
R8055 DIN6 DIN6.n2 14.2776
R8056 DIN6.n2 DIN6 5.8885
R8057 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t14 738.899
R8058 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t10 241.536
R8059 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t19 232.214
R8060 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t8 232.214
R8061 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t9 229.369
R8062 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t20 229.369
R8063 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t5 229.369
R8064 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t13 212.081
R8065 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t11 212.081
R8066 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 203.922
R8067 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 186.001
R8068 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t7 169.237
R8069 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t12 159.915
R8070 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t4 159.915
R8071 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t15 157.07
R8072 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t6 157.07
R8073 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t16 157.07
R8074 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 155.88
R8075 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 154.065
R8076 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 152.712
R8077 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 152.475
R8078 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 152
R8079 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 152
R8080 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t18 139.78
R8081 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t17 139.78
R8082 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 101.49
R8083 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 61.346
R8084 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t1 26.5955
R8085 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t0 26.5955
R8086 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t3 24.9236
R8087 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t2 24.9236
R8088 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 23.417
R8089 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 21.961
R8090 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 20.0025
R8091 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 18.2158
R8092 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 15.6884
R8093 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y 13.5685
R8094 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 12.4213
R8095 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[0] 11.8734
R8096 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 10.9817
R8097 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y 10.7525
R8098 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 10.2234
R8099 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 9.77342
R8100 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 9.64425
R8101 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 9.30224
R8102 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x2.C 6.98232
R8103 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y 6.6565
R8104 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x1.B 5.92643
R8105 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.B 5.45235
R8106 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.B 5.21532
R8107 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 5.04292
R8108 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 4.91925
R8109 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 3.8405
R8110 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.A 3.0725
R8111 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.A 2.68437
R8112 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 2.5605
R8113 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 2.30909
R8114 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y 1.93989
R8115 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 1.42823
R8116 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.A 0.970197
R8117 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 0.623547
R8118 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[6] 0.451672
R8119 a_43890_2518.t0 a_43890_2518.t1 49.8467
R8120 a_41529_20308.t0 a_41529_20308.t1 65.941
R8121 a_41787_20308.t0 a_41787_20308.t1 65.941
R8122 DIN4.n1 DIN4.t0 212.081
R8123 DIN4.n0 DIN4.t3 212.081
R8124 DIN4.n2 DIN4.n1 183.185
R8125 DIN4.n1 DIN4.t2 139.78
R8126 DIN4.n0 DIN4.t1 139.78
R8127 DIN4.n1 DIN4.n0 61.346
R8128 DIN4 DIN4.n2 14.2776
R8129 DIN4.n2 DIN4 5.8885
R8130 top_segment_1_0.rseg_1_v3_1.v7 top_segment_1_0.rseg_1_v3_1.v7.t1 248.075
R8131 top_segment_1_0.rseg_1_v3_1.v7.n0 top_segment_1_0.rseg_1_v3_1.v7.t2 10.5773
R8132 top_segment_1_0.rseg_1_v3_1.v7.n0 top_segment_1_0.rseg_1_v3_1.v7.t0 10.5739
R8133 top_segment_1_0.rseg_1_v3_1.v7 top_segment_1_0.rseg_1_v3_1.v7.n0 4.31612
R8134 top_segment_1_0.rseg_1_v3_1.v20 top_segment_1_0.rseg_1_v3_1.v20.t0 246.501
R8135 top_segment_1_0.rseg_1_v3_1.v20.n0 top_segment_1_0.rseg_1_v3_1.v20.t2 10.5309
R8136 top_segment_1_0.rseg_1_v3_1.v20.n0 top_segment_1_0.rseg_1_v3_1.v20.t1 10.5285
R8137 top_segment_1_0.rseg_1_v3_1.v20 top_segment_1_0.rseg_1_v3_1.v20.n0 2.14784
R8138 top_segment_1_0.rseg_1_v3_1.v48.n0 top_segment_1_0.rseg_1_v3_1.v48.t2 241.547
R8139 top_segment_1_0.rseg_1_v3_1.v48.t0 top_segment_1_0.rseg_1_v3_1.v48.n0 12.1331
R8140 top_segment_1_0.rseg_1_v3_1.v48.n0 top_segment_1_0.rseg_1_v3_1.v48.t1 12.0758
R8141 a_41787_17460.t0 a_41787_17460.t1 65.941
R8142 a_29589_6674.n2 a_29589_6674.t3 246.612
R8143 a_29589_6674.n0 a_29589_6674.t4 242.863
R8144 a_29589_6674.n0 a_29589_6674.t1 239.639
R8145 a_29589_6674.n1 a_29589_6674.t2 239.326
R8146 a_29589_6674.t0 a_29589_6674.n2 239.326
R8147 a_29589_6674.n2 a_29589_6674.n1 6.788
R8148 a_29589_6674.n1 a_29589_6674.n0 3.04425
R8149 top_segment_2_0.rseg_2_v3_0.v34.n0 top_segment_2_0.rseg_2_v3_0.v34.t2 237.841
R8150 top_segment_2_0.rseg_2_v3_0.v34.t0 top_segment_2_0.rseg_2_v3_0.v34.n0 10.7808
R8151 top_segment_2_0.rseg_2_v3_0.v34.n0 top_segment_2_0.rseg_2_v3_0.v34.t1 10.6951
R8152 top_segment_2_0.rseg_2_v3_0.v33.n0 top_segment_2_0.rseg_2_v3_0.v33.t2 237.419
R8153 top_segment_2_0.rseg_2_v3_0.v33.n0 top_segment_2_0.rseg_2_v3_0.v33.t1 10.6247
R8154 top_segment_2_0.rseg_2_v3_0.v33.t0 top_segment_2_0.rseg_2_v3_0.v33.n0 10.5295
R8155 top_segment_2_0.DEC0[1].n17 top_segment_2_0.DEC0[1].t0 334.771
R8156 top_segment_2_0.DEC0[1].n8 top_segment_2_0.DEC0[1].t4 213.218
R8157 top_segment_2_0.DEC0[1].n8 top_segment_2_0.DEC0[1].t11 212.554
R8158 top_segment_2_0.DEC0[1].n9 top_segment_2_0.DEC0[1].t2 212.554
R8159 top_segment_2_0.DEC0[1].n10 top_segment_2_0.DEC0[1].t14 212.554
R8160 top_segment_2_0.DEC0[1].n11 top_segment_2_0.DEC0[1].t18 212.554
R8161 top_segment_2_0.DEC0[1].n12 top_segment_2_0.DEC0[1].t3 212.554
R8162 top_segment_2_0.DEC0[1].n13 top_segment_2_0.DEC0[1].t16 212.554
R8163 top_segment_2_0.DEC0[1].n14 top_segment_2_0.DEC0[1].t6 212.554
R8164 top_segment_2_0.DEC0[1].n15 top_segment_2_0.DEC0[1].t13 212.554
R8165 top_segment_2_0.DEC0[1].n7 top_segment_2_0.DEC0[1].t19 212.554
R8166 top_segment_2_0.DEC0[1].n6 top_segment_2_0.DEC0[1].t8 212.554
R8167 top_segment_2_0.DEC0[1].n5 top_segment_2_0.DEC0[1].t15 212.554
R8168 top_segment_2_0.DEC0[1].n4 top_segment_2_0.DEC0[1].t5 212.554
R8169 top_segment_2_0.DEC0[1].n3 top_segment_2_0.DEC0[1].t9 212.554
R8170 top_segment_2_0.DEC0[1].n2 top_segment_2_0.DEC0[1].t21 212.554
R8171 top_segment_2_0.DEC0[1].n1 top_segment_2_0.DEC0[1].t7 212.554
R8172 top_segment_2_0.DEC0[1].n0 top_segment_2_0.DEC0[1].t17 212.554
R8173 top_segment_2_0.DEC0[1].n20 top_segment_2_0.DEC0[1].t10 131.306
R8174 top_segment_2_0.DEC0[1].n18 top_segment_2_0.DEC0[1].t12 126.278
R8175 top_segment_2_0.DEC0[1].n18 top_segment_2_0.DEC0[1].t20 125.566
R8176 top_segment_2_0.DEC0[1].n17 top_segment_2_0.DEC0[1].t1 87.8231
R8177 top_segment_2_0.DEC0[1] top_segment_2_0.DEC0[1].n16 71.2205
R8178 top_segment_2_0.DEC0[1] top_segment_2_0.DEC0[1].n20 5.12863
R8179 top_segment_2_0.DEC0[1].n19 top_segment_2_0.DEC0[1].n18 4.68383
R8180 top_segment_2_0.DEC0[1].n15 top_segment_2_0.DEC0[1].n14 0.663962
R8181 top_segment_2_0.DEC0[1].n14 top_segment_2_0.DEC0[1].n13 0.663962
R8182 top_segment_2_0.DEC0[1].n13 top_segment_2_0.DEC0[1].n12 0.663962
R8183 top_segment_2_0.DEC0[1].n12 top_segment_2_0.DEC0[1].n11 0.663962
R8184 top_segment_2_0.DEC0[1].n11 top_segment_2_0.DEC0[1].n10 0.663962
R8185 top_segment_2_0.DEC0[1].n10 top_segment_2_0.DEC0[1].n9 0.663962
R8186 top_segment_2_0.DEC0[1].n9 top_segment_2_0.DEC0[1].n8 0.663962
R8187 top_segment_2_0.DEC0[1].n1 top_segment_2_0.DEC0[1].n0 0.663962
R8188 top_segment_2_0.DEC0[1].n2 top_segment_2_0.DEC0[1].n1 0.663962
R8189 top_segment_2_0.DEC0[1].n3 top_segment_2_0.DEC0[1].n2 0.663962
R8190 top_segment_2_0.DEC0[1].n4 top_segment_2_0.DEC0[1].n3 0.663962
R8191 top_segment_2_0.DEC0[1].n5 top_segment_2_0.DEC0[1].n4 0.663962
R8192 top_segment_2_0.DEC0[1].n6 top_segment_2_0.DEC0[1].n5 0.663962
R8193 top_segment_2_0.DEC0[1].n7 top_segment_2_0.DEC0[1].n6 0.663962
R8194 top_segment_2_0.DEC0[1].n19 top_segment_2_0.DEC0[1].n17 0.608192
R8195 top_segment_2_0.DEC0[1].n16 top_segment_2_0.DEC0[1].n7 0.542052
R8196 top_segment_2_0.DEC0[1].n0 top_segment_2_0.DEC0[1] 0.238481
R8197 top_segment_2_0.DEC0[1].n20 top_segment_2_0.DEC0[1].n19 0.177583
R8198 top_segment_2_0.DEC0[1].n16 top_segment_2_0.DEC0[1].n15 0.10936
R8199 a_19646_19162.n1 a_19646_19162.t1 251.536
R8200 a_19646_19162.n0 a_19646_19162.t3 250.017
R8201 a_19646_19162.t0 a_19646_19162.n1 241.447
R8202 a_19646_19162.n0 a_19646_19162.t2 239.1
R8203 a_19646_19162.n1 a_19646_19162.n0 1.51925
R8204 top_segment_2_0.rseg_2_v3_0.v30.t0 top_segment_2_0.rseg_2_v3_0.v30.n0 237.898
R8205 top_segment_2_0.rseg_2_v3_0.v30.n0 top_segment_2_0.rseg_2_v3_0.v30.t2 10.786
R8206 top_segment_2_0.rseg_2_v3_0.v30.n0 top_segment_2_0.rseg_2_v3_0.v30.t1 10.6951
R8207 a_41271_19226.t0 a_41271_19226.t1 65.941
R8208 top_segment_3_0.b[6].n2 top_segment_3_0.b[6].n1 863.124
R8209 top_segment_3_0.b[6].n1 top_segment_3_0.b[6].n0 585
R8210 top_segment_3_0.b[6] top_segment_3_0.b[6].t1 495.469
R8211 top_segment_3_0.b[6].t0 top_segment_3_0.b[6] 291.983
R8212 top_segment_3_0.b[6].n13 top_segment_3_0.b[6].t0 285
R8213 top_segment_3_0.b[6].n3 top_segment_3_0.b[6].t2 217.555
R8214 top_segment_3_0.b[6].n3 top_segment_3_0.b[6].t7 216.893
R8215 top_segment_3_0.b[6].n4 top_segment_3_0.b[6].t8 216.893
R8216 top_segment_3_0.b[6].n5 top_segment_3_0.b[6].t3 216.893
R8217 top_segment_3_0.b[6].n6 top_segment_3_0.b[6].t9 216.893
R8218 top_segment_3_0.b[6].n7 top_segment_3_0.b[6].t4 216.893
R8219 top_segment_3_0.b[6].n8 top_segment_3_0.b[6].t6 216.893
R8220 top_segment_3_0.b[6].n9 top_segment_3_0.b[6].t10 216.893
R8221 top_segment_3_0.b[6].n10 top_segment_3_0.b[6].t5 216.893
R8222 top_segment_3_0.b[6].n1 top_segment_3_0.b[6].t1 140.738
R8223 top_segment_3_0.b[6] top_segment_3_0.b[6].n11 79.1581
R8224 top_segment_3_0.b[6].n12 top_segment_3_0.b[6] 14.3755
R8225 top_segment_3_0.b[6].n13 top_segment_3_0.b[6] 12.4126
R8226 top_segment_3_0.b[6].n2 top_segment_3_0.b[6] 11.6369
R8227 top_segment_3_0.b[6].n0 top_segment_3_0.b[6] 10.1408
R8228 top_segment_3_0.b[6].n12 top_segment_3_0.b[6] 8.53383
R8229 top_segment_3_0.b[6] top_segment_3_0.b[6].n12 5.81868
R8230 top_segment_3_0.b[6].n0 top_segment_3_0.b[6] 2.16154
R8231 top_segment_3_0.b[6] top_segment_3_0.b[6].n13 1.93989
R8232 top_segment_3_0.b[6] top_segment_3_0.b[6].n2 0.665435
R8233 top_segment_3_0.b[6].n10 top_segment_3_0.b[6].n9 0.663962
R8234 top_segment_3_0.b[6].n9 top_segment_3_0.b[6].n8 0.663962
R8235 top_segment_3_0.b[6].n8 top_segment_3_0.b[6].n7 0.663962
R8236 top_segment_3_0.b[6].n7 top_segment_3_0.b[6].n6 0.663962
R8237 top_segment_3_0.b[6].n6 top_segment_3_0.b[6].n5 0.663962
R8238 top_segment_3_0.b[6].n5 top_segment_3_0.b[6].n4 0.663962
R8239 top_segment_3_0.b[6].n4 top_segment_3_0.b[6].n3 0.663962
R8240 top_segment_3_0.b[6].n11 top_segment_3_0.b[6].n10 0.284841
R8241 top_segment_3_0.b[6].n11 top_segment_3_0.b[6] 0.0250536
R8242 a_15162_6674.n0 a_15162_6674.t3 672.396
R8243 a_15162_6674.t0 a_15162_6674.n2 669.848
R8244 a_15162_6674.n2 a_15162_6674.t4 666.222
R8245 a_15162_6674.n0 a_15162_6674.t2 665.909
R8246 a_15162_6674.n1 a_15162_6674.t1 665.909
R8247 a_15162_6674.n1 a_15162_6674.n0 6.63383
R8248 a_15162_6674.n2 a_15162_6674.n1 3.01508
R8249 top_segment_4_1.V0.n1 top_segment_4_1.V0.t3 668.534
R8250 top_segment_4_1.V0.n0 top_segment_4_1.V0.t1 668.481
R8251 top_segment_4_1.V0.n0 top_segment_4_1.V0.t2 11.7556
R8252 top_segment_4_1.V0.t0 top_segment_4_1.V0.n1 10.6569
R8253 top_segment_4_1.V0.n1 top_segment_4_1.V0.n0 5.86455
R8254 a_13645_18854.t0 a_13645_18854.n0 670.881
R8255 a_13645_18854.n0 a_13645_18854.t2 668.149
R8256 a_13645_18854.n0 a_13645_18854.t1 665.133
R8257 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t1 675.814
R8258 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t0 10.7162
R8259 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t2 10.6712
R8260 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.n0 2.05317
R8261 VH2.n0 VH2.t2 244.607
R8262 VH2.n2 VH2.t3 239.264
R8263 VH2.n1 VH2.t1 239.264
R8264 VH2.n0 VH2.t0 234.399
R8265 VH2.n1 VH2.n0 6.0755
R8266 VH2 VH2.n1 1.09842
R8267 VH2 VH2.n2 0.110917
R8268 VH2.n2 VH2 0.063
R8269 a_22176_17121.n0 a_22176_17121.t1 241.998
R8270 a_22176_17121.t0 a_22176_17121.n3 239.899
R8271 a_22176_17121.n3 a_22176_17121.t3 239.264
R8272 a_22176_17121.n2 a_22176_17121.t4 239.065
R8273 a_22176_17121.n1 a_22176_17121.t5 239.065
R8274 a_22176_17121.n0 a_22176_17121.t2 239.065
R8275 a_22176_17121.n1 a_22176_17121.n0 2.93383
R8276 a_22176_17121.n2 a_22176_17121.n1 2.93383
R8277 a_22176_17121.n3 a_22176_17121.n2 2.7755
R8278 a_17271_7938.n0 a_17271_7938.t1 670.153
R8279 a_17271_7938.n0 a_17271_7938.t2 669.817
R8280 a_17271_7938.t0 a_17271_7938.n0 666.441
R8281 a_42802_2150.t0 a_42802_2150.t1 49.8467
R8282 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n2 271.668
R8283 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t2 258.846
R8284 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t4 228.649
R8285 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n5 224.775
R8286 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t3 156.35
R8287 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n0 152
R8288 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n1 35.7621
R8289 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t1 26.5955
R8290 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.t0 26.5955
R8291 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 6.13383
R8292 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n4 3.76521
R8293 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n3 3.03935
R8294 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 2.30266
R8295 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.921363
R8296 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A 0.368845
R8297 a_22406_19162.n1 a_22406_19162.t3 248.969
R8298 a_22406_19162.n0 a_22406_19162.t2 246.287
R8299 a_22406_19162.n0 a_22406_19162.t1 241.666
R8300 a_22406_19162.t0 a_22406_19162.n1 238.881
R8301 a_22406_19162.n1 a_22406_19162.n0 2.68175
R8302 top_segment_2_0.V0.n0 top_segment_2_0.V0.t0 237.625
R8303 top_segment_2_0.V0.n1 top_segment_2_0.V0.t2 15.5067
R8304 top_segment_2_0.V0.n0 top_segment_2_0.V0.t1 10.6569
R8305 top_segment_2_0.V0.n1 top_segment_2_0.V0.n0 2.49239
R8306 top_segment_2_0.V0 top_segment_2_0.V0.n1 0.252408
R8307 a_33403_7938.n0 a_33403_7938.t2 246.133
R8308 a_33403_7938.n0 a_33403_7938.t1 244.286
R8309 a_33403_7938.t0 a_33403_7938.n0 238.756
R8310 top_segment_3_0.rseg_3_v3_0.v10.n0 top_segment_3_0.rseg_3_v3_0.v10.t2 680.375
R8311 top_segment_3_0.rseg_3_v3_0.v10.n0 top_segment_3_0.rseg_3_v3_0.v10.t1 10.7835
R8312 top_segment_3_0.rseg_3_v3_0.v10.t0 top_segment_3_0.rseg_3_v3_0.v10.n0 10.6741
R8313 top_segment_3_0.rseg_3_v3_0.v9.n0 top_segment_3_0.rseg_3_v3_0.v9.t2 677.731
R8314 top_segment_3_0.rseg_3_v3_0.v9.t0 top_segment_3_0.rseg_3_v3_0.v9.n0 10.7394
R8315 top_segment_3_0.rseg_3_v3_0.v9.n0 top_segment_3_0.rseg_3_v3_0.v9.t1 10.6292
R8316 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t4 757.36
R8317 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t5 212.081
R8318 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t6 212.081
R8319 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 203.923
R8320 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 186.001
R8321 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t7 139.78
R8322 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t8 139.78
R8323 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 101.49
R8324 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 61.346
R8325 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t1 26.5955
R8326 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t2 26.5955
R8327 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t3 24.9236
R8328 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t0 24.9236
R8329 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 13.5685
R8330 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 10.7525
R8331 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 9.64425
R8332 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 9.30224
R8333 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y 6.6565
R8334 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y 5.04292
R8335 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y 3.8405
R8336 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.A 3.0725
R8337 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y 2.5605
R8338 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 1.93989
R8339 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t4 766.463
R8340 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 203.923
R8341 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 101.49
R8342 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t0 26.5955
R8343 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t1 26.5955
R8344 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t2 24.9236
R8345 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t3 24.9236
R8346 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y 13.0565
R8347 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y 10.7525
R8348 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y 6.6565
R8349 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 5.04292
R8350 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 4.3525
R8351 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 2.5605
R8352 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y 1.93989
R8353 a_18899_9019.n0 a_18899_9019.t1 668.659
R8354 a_18899_9019.n0 a_18899_9019.t2 668.024
R8355 a_18899_9019.t0 a_18899_9019.n0 665.667
R8356 a_35435_18774.n4 a_35435_18774.t0 239.399
R8357 a_35435_18774.t1 a_35435_18774.n4 227.651
R8358 a_35435_18774.n0 a_35435_18774.t5 222.332
R8359 a_35435_18774.n2 a_35435_18774.t3 222.332
R8360 a_35435_18774.n1 a_35435_18774.t7 111.007
R8361 a_35435_18774.n3 a_35435_18774.t6 111.007
R8362 a_35435_18774.n0 a_35435_18774.t4 108.365
R8363 a_35435_18774.n2 a_35435_18774.t2 108.365
R8364 a_35435_18774.n1 a_35435_18774.n0 2.64217
R8365 a_35435_18774.n3 a_35435_18774.n2 2.64217
R8366 a_35435_18774.n3 a_35435_18774.n1 0.817167
R8367 a_35435_18774.n4 a_35435_18774.n3 0.302583
R8368 a_42245_8754.t0 a_42245_8754.n0 228.04
R8369 a_42245_8754.n0 a_42245_8754.t2 145.648
R8370 a_42245_8754.n0 a_42245_8754.t1 83.2159
R8371 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t4 241.536
R8372 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n5 224.775
R8373 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t3 169.237
R8374 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n1 153.032
R8375 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t1 132.067
R8376 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n2 32.3107
R8377 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t0 26.5955
R8378 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.t2 26.5955
R8379 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 24.8072
R8380 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n4 3.76521
R8381 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n0 2.77619
R8382 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n3 1.38179
R8383 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 1.17559
R8384 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.921363
R8385 top_segment_4_1.bb1.n2 top_segment_4_1.bb1.n1 863.124
R8386 top_segment_4_1.bb1.n1 top_segment_4_1.bb1.n0 585
R8387 top_segment_4_1.bb1 top_segment_4_1.bb1.t1 495.469
R8388 top_segment_4_1.bb1 top_segment_4_1.bb1.t0 291.983
R8389 top_segment_4_1.bb1.t0 top_segment_4_1.bb1.n10 285
R8390 top_segment_4_1.bb1.n3 top_segment_4_1.bb1.t2 216.893
R8391 top_segment_4_1.bb1 top_segment_4_1.bb1.t6 213.042
R8392 top_segment_4_1.bb1.n4 top_segment_4_1.bb1.t3 212.393
R8393 top_segment_4_1.bb1.n5 top_segment_4_1.bb1.t5 208.054
R8394 top_segment_4_1.bb1.n8 top_segment_4_1.bb1.n7 152
R8395 top_segment_4_1.bb1.n1 top_segment_4_1.bb1.t1 140.738
R8396 top_segment_4_1.bb1.n7 top_segment_4_1.bb1.t4 114.031
R8397 top_segment_4_1.bb1.n7 top_segment_4_1.bb1.t7 81.5883
R8398 top_segment_4_1.bb1.n6 top_segment_4_1.bb1.n4 43.6755
R8399 top_segment_4_1.bb1 top_segment_4_1.bb1.n6 25.5255
R8400 top_segment_4_1.bb1.n8 top_segment_4_1.bb1 16.7132
R8401 top_segment_4_1.bb1.n9 top_segment_4_1.bb1 13.7979
R8402 top_segment_4_1.bb1 top_segment_4_1.bb1.n9 13.1884
R8403 top_segment_4_1.bb1 top_segment_4_1.bb1.n10 12.4126
R8404 top_segment_4_1.bb1.n2 top_segment_4_1.bb1 11.6369
R8405 top_segment_4_1.bb1.n6 top_segment_4_1.bb1.n5 11.0276
R8406 top_segment_4_1.bb1.n0 top_segment_4_1.bb1 10.1408
R8407 top_segment_4_1.bb1.n4 top_segment_4_1.bb1.n3 5.16396
R8408 top_segment_4_1.bb1.n5 top_segment_4_1.bb1 4.67598
R8409 top_segment_4_1.bb1.n0 top_segment_4_1.bb1 2.16154
R8410 top_segment_4_1.bb1.n9 top_segment_4_1.bb1 2.16154
R8411 top_segment_4_1.bb1.n10 top_segment_4_1.bb1 1.93989
R8412 top_segment_4_1.bb1 top_segment_4_1.bb1.n8 1.16414
R8413 top_segment_4_1.bb1 top_segment_4_1.bb1.n2 0.665435
R8414 top_segment_4_1.bb1.n9 top_segment_4_1.bb1 0.582318
R8415 top_segment_4_1.bb1.n3 top_segment_4_1.bb1 0.166365
R8416 a_18319_9019.n0 a_18319_9019.t2 666.712
R8417 a_18319_9019.t0 a_18319_9019.n0 666.096
R8418 a_18319_9019.n0 a_18319_9019.t1 665.505
R8419 a_33116_9019.n0 a_33116_9019.t1 240.108
R8420 a_33116_9019.t0 a_33116_9019.n0 239.733
R8421 a_33116_9019.n0 a_33116_9019.t2 238.899
R8422 a_41271_17802.t0 a_41271_17802.t1 65.941
R8423 top_segment_1_0.rseg_1_v3_1.v59 top_segment_1_0.rseg_1_v3_1.v59.t1 248.95
R8424 top_segment_1_0.rseg_1_v3_1.v59.n0 top_segment_1_0.rseg_1_v3_1.v59.t0 10.6701
R8425 top_segment_1_0.rseg_1_v3_1.v59.n0 top_segment_1_0.rseg_1_v3_1.v59.t2 10.5739
R8426 top_segment_1_0.rseg_1_v3_1.v59 top_segment_1_0.rseg_1_v3_1.v59.n0 2.77016
R8427 top_segment_1_0.rseg_1_v3_1.v60 top_segment_1_0.rseg_1_v3_1.v60.t1 249.148
R8428 top_segment_1_0.rseg_1_v3_1.v60.n0 top_segment_1_0.rseg_1_v3_1.v60.t2 10.6247
R8429 top_segment_1_0.rseg_1_v3_1.v60.n0 top_segment_1_0.rseg_1_v3_1.v60.t0 10.5295
R8430 top_segment_1_0.rseg_1_v3_1.v60 top_segment_1_0.rseg_1_v3_1.v60.n0 2.09277
R8431 a_21026_19162.n1 a_21026_19162.t1 250.619
R8432 a_21026_19162.n0 a_21026_19162.t2 249.733
R8433 a_21026_19162.t0 a_21026_19162.n1 240.531
R8434 a_21026_19162.n0 a_21026_19162.t3 240.016
R8435 a_21026_19162.n1 a_21026_19162.n0 0.885917
R8436 top_segment_2_0.rseg_2_v3_0.v9.n0 top_segment_2_0.rseg_2_v3_0.v9.t1 240.44
R8437 top_segment_2_0.rseg_2_v3_0.v9.t0 top_segment_2_0.rseg_2_v3_0.v9.n0 10.534
R8438 top_segment_2_0.rseg_2_v3_0.v9.n0 top_segment_2_0.rseg_2_v3_0.v9.t2 10.5285
R8439 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t6 739.265
R8440 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t5 230.155
R8441 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t9 229.369
R8442 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t12 212.081
R8443 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t11 212.081
R8444 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 203.922
R8445 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 186.001
R8446 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 157.927
R8447 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t8 157.856
R8448 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t10 157.07
R8449 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 152
R8450 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t7 139.78
R8451 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t4 139.78
R8452 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 101.49
R8453 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 61.346
R8454 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t3 26.5955
R8455 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t0 26.5955
R8456 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t1 24.9236
R8457 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t2 24.9236
R8458 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 19.6746
R8459 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 19.6318
R8460 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.B 14.4147
R8461 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y 13.5685
R8462 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[1] 11.5193
R8463 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y 10.7525
R8464 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 9.64425
R8465 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 9.30224
R8466 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y 6.6565
R8467 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 5.04292
R8468 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 3.8405
R8469 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.A 3.0725
R8470 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 2.5605
R8471 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.A 2.13383
R8472 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y 1.93989
R8473 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t6 739.449
R8474 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t7 230.155
R8475 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t4 229.369
R8476 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 203.922
R8477 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 157.927
R8478 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t8 157.856
R8479 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t5 157.07
R8480 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 152
R8481 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 101.49
R8482 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 28.9524
R8483 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t1 26.5955
R8484 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t0 26.5955
R8485 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t3 24.9236
R8486 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t2 24.9236
R8487 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 14.4113
R8488 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y 13.0565
R8489 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 12.5635
R8490 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[1] 12.4026
R8491 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y 10.7525
R8492 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.B 7.11161
R8493 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y 6.6565
R8494 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 5.04292
R8495 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 4.3525
R8496 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 2.5605
R8497 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.A 2.13383
R8498 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y 1.93989
R8499 top_segment_1_0.rseg_1_v3_1.v29 top_segment_1_0.rseg_1_v3_1.v29.t0 249.321
R8500 top_segment_1_0.rseg_1_v3_1.v29.n0 top_segment_1_0.rseg_1_v3_1.v29.t1 10.6701
R8501 top_segment_1_0.rseg_1_v3_1.v29.n0 top_segment_1_0.rseg_1_v3_1.v29.t2 10.5739
R8502 top_segment_1_0.rseg_1_v3_1.v29 top_segment_1_0.rseg_1_v3_1.v29.n0 1.54779
R8503 a_29865_6674.n2 a_29865_6674.t3 246.794
R8504 a_29865_6674.n0 a_29865_6674.t4 243.439
R8505 a_29865_6674.n0 a_29865_6674.t1 239.809
R8506 a_29865_6674.n1 a_29865_6674.t2 239.51
R8507 a_29865_6674.t0 a_29865_6674.n2 239.51
R8508 a_29865_6674.n2 a_29865_6674.n1 6.788
R8509 a_29865_6674.n1 a_29865_6674.n0 2.65258
R8510 a_20474_19162.n1 a_20474_19162.t1 251.352
R8511 a_20474_19162.n0 a_20474_19162.t3 248.684
R8512 a_20474_19162.t0 a_20474_19162.n1 241.264
R8513 a_20474_19162.n0 a_20474_19162.t2 239.282
R8514 a_20474_19162.n1 a_20474_19162.n0 2.66925
R8515 top_segment_2_0.rseg_2_v3_0.v29.t0 top_segment_2_0.rseg_2_v3_0.v29.n0 238.269
R8516 top_segment_2_0.rseg_2_v3_0.v29.n0 top_segment_2_0.rseg_2_v3_0.v29.t2 10.7341
R8517 top_segment_2_0.rseg_2_v3_0.v29.n0 top_segment_2_0.rseg_2_v3_0.v29.t1 10.6516
R8518 a_41271_20308.t0 a_41271_20308.t1 65.941
R8519 DIN1.n1 DIN1.t3 212.081
R8520 DIN1.n0 DIN1.t2 212.081
R8521 DIN1.n2 DIN1.n1 183.185
R8522 DIN1.n1 DIN1.t1 139.78
R8523 DIN1.n0 DIN1.t0 139.78
R8524 DIN1.n1 DIN1.n0 61.346
R8525 DIN1 DIN1.n2 14.2776
R8526 DIN1.n2 DIN1 5.8885
R8527 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t2 672.309
R8528 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t1 10.7857
R8529 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.t0 10.6946
R8530 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19.n0 1.3567
R8531 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t2 673.259
R8532 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t1 10.7368
R8533 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.t0 10.6531
R8534 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18.n0 0.682657
R8535 a_14140_5238.n0 a_14140_5238.t1 673.193
R8536 a_14140_5238.n1 a_14140_5238.t4 672.821
R8537 a_14140_5238.t0 a_14140_5238.n2 670.087
R8538 a_14140_5238.n1 a_14140_5238.t3 666.399
R8539 a_14140_5238.n0 a_14140_5238.t2 666.399
R8540 a_14140_5238.n2 a_14140_5238.n1 4.99842
R8541 a_14140_5238.n2 a_14140_5238.n0 1.563
R8542 top_segment_2_0.DEC1[1].n4 top_segment_2_0.DEC1[1].t1 334.771
R8543 top_segment_2_0.DEC1[1].n1 top_segment_2_0.DEC1[1].t3 213.218
R8544 top_segment_2_0.DEC1[1] top_segment_2_0.DEC1[1].t6 212.989
R8545 top_segment_2_0.DEC1[1].n1 top_segment_2_0.DEC1[1].t5 212.554
R8546 top_segment_2_0.DEC1[1].n0 top_segment_2_0.DEC1[1].t4 212.554
R8547 top_segment_2_0.DEC1[1].n3 top_segment_2_0.DEC1[1].t9 208.054
R8548 top_segment_2_0.DEC1[1].n7 top_segment_2_0.DEC1[1].t8 131.306
R8549 top_segment_2_0.DEC1[1].n5 top_segment_2_0.DEC1[1].t2 126.278
R8550 top_segment_2_0.DEC1[1].n5 top_segment_2_0.DEC1[1].t7 125.566
R8551 top_segment_2_0.DEC1[1].n4 top_segment_2_0.DEC1[1].t0 87.8231
R8552 top_segment_2_0.DEC1[1] top_segment_2_0.DEC1[1].n3 56.8068
R8553 top_segment_2_0.DEC1[1] top_segment_2_0.DEC1[1].n7 5.12863
R8554 top_segment_2_0.DEC1[1].n6 top_segment_2_0.DEC1[1].n5 4.68383
R8555 top_segment_2_0.DEC1[1].n3 top_segment_2_0.DEC1[1].n2 4.5005
R8556 top_segment_2_0.DEC1[1].n2 top_segment_2_0.DEC1[1].n0 0.663962
R8557 top_segment_2_0.DEC1[1].n2 top_segment_2_0.DEC1[1].n1 0.663962
R8558 top_segment_2_0.DEC1[1].n6 top_segment_2_0.DEC1[1].n4 0.608192
R8559 top_segment_2_0.DEC1[1].n0 top_segment_2_0.DEC1[1] 0.228865
R8560 top_segment_2_0.DEC1[1].n7 top_segment_2_0.DEC1[1].n6 0.177583
R8561 a_41529_19568.t0 a_41529_19568.t1 65.941
R8562 a_41787_19568.t0 a_41787_19568.t1 65.941
R8563 a_42271_8360.t0 a_42271_8360.t1 55.3905
R8564 a_42271_15844.t0 a_42271_15844.t1 55.3905
R8565 top_segment_1_0.rseg_1_v3_1.v17.t0 top_segment_1_0.rseg_1_v3_1.v17.n0 236.649
R8566 top_segment_1_0.rseg_1_v3_1.v17.n0 top_segment_1_0.rseg_1_v3_1.v17.t2 10.6701
R8567 top_segment_1_0.rseg_1_v3_1.v17.n0 top_segment_1_0.rseg_1_v3_1.v17.t1 10.5739
R8568 a_13495_17684.t0 a_13495_17684.n0 671.708
R8569 a_13495_17684.n0 a_13495_17684.t1 667.766
R8570 a_13495_17684.n0 a_13495_17684.t2 666.221
R8571 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t1 675.904
R8572 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t0 10.7856
R8573 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.t2 10.6951
R8574 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13.n0 1.35718
R8575 DIN0.n1 DIN0.t1 212.081
R8576 DIN0.n0 DIN0.t0 212.081
R8577 DIN0.n2 DIN0.n1 183.185
R8578 DIN0.n1 DIN0.t3 139.78
R8579 DIN0.n0 DIN0.t2 139.78
R8580 DIN0.n1 DIN0.n0 61.346
R8581 DIN0 DIN0.n2 14.2776
R8582 DIN0.n2 DIN0 5.8885
R8583 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t7 761.269
R8584 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t5 212.081
R8585 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t4 212.081
R8586 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 203.922
R8587 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 186.001
R8588 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t8 139.78
R8589 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t6 139.78
R8590 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 101.49
R8591 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 61.346
R8592 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t1 26.5955
R8593 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t0 26.5955
R8594 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t3 24.9236
R8595 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t2 24.9236
R8596 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y 13.5685
R8597 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y 10.7525
R8598 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 9.64425
R8599 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 9.30224
R8600 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y 6.6565
R8601 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 5.04292
R8602 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 3.8405
R8603 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.A 3.0725
R8604 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 2.5605
R8605 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y 1.93989
R8606 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t1 227.856
R8607 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R8608 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t4 140.163
R8609 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t2 114.031
R8610 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t0 83.3993
R8611 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.t3 81.5883
R8612 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R8613 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R8614 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R8615 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R8616 SH[2].n2 SH[2].n1 863.124
R8617 SH[2].n1 SH[2].n0 585
R8618 SH[2] SH[2].t1 495.469
R8619 SH[2].n3 SH[2].t0 141.189
R8620 SH[2].n1 SH[2].t1 140.738
R8621 SH[2] SH[2].n4 14.5776
R8622 SH[2].n2 SH[2] 11.6369
R8623 SH[2].n0 SH[2] 10.1408
R8624 SH[2].n4 SH[2] 8.14595
R8625 SH[2] SH[2].n3 7.94225
R8626 SH[2].n4 SH[2] 6.20656
R8627 SH[2].n3 SH[2] 6.14988
R8628 SH[2].n0 SH[2] 2.16154
R8629 SH[2] SH[2].n2 0.665435
R8630 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t3 232.214
R8631 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n0 191.1
R8632 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t4 159.915
R8633 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n1 152
R8634 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t1 140.53
R8635 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n3 46.4787
R8636 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n2 36.7299
R8637 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t0 26.5955
R8638 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.t2 26.5955
R8639 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 16.5652
R8640 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n4 9.03579
R8641 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 2.27147
R8642 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A 1.72748
R8643 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t1 227.856
R8644 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n2 152.333
R8645 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t2 140.382
R8646 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t4 114.031
R8647 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t0 83.3993
R8648 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.t3 81.5883
R8649 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n3 14.4422
R8650 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n1 7.56882
R8651 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n0 5.08175
R8652 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R8653 a_42781_9944.t0 a_42781_9944.t1 114.052
R8654 a_42245_7764.n0 a_42245_7764.t1 228.04
R8655 a_42245_7764.n0 a_42245_7764.t2 145.648
R8656 a_42245_7764.t0 a_42245_7764.n0 83.2159
R8657 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t1 227.856
R8658 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R8659 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t4 140.163
R8660 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t2 114.031
R8661 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t0 83.3993
R8662 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.t3 81.5883
R8663 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R8664 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R8665 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R8666 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R8667 a_42271_7924.t0 a_42271_7924.t1 55.3905
R8668 a_13864_5238.n0 a_13864_5238.t1 673.01
R8669 a_13864_5238.n1 a_13864_5238.t4 672.638
R8670 a_13864_5238.t0 a_13864_5238.n2 670.662
R8671 a_13864_5238.n1 a_13864_5238.t3 666.216
R8672 a_13864_5238.n0 a_13864_5238.t2 666.216
R8673 a_13864_5238.n2 a_13864_5238.n1 5.39008
R8674 a_13864_5238.n2 a_13864_5238.n0 1.17133
R8675 a_20740_17121.n0 a_20740_17121.t1 244.489
R8676 a_20740_17121.n2 a_20740_17121.t2 242.548
R8677 a_20740_17121.n0 a_20740_17121.t3 239.614
R8678 a_20740_17121.n1 a_20740_17121.t4 239.614
R8679 a_20740_17121.t0 a_20740_17121.n2 239.614
R8680 a_20740_17121.n2 a_20740_17121.n1 2.93383
R8681 a_20740_17121.n1 a_20740_17121.n0 2.93383
R8682 a_21854_19162.n2 a_21854_19162.t4 249.702
R8683 a_21854_19162.n0 a_21854_19162.t1 248.171
R8684 a_21854_19162.n1 a_21854_19162.t2 240.933
R8685 a_21854_19162.n0 a_21854_19162.t3 240.933
R8686 a_21854_19162.t0 a_21854_19162.n2 239.614
R8687 a_21854_19162.n2 a_21854_19162.n1 0.898417
R8688 a_21854_19162.n1 a_21854_19162.n0 0.633833
R8689 a_27153_5238.n2 a_27153_5238.t3 248.102
R8690 a_27153_5238.n0 a_27153_5238.t4 246.119
R8691 a_27153_5238.n1 a_27153_5238.t2 245.203
R8692 a_27153_5238.n0 a_27153_5238.t1 239.45
R8693 a_27153_5238.t0 a_27153_5238.n2 239.45
R8694 a_27153_5238.n2 a_27153_5238.n1 6.32758
R8695 a_27153_5238.n1 a_27153_5238.n0 0.69425
R8696 top_segment_4_1.bb0.n2 top_segment_4_1.bb0.n1 863.124
R8697 top_segment_4_1.bb0.n1 top_segment_4_1.bb0.n0 585
R8698 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y top_segment_4_1.bb0.t1 495.469
R8699 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y top_segment_4_1.bb0.t0 291.983
R8700 top_segment_4_1.bb0.t0 top_segment_4_1.bb0.n8 285
R8701 top_segment_4_1.bb0.n4 top_segment_4_1.bb0.t2 255.121
R8702 top_segment_4_1.bb0.n3 top_segment_4_1.bb0.t5 208.054
R8703 top_segment_4_1.bb0.n6 top_segment_4_1.bb0.n5 152
R8704 top_segment_4_1.bb0.n1 top_segment_4_1.bb0.t1 140.738
R8705 top_segment_4_1.bb0.n5 top_segment_4_1.bb0.t3 114.031
R8706 top_segment_4_1.bb0.n5 top_segment_4_1.bb0.t4 81.5883
R8707 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.bb[0] top_segment_4_1.bb0.n4 29.0609
R8708 top_segment_4_1.bb0.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUTB 16.7132
R8709 top_segment_4_1.bb0.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.A 13.7979
R8710 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y top_segment_4_1.bb0.n7 13.1884
R8711 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y top_segment_4_1.bb0.n8 12.4126
R8712 top_segment_4_1.bb0.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 11.6369
R8713 top_segment_4_1.bb0.n4 top_segment_4_1.bb0.n3 10.6609
R8714 top_segment_4_1.bb0.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 10.1408
R8715 top_segment_4_1.bb0.n3 top_segment_1_0.bb[0] 4.5606
R8716 top_segment_4_1.bb0.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 2.16154
R8717 top_segment_4_1.bb0.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 2.16154
R8718 top_segment_4_1.bb0.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 1.93989
R8719 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.A top_segment_4_1.bb0.n6 1.16414
R8720 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y top_segment_4_1.bb0.n2 0.665435
R8721 top_segment_4_1.bb0.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y 0.582318
R8722 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUTB top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.bb[0] 0.185917
R8723 VS4.n0 VS4.t0 665.933
R8724 VS4.n0 VS4.t1 665.299
R8725 VS4 VS4.n0 0.063
R8726 a_18015_9019.n0 a_18015_9019.t2 666.692
R8727 a_18015_9019.n0 a_18015_9019.t1 666.317
R8728 a_18015_9019.t0 a_18015_9019.n0 665.484
R8729 top_segment_1_0.rseg_1_v3_1.v1.n0 top_segment_1_0.rseg_1_v3_1.v1.t2 236.657
R8730 top_segment_1_0.rseg_1_v3_1.v1.n0 top_segment_1_0.rseg_1_v3_1.v1.t1 10.6906
R8731 top_segment_1_0.rseg_1_v3_1.v1.t0 top_segment_1_0.rseg_1_v3_1.v1.n0 10.5739
R8732 a_42781_7964.t0 a_42781_7964.t1 114.052
R8733 a_41271_18144.t0 a_41271_18144.t1 65.941
R8734 a_27981_5238.n2 a_27981_5238.t3 248.653
R8735 a_27981_5238.n0 a_27981_5238.t4 246.668
R8736 a_27981_5238.n1 a_27981_5238.t2 243.488
R8737 a_27981_5238.n0 a_27981_5238.t1 240
R8738 a_27981_5238.t0 a_27981_5238.n2 240
R8739 a_27981_5238.n2 a_27981_5238.n1 5.15258
R8740 a_27981_5238.n1 a_27981_5238.n0 1.86925
R8741 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t0 676.005
R8742 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t2 10.7345
R8743 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.t1 10.6512
R8744 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46.n0 0.683611
R8745 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t4 241.536
R8746 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n5 224.775
R8747 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t3 169.237
R8748 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n2 152
R8749 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t1 132.067
R8750 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n3 31.596
R8751 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t0 26.5955
R8752 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.t2 26.5955
R8753 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 22.9652
R8754 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n0 4.15748
R8755 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 3.87418
R8756 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n1 3.76521
R8757 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n4 2.63579
R8758 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 1.17559
R8759 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.921363
R8760 a_43570_18700.t0 a_43570_18700.t1 49.8467
R8761 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t2 663.232
R8762 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t1 10.6713
R8763 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v17.n0 10.5739
R8764 top_segment_1_0.rseg_1_v3_1.v24 top_segment_1_0.rseg_1_v3_1.v24.t0 249.738
R8765 top_segment_1_0.rseg_1_v3_1.v24.n0 top_segment_1_0.rseg_1_v3_1.v24.t2 13.5018
R8766 top_segment_1_0.rseg_1_v3_1.v24.n0 top_segment_1_0.rseg_1_v3_1.v24.t1 10.7924
R8767 top_segment_1_0.rseg_1_v3_1.v24 top_segment_1_0.rseg_1_v3_1.v24.n0 4.72836
R8768 top_segment_2_0.rseg_2_v3_0.v11.n0 top_segment_2_0.rseg_2_v3_0.v11.t2 239.53
R8769 top_segment_2_0.rseg_2_v3_0.v11.t0 top_segment_2_0.rseg_2_v3_0.v11.n0 10.534
R8770 top_segment_2_0.rseg_2_v3_0.v11.n0 top_segment_2_0.rseg_2_v3_0.v11.t1 10.5285
R8771 top_segment_1_0.rseg_1_v3_1.v52 top_segment_1_0.rseg_1_v3_1.v52.t2 246.18
R8772 top_segment_1_0.rseg_1_v3_1.v52.n0 top_segment_1_0.rseg_1_v3_1.v52.t0 10.5306
R8773 top_segment_1_0.rseg_1_v3_1.v52.n0 top_segment_1_0.rseg_1_v3_1.v52.t1 10.5285
R8774 top_segment_1_0.rseg_1_v3_1.v52 top_segment_1_0.rseg_1_v3_1.v52.n0 2.14387
R8775 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t1 674.658
R8776 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t0 10.7625
R8777 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t2 10.7309
R8778 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.n0 4.09058
R8779 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t4 769.742
R8780 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 203.923
R8781 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 101.49
R8782 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t1 26.5955
R8783 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t0 26.5955
R8784 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t3 24.9236
R8785 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t2 24.9236
R8786 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y 13.0565
R8787 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y 10.7525
R8788 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y 6.6565
R8789 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 5.04292
R8790 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 4.3525
R8791 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 2.5605
R8792 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y 1.93989
R8793 a_42781_10300.t0 a_42781_10300.t1 114.052
R8794 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t2 675.741
R8795 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t0 10.7136
R8796 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t1 10.6722
R8797 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.n0 2.0546
R8798 a_41938_2146.t0 a_41938_2146.t1 49.8467
R8799 top_segment_1_0.rseg_1_v3_1.v4 top_segment_1_0.rseg_1_v3_1.v4.t1 247.869
R8800 top_segment_1_0.rseg_1_v3_1.v4.n0 top_segment_1_0.rseg_1_v3_1.v4.t2 10.5339
R8801 top_segment_1_0.rseg_1_v3_1.v4.n0 top_segment_1_0.rseg_1_v3_1.v4.t0 10.5295
R8802 top_segment_1_0.rseg_1_v3_1.v4 top_segment_1_0.rseg_1_v3_1.v4.n0 2.21785
R8803 top_segment_2_0.rseg_2_v3_0.v46.n0 top_segment_2_0.rseg_2_v3_0.v46.t2 238.37
R8804 top_segment_2_0.rseg_2_v3_0.v46.n0 top_segment_2_0.rseg_2_v3_0.v46.t1 10.7799
R8805 top_segment_2_0.rseg_2_v3_0.v46.t0 top_segment_2_0.rseg_2_v3_0.v46.n0 10.7013
R8806 a_41271_19568.t0 a_41271_19568.t1 65.941
R8807 a_14165_17684.n0 a_14165_17684.t2 671.716
R8808 a_14165_17684.n0 a_14165_17684.t1 667.361
R8809 a_14165_17684.t0 a_14165_17684.n0 666.032
R8810 a_22682_19162.n1 a_22682_19162.t3 249.153
R8811 a_22682_19162.n0 a_22682_19162.t1 247.62
R8812 a_22682_19162.n0 a_22682_19162.t2 241.482
R8813 a_22682_19162.t0 a_22682_19162.n1 239.065
R8814 a_22682_19162.n1 a_22682_19162.n0 1.53175
R8815 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t1 227.856
R8816 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n0 153.165
R8817 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t3 140.163
R8818 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t4 114.031
R8819 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t0 83.3993
R8820 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.t2 81.5883
R8821 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n2 21.9959
R8822 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 10.1408
R8823 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n3 5.81868
R8824 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A.n1 5.3005
R8825 SH[4].n2 SH[4].n1 863.124
R8826 SH[4].n1 SH[4].n0 585
R8827 SH[4] SH[4].t1 495.469
R8828 SH[4].n3 SH[4].t0 141.189
R8829 SH[4].n1 SH[4].t1 140.738
R8830 SH[4] SH[4].n4 14.5776
R8831 SH[4].n2 SH[4] 11.6369
R8832 SH[4].n0 SH[4] 10.1408
R8833 SH[4].n4 SH[4] 8.14595
R8834 SH[4] SH[4].n3 7.94225
R8835 SH[4].n4 SH[4] 6.20656
R8836 SH[4].n3 SH[4] 6.14988
R8837 SH[4].n0 SH[4] 2.16154
R8838 SH[4] SH[4].n2 0.665435
R8839 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t1 667.052
R8840 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.n0 10.6701
R8841 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v15.t2 10.5739
R8842 a_15990_6674.n0 a_15990_6674.t3 672.947
R8843 a_15990_6674.t0 a_15990_6674.n2 671.573
R8844 a_15990_6674.n2 a_15990_6674.t4 666.919
R8845 a_15990_6674.n0 a_15990_6674.t2 666.46
R8846 a_15990_6674.n1 a_15990_6674.t1 666.46
R8847 a_15990_6674.n1 a_15990_6674.n0 6.63383
R8848 a_15990_6674.n2 a_15990_6674.n1 1.84008
R8849 top_segment_2_0.rseg_2_v3_0.v24.t0 top_segment_2_0.rseg_2_v3_0.v24.n0 240.931
R8850 top_segment_2_0.rseg_2_v3_0.v24.n0 top_segment_2_0.rseg_2_v3_0.v24.t1 13.8869
R8851 top_segment_2_0.rseg_2_v3_0.v24.n0 top_segment_2_0.rseg_2_v3_0.v24.t2 10.8444
R8852 top_segment_1_0.rseg_1_v3_1.v45 top_segment_1_0.rseg_1_v3_1.v45.t1 249.321
R8853 top_segment_1_0.rseg_1_v3_1.v45.n0 top_segment_1_0.rseg_1_v3_1.v45.t2 10.6671
R8854 top_segment_1_0.rseg_1_v3_1.v45.n0 top_segment_1_0.rseg_1_v3_1.v45.t0 10.5769
R8855 top_segment_1_0.rseg_1_v3_1.v45 top_segment_1_0.rseg_1_v3_1.v45.n0 1.55078
R8856 DIN9.n1 DIN9.t3 212.081
R8857 DIN9.n0 DIN9.t1 212.081
R8858 DIN9.n2 DIN9.n1 183.185
R8859 DIN9.n1 DIN9.t2 139.78
R8860 DIN9.n0 DIN9.t0 139.78
R8861 DIN9.n1 DIN9.n0 61.346
R8862 DIN9 DIN9.n2 14.2776
R8863 DIN9.n2 DIN9 5.8885
R8864 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t3 593.165
R8865 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 237.577
R8866 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t1 140.53
R8867 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t0 26.5955
R8868 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.t2 26.5955
R8869 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 16.5652
R8870 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 9.03579
R8871 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 1.72748
R8872 DIN3.n1 DIN3.t0 212.081
R8873 DIN3.n0 DIN3.t3 212.081
R8874 DIN3.n2 DIN3.n1 183.185
R8875 DIN3.n1 DIN3.t2 139.78
R8876 DIN3.n0 DIN3.t1 139.78
R8877 DIN3.n1 DIN3.n0 61.346
R8878 DIN3 DIN3.n2 14.3234
R8879 DIN3.n2 DIN3 5.8885
R8880 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t6 752.088
R8881 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t5 212.081
R8882 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t4 212.081
R8883 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 203.922
R8884 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 186.001
R8885 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t8 139.78
R8886 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t7 139.78
R8887 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 101.49
R8888 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 61.346
R8889 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t0 26.5955
R8890 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t1 26.5955
R8891 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t3 24.9236
R8892 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t2 24.9236
R8893 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y 13.5685
R8894 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y 10.7525
R8895 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 9.64425
R8896 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 9.30224
R8897 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y 6.6565
R8898 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 5.04292
R8899 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 3.8405
R8900 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.A 3.0725
R8901 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 2.5605
R8902 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y 1.93989
R8903 a_25891_5238.n2 a_25891_5238.t3 247.369
R8904 a_25891_5238.n0 a_25891_5238.t4 245.386
R8905 a_25891_5238.n1 a_25891_5238.t2 244.766
R8906 a_25891_5238.n0 a_25891_5238.t1 238.716
R8907 a_25891_5238.t0 a_25891_5238.n2 238.716
R8908 a_25891_5238.n1 a_25891_5238.n0 5.07133
R8909 a_25891_5238.n2 a_25891_5238.n1 1.9505
R8910 top_segment_2_0.rseg_2_v3_0.v18.t0 top_segment_2_0.rseg_2_v3_0.v18.n0 238.254
R8911 top_segment_2_0.rseg_2_v3_0.v18.n0 top_segment_2_0.rseg_2_v3_0.v18.t1 10.5761
R8912 top_segment_2_0.rseg_2_v3_0.v18.n0 top_segment_2_0.rseg_2_v3_0.v18.t2 10.5739
R8913 top_segment_2_0.rseg_2_v3_0.v19.t0 top_segment_2_0.rseg_2_v3_0.v19.n0 248.799
R8914 top_segment_2_0.rseg_2_v3_0.v19.n0 top_segment_2_0.rseg_2_v3_0.v19.t1 10.6674
R8915 top_segment_2_0.rseg_2_v3_0.v19.n0 top_segment_2_0.rseg_2_v3_0.v19.t2 10.5285
R8916 a_12878_5238.n0 a_12878_5238.t1 672.461
R8917 a_12878_5238.n1 a_12878_5238.t4 672.087
R8918 a_12878_5238.t0 a_12878_5238.n2 671.755
R8919 a_12878_5238.n1 a_12878_5238.t3 665.667
R8920 a_12878_5238.n0 a_12878_5238.t2 665.667
R8921 a_12878_5238.n2 a_12878_5238.n0 5.39008
R8922 a_12878_5238.n2 a_12878_5238.n1 1.17133
R8923 a_43570_18976.t0 a_43570_18976.t1 49.8467
R8924 top_segment_1_0.rseg_1_v3_1.v57 top_segment_1_0.rseg_1_v3_1.v57.t1 249.345
R8925 top_segment_1_0.rseg_1_v3_1.v57.n0 top_segment_1_0.rseg_1_v3_1.v57.t0 10.575
R8926 top_segment_1_0.rseg_1_v3_1.v57.n0 top_segment_1_0.rseg_1_v3_1.v57.t2 10.5739
R8927 top_segment_1_0.rseg_1_v3_1.v57 top_segment_1_0.rseg_1_v3_1.v57.n0 4.20587
R8928 top_segment_1_0.rseg_1_v3_1.v58 top_segment_1_0.rseg_1_v3_1.v58.t2 249.886
R8929 top_segment_1_0.rseg_1_v3_1.v58.n0 top_segment_1_0.rseg_1_v3_1.v58.t1 10.6247
R8930 top_segment_1_0.rseg_1_v3_1.v58.n0 top_segment_1_0.rseg_1_v3_1.v58.t0 10.5295
R8931 top_segment_1_0.rseg_1_v3_1.v58 top_segment_1_0.rseg_1_v3_1.v58.n0 3.48476
R8932 top_segment_3_0.rseg_3_v3_0.v14.n0 top_segment_3_0.rseg_3_v3_0.v14.t2 678.111
R8933 top_segment_3_0.rseg_3_v3_0.v14.n0 top_segment_3_0.rseg_3_v3_0.v14.t1 10.7803
R8934 top_segment_3_0.rseg_3_v3_0.v14.t0 top_segment_3_0.rseg_3_v3_0.v14.n0 10.7023
R8935 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t0 675.843
R8936 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t1 10.7383
R8937 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.t2 10.6478
R8938 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30.n0 0.682179
R8939 top_segment_1_0.rseg_1_v3_1.v5 top_segment_1_0.rseg_1_v3_1.v5.t0 246.63
R8940 top_segment_1_0.rseg_1_v3_1.v5.n0 top_segment_1_0.rseg_1_v3_1.v5.t2 10.5795
R8941 top_segment_1_0.rseg_1_v3_1.v5.n0 top_segment_1_0.rseg_1_v3_1.v5.t1 10.5739
R8942 top_segment_1_0.rseg_1_v3_1.v5 top_segment_1_0.rseg_1_v3_1.v5.n0 2.90483
R8943 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t1 674.658
R8944 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t0 10.7657
R8945 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t2 10.7357
R8946 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.n0 4.09773
R8947 top_segment_3_0.rseg_3_v3_0.v11.n0 top_segment_3_0.rseg_3_v3_0.v11.t2 677.365
R8948 top_segment_3_0.rseg_3_v3_0.v11.t0 top_segment_3_0.rseg_3_v3_0.v11.n0 10.791
R8949 top_segment_3_0.rseg_3_v3_0.v11.n0 top_segment_3_0.rseg_3_v3_0.v11.t1 10.6292
R8950 a_42271_9350.t0 a_42271_9350.t1 55.3905
R8951 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[2] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t2 753.312
R8952 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n0 268.349
R8953 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t0 268.077
R8954 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.t1 230.518
R8955 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n1 27.3291
R8956 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[2] 12.4649
R8957 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.Y 11.6875
R8958 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n2 7.23528
R8959 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.Y 5.04292
R8960 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.IN.n0 3.68535
R8961 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[2] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[2] 0.90675
R8962 a_42781_7330.t0 a_42781_7330.t1 114.052
R8963 a_41938_3162.t0 a_41938_3162.t1 49.8467
R8964 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t3 241.536
R8965 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n2 195.704
R8966 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t4 169.237
R8967 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n0 152
R8968 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t2 140.53
R8969 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n3 41.8732
R8970 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n1 28.2143
R8971 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t1 26.5955
R8972 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.t0 26.5955
R8973 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 16.5652
R8974 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n4 9.03579
R8975 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 1.87783
R8976 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 1.72748
R8977 a_42781_14894.t0 a_42781_14894.t1 114.052
R8978 a_41714_2426.t0 a_41714_2426.t1 49.8467
R8979 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t3 230.363
R8980 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n2 201.161
R8981 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t4 158.064
R8982 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n3 155.328
R8983 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t1 132.067
R8984 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n4 29.1319
R8985 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t0 26.5955
R8986 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.t2 26.5955
R8987 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n5 23.616
R8988 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n0 4.15748
R8989 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n1 3.76521
R8990 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 3.0725
R8991 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 1.17559
R8992 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.921363
R8993 a_14867_17684.t0 a_14867_17684.n0 671.341
R8994 a_14867_17684.n0 a_14867_17684.t1 666.413
R8995 a_14867_17684.n0 a_14867_17684.t2 665.855
R8996 a_43570_20400.t0 a_43570_20400.t1 49.8467
R8997 a_16279_17684.t0 a_16279_17684.n0 667.216
R8998 a_16279_17684.n0 a_16279_17684.t1 666.692
R8999 a_16279_17684.n0 a_16279_17684.t2 665.433
R9000 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t1 334.822
R9001 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t4 126.27
R9002 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t2 125.558
R9003 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t3 125.558
R9004 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n1 5.73592
R9005 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n2 5.66196
R9006 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n0 0.713
R9007 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t0 0.197295
R9008 a_41787_20650.t0 a_41787_20650.t1 65.941
R9009 a_32733_7938.n0 a_32733_7938.t2 245.316
R9010 a_32733_7938.t0 a_32733_7938.n0 243.361
R9011 a_32733_7938.n0 a_32733_7938.t1 239.308
R9012 a_42781_11290.t0 a_42781_11290.t1 114.052
R9013 a_42245_10734.n0 a_42245_10734.t1 228.04
R9014 a_42245_10734.n0 a_42245_10734.t2 145.648
R9015 a_42245_10734.t0 a_42245_10734.n0 83.2159
R9016 a_23234_19162.n1 a_23234_19162.t1 249.886
R9017 a_23234_19162.n0 a_23234_19162.t3 247.333
R9018 a_23234_19162.n0 a_23234_19162.t2 240.75
R9019 a_23234_19162.t0 a_23234_19162.n1 239.798
R9020 a_23234_19162.n1 a_23234_19162.n0 2.55258
R9021 top_segment_2_0.rseg_2_v3_0.v21.n0 top_segment_2_0.rseg_2_v3_0.v21.t1 239.279
R9022 top_segment_2_0.rseg_2_v3_0.v21.n0 top_segment_2_0.rseg_2_v3_0.v21.t2 10.68
R9023 top_segment_2_0.rseg_2_v3_0.v21.t0 top_segment_2_0.rseg_2_v3_0.v21.n0 10.5763
R9024 a_43570_20124.t0 a_43570_20124.t1 49.8467
R9025 a_13771_17684.t0 a_13771_17684.n0 671.891
R9026 a_13771_17684.n0 a_13771_17684.t1 666.433
R9027 a_13771_17684.n0 a_13771_17684.t2 666.404
R9028 a_21016_17121.n3 a_21016_17121.t3 242.364
R9029 a_21016_17121.n0 a_21016_17121.t2 240.264
R9030 a_21016_17121.n0 a_21016_17121.t1 239.631
R9031 a_21016_17121.n1 a_21016_17121.t4 239.431
R9032 a_21016_17121.n2 a_21016_17121.t5 239.431
R9033 a_21016_17121.t0 a_21016_17121.n3 239.431
R9034 a_21016_17121.n1 a_21016_17121.n0 4.04217
R9035 a_21016_17121.n3 a_21016_17121.n2 2.93383
R9036 a_21016_17121.n2 a_21016_17121.n1 2.93383
R9037 a_22958_19162.n1 a_22958_19162.t1 249.518
R9038 a_22958_19162.n0 a_22958_19162.t3 249.325
R9039 a_22958_19162.n0 a_22958_19162.t2 241.115
R9040 a_22958_19162.t0 a_22958_19162.n1 239.431
R9041 a_22958_19162.n1 a_22958_19162.n0 0.19425
R9042 a_20198_19162.n1 a_20198_19162.t1 251.719
R9043 a_20198_19162.n0 a_20198_19162.t3 248.475
R9044 a_20198_19162.t0 a_20198_19162.n1 241.631
R9045 a_20198_19162.n0 a_20198_19162.t2 238.916
R9046 a_20198_19162.n1 a_20198_19162.n0 3.24425
R9047 top_segment_2_0.rseg_2_v3_0.v47.n0 top_segment_2_0.rseg_2_v3_0.v47.t2 237.56
R9048 top_segment_2_0.rseg_2_v3_0.v47.t0 top_segment_2_0.rseg_2_v3_0.v47.n0 10.5738
R9049 top_segment_2_0.rseg_2_v3_0.v47.n0 top_segment_2_0.rseg_2_v3_0.v47.t1 10.5285
R9050 a_30141_6674.n2 a_30141_6674.t3 246.978
R9051 a_30141_6674.n0 a_30141_6674.t4 244.013
R9052 a_30141_6674.n0 a_30141_6674.t1 240.072
R9053 a_30141_6674.n1 a_30141_6674.t2 239.692
R9054 a_30141_6674.t0 a_30141_6674.n2 239.692
R9055 a_30141_6674.n2 a_30141_6674.n1 6.788
R9056 a_30141_6674.n1 a_30141_6674.n0 2.26092
R9057 a_41529_19966.t0 a_41529_19966.t1 65.941
R9058 a_41787_19966.t0 a_41787_19966.t1 65.941
R9059 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t5 754.659
R9060 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t7 212.081
R9061 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t6 212.081
R9062 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 203.923
R9063 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 186.001
R9064 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t4 139.78
R9065 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t8 139.78
R9066 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 101.49
R9067 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 61.346
R9068 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t1 26.5955
R9069 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t2 26.5955
R9070 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t3 24.9236
R9071 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t0 24.9236
R9072 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 13.5685
R9073 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 10.7525
R9074 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 9.64425
R9075 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 9.30224
R9076 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y 6.6565
R9077 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y 5.04292
R9078 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y 3.8405
R9079 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.A 3.0725
R9080 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y 2.5605
R9081 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 1.93989
R9082 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t4 762.88
R9083 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 203.923
R9084 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 101.49
R9085 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t1 26.5955
R9086 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t0 26.5955
R9087 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t2 24.9236
R9088 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t3 24.9236
R9089 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y 13.0565
R9090 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y 10.7525
R9091 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y 6.6565
R9092 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 5.04292
R9093 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 4.3525
R9094 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 2.5605
R9095 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y 1.93989
R9096 a_34304_9019.n0 a_34304_9019.t1 241.258
R9097 a_34304_9019.t0 a_34304_9019.n0 240.909
R9098 a_34304_9019.n0 a_34304_9019.t2 238.899
R9099 top_segment_1_0.rseg_1_v3_1.v55 top_segment_1_0.rseg_1_v3_1.v55.t2 248.075
R9100 top_segment_1_0.rseg_1_v3_1.v55.n0 top_segment_1_0.rseg_1_v3_1.v55.t0 10.6701
R9101 top_segment_1_0.rseg_1_v3_1.v55.n0 top_segment_1_0.rseg_1_v3_1.v55.t1 10.5739
R9102 top_segment_1_0.rseg_1_v3_1.v55 top_segment_1_0.rseg_1_v3_1.v55.n0 4.16691
R9103 top_segment_1_0.rseg_1_v3_1.v54 top_segment_1_0.rseg_1_v3_1.v54.t2 246.798
R9104 top_segment_1_0.rseg_1_v3_1.v54.n0 top_segment_1_0.rseg_1_v3_1.v54.t1 10.6247
R9105 top_segment_1_0.rseg_1_v3_1.v54.n0 top_segment_1_0.rseg_1_v3_1.v54.t0 10.5295
R9106 top_segment_1_0.rseg_1_v3_1.v54 top_segment_1_0.rseg_1_v3_1.v54.n0 3.49191
R9107 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t2 158.273
R9108 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t0 141.358
R9109 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t3 140.304
R9110 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t1 139.566
R9111 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n0 8.02027
R9112 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n1 0.063
R9113 top_segment_2_0.rseg_2_v3_0.v20.n0 top_segment_2_0.rseg_2_v3_0.v20.t1 239.094
R9114 top_segment_2_0.rseg_2_v3_0.v20.t0 top_segment_2_0.rseg_2_v3_0.v20.n0 10.6701
R9115 top_segment_2_0.rseg_2_v3_0.v20.n0 top_segment_2_0.rseg_2_v3_0.v20.t2 10.5739
R9116 a_42245_12714.t0 a_42245_12714.n0 228.04
R9117 a_42245_12714.n0 a_42245_12714.t2 145.648
R9118 a_42245_12714.n0 a_42245_12714.t1 83.2159
R9119 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t1 227.856
R9120 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n2 152.333
R9121 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t2 140.382
R9122 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t3 114.031
R9123 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t0 83.3993
R9124 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.t4 81.5883
R9125 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n3 14.4422
R9126 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/buff_hvl_0.IN top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n1 7.56882
R9127 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n0 5.08175
R9128 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.OUTP.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.A 0.831669
R9129 a_42271_12874.t0 a_42271_12874.t1 55.3905
R9130 a_43570_19252.t0 a_43570_19252.t1 49.8467
R9131 a_42781_11924.t0 a_42781_11924.t1 114.052
R9132 a_41714_3622.t0 a_41714_3622.t1 49.8467
R9133 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t2 673.212
R9134 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t1 10.7631
R9135 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t0 10.7147
R9136 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.n0 2.72674
R9137 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t1 673.273
R9138 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t2 10.7798
R9139 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.t0 10.6302
R9140 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6.n0 3.43753
R9141 top_segment_3_0.rseg_3_v3_0.v6.t0 top_segment_3_0.rseg_3_v3_0.v6.n0 679.191
R9142 top_segment_3_0.rseg_3_v3_0.v6.n0 top_segment_3_0.rseg_3_v3_0.v6.t1 10.7575
R9143 top_segment_3_0.rseg_3_v3_0.v6.n0 top_segment_3_0.rseg_3_v3_0.v6.t2 10.7275
R9144 top_segment_3_0.rseg_3_v3_0.v7.t0 top_segment_3_0.rseg_3_v3_0.v7.n0 680.072
R9145 top_segment_3_0.rseg_3_v3_0.v7.n0 top_segment_3_0.rseg_3_v3_0.v7.t2 10.7276
R9146 top_segment_3_0.rseg_3_v3_0.v7.n0 top_segment_3_0.rseg_3_v3_0.v7.t1 10.6922
R9147 top_segment_4_1.b0.n2 top_segment_4_1.b0.n1 863.124
R9148 top_segment_4_1.b0.n1 top_segment_4_1.b0.n0 585
R9149 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y top_segment_4_1.b0.t1 495.469
R9150 top_segment_4_1.b0.t0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 291.983
R9151 top_segment_4_1.b0.n6 top_segment_4_1.b0.t0 285
R9152 top_segment_4_1.b0.n4 top_segment_4_1.b0.t3 254.05
R9153 top_segment_4_1.b0.n3 top_segment_4_1.b0.t2 208.054
R9154 top_segment_4_1.b0.n1 top_segment_4_1.b0.t1 140.738
R9155 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.b[0] top_segment_4_1.b0.n4 29.688
R9156 top_segment_4_1.b0.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUT 14.3755
R9157 top_segment_4_1.b0.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 12.4126
R9158 top_segment_4_1.b0.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 11.6369
R9159 top_segment_4_1.b0.n4 top_segment_4_1.b0.n3 10.8443
R9160 top_segment_4_1.b0.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 10.1408
R9161 top_segment_4_1.b0.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 8.53383
R9162 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y top_segment_4_1.b0.n5 5.81868
R9163 top_segment_4_1.b0.n3 top_segment_1_0.b[0] 4.71204
R9164 top_segment_4_1.b0.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y 2.16154
R9165 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y top_segment_4_1.b0.n6 1.93989
R9166 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y top_segment_4_1.b0.n2 0.665435
R9167 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUT top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.b[0] 0.19425
R9168 top_segment_3_0.rseg_3_v3_0.v8.t0 top_segment_3_0.rseg_3_v3_0.v8.n1 676.072
R9169 top_segment_3_0.rseg_3_v3_0.v8.n1 top_segment_3_0.rseg_3_v3_0.v8.t3 672.926
R9170 top_segment_3_0.rseg_3_v3_0.v8.n0 top_segment_3_0.rseg_3_v3_0.v8.t1 13.884
R9171 top_segment_3_0.rseg_3_v3_0.v8.n0 top_segment_3_0.rseg_3_v3_0.v8.t2 10.7934
R9172 top_segment_3_0.rseg_3_v3_0.v8.n1 top_segment_3_0.rseg_3_v3_0.v8.n0 5.03253
R9173 a_41271_18542.t0 a_41271_18542.t1 65.941
R9174 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t3 230.363
R9175 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n0 203.147
R9176 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t4 158.064
R9177 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n1 152
R9178 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t2 140.53
R9179 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n3 34.4304
R9180 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t1 26.5955
R9181 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.t0 26.5955
R9182 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n2 24.0657
R9183 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 16.5652
R9184 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n4 9.03579
R9185 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 3.2005
R9186 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 1.72748
R9187 top_segment_1_0.rseg_1_v3_1.v3 top_segment_1_0.rseg_1_v3_1.v3.t2 245.726
R9188 top_segment_1_0.rseg_1_v3_1.v3.n0 top_segment_1_0.rseg_1_v3_1.v3.t0 10.5816
R9189 top_segment_1_0.rseg_1_v3_1.v3.n0 top_segment_1_0.rseg_1_v3_1.v3.t1 10.5739
R9190 top_segment_1_0.rseg_1_v3_1.v3 top_segment_1_0.rseg_1_v3_1.v3.n0 1.48638
R9191 top_segment_3_0.V0.n1 top_segment_3_0.V0.t0 668.619
R9192 top_segment_3_0.V0.n0 top_segment_3_0.V0.t3 238.077
R9193 top_segment_3_0.V0.n1 top_segment_3_0.V0.t2 12.4069
R9194 top_segment_3_0.V0.n0 top_segment_3_0.V0.t1 10.6569
R9195 top_segment_2_0.V48 top_segment_3_0.V0.n0 1.29821
R9196 top_segment_2_0.V48 top_segment_3_0.V0.n1 0.397447
R9197 top_segment_2_0.DEC1[2].n4 top_segment_2_0.DEC1[2].t1 334.788
R9198 top_segment_2_0.DEC1[2].n1 top_segment_2_0.DEC1[2].t9 213.218
R9199 top_segment_2_0.DEC1[2] top_segment_2_0.DEC1[2].t6 212.982
R9200 top_segment_2_0.DEC1[2].n1 top_segment_2_0.DEC1[2].t2 212.554
R9201 top_segment_2_0.DEC1[2].n0 top_segment_2_0.DEC1[2].t4 212.554
R9202 top_segment_2_0.DEC1[2].n3 top_segment_2_0.DEC1[2].t7 208.054
R9203 top_segment_2_0.DEC1[2].n6 top_segment_2_0.DEC1[2].t8 126.27
R9204 top_segment_2_0.DEC1[2].n6 top_segment_2_0.DEC1[2].t3 125.558
R9205 top_segment_2_0.DEC1[2].n5 top_segment_2_0.DEC1[2].t5 121.127
R9206 top_segment_2_0.DEC1[2].n4 top_segment_2_0.DEC1[2].t0 87.8063
R9207 top_segment_2_0.DEC1[2] top_segment_2_0.DEC1[2].n3 60.0689
R9208 top_segment_2_0.DEC1[2].n7 top_segment_2_0.DEC1[2].n6 5.73592
R9209 top_segment_2_0.DEC1[2] top_segment_2_0.DEC1[2].n7 5.388
R9210 top_segment_2_0.DEC1[2].n3 top_segment_2_0.DEC1[2].n2 4.5005
R9211 top_segment_2_0.DEC1[2].n2 top_segment_2_0.DEC1[2].n0 0.663962
R9212 top_segment_2_0.DEC1[2].n2 top_segment_2_0.DEC1[2].n1 0.663962
R9213 top_segment_2_0.DEC1[2].n5 top_segment_2_0.DEC1[2].n4 0.322615
R9214 top_segment_2_0.DEC1[2].n0 top_segment_2_0.DEC1[2] 0.236077
R9215 top_segment_2_0.DEC1[2].n7 top_segment_2_0.DEC1[2].n5 0.177583
R9216 top_segment_1_0.rseg_1_v3_1.v44 top_segment_1_0.rseg_1_v3_1.v44.t0 249.209
R9217 top_segment_1_0.rseg_1_v3_1.v44.n0 top_segment_1_0.rseg_1_v3_1.v44.t1 10.5296
R9218 top_segment_1_0.rseg_1_v3_1.v44.n0 top_segment_1_0.rseg_1_v3_1.v44.t2 10.5285
R9219 top_segment_1_0.rseg_1_v3_1.v44 top_segment_1_0.rseg_1_v3_1.v44.n0 2.13671
R9220 a_42609_18861.t0 a_42609_18861.t1 129.28
R9221 a_42271_13310.t0 a_42271_13310.t1 55.3905
R9222 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t0 676.712
R9223 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t1 10.7718
R9224 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t2 10.6268
R9225 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.n0 3.43316
R9226 top_segment_1_0.rseg_1_v3_1.v16.t0 top_segment_1_0.rseg_1_v3_1.v16.n0 241.547
R9227 top_segment_1_0.rseg_1_v3_1.v16.n0 top_segment_1_0.rseg_1_v3_1.v16.t1 12.2056
R9228 top_segment_1_0.rseg_1_v3_1.v16.n0 top_segment_1_0.rseg_1_v3_1.v16.t2 12.0758
R9229 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[2] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t7 752.615
R9230 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n5 258.363
R9231 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t6 230.576
R9232 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n4 202.094
R9233 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t5 158.275
R9234 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n0 152
R9235 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t2 126.469
R9236 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n6 62.4946
R9237 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t1 32.5055
R9238 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t0 32.5055
R9239 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t3 26.5955
R9240 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.t4 26.5955
R9241 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[2] 13.6567
R9242 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n1 12.0102
R9243 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n2 9.82192
R9244 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_3.A 6.66717
R9245 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n3 6.51278
R9246 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/lvsf_0.INB.n7 4.04261
R9247 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[2] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[2] 0.853179
R9248 a_12602_5238.n0 a_12602_5238.t1 672.278
R9249 a_12602_5238.n1 a_12602_5238.t4 671.904
R9250 a_12602_5238.t0 a_12602_5238.n2 671.547
R9251 a_12602_5238.n1 a_12602_5238.t3 665.484
R9252 a_12602_5238.n0 a_12602_5238.t2 665.484
R9253 a_12602_5238.n2 a_12602_5238.n0 4.99842
R9254 a_12602_5238.n2 a_12602_5238.n1 1.563
R9255 top_segment_2_0.rseg_2_v3_0.v17.t0 top_segment_2_0.rseg_2_v3_0.v17.n0 242.349
R9256 top_segment_2_0.rseg_2_v3_0.v17.n0 top_segment_2_0.rseg_2_v3_0.v17.t2 10.6919
R9257 top_segment_2_0.rseg_2_v3_0.v17.n0 top_segment_2_0.rseg_2_v3_0.v17.t1 10.5285
R9258 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t1 675.904
R9259 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t0 10.7766
R9260 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.t2 10.6951
R9261 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45.n0 1.35956
R9262 top_segment_1_0.rseg_1_v3_1.v51 top_segment_1_0.rseg_1_v3_1.v51.t2 245.726
R9263 top_segment_1_0.rseg_1_v3_1.v51.n0 top_segment_1_0.rseg_1_v3_1.v51.t0 10.575
R9264 top_segment_1_0.rseg_1_v3_1.v51.n0 top_segment_1_0.rseg_1_v3_1.v51.t1 10.5739
R9265 top_segment_1_0.rseg_1_v3_1.v51 top_segment_1_0.rseg_1_v3_1.v51.n0 1.5626
R9266 a_41271_19966.t0 a_41271_19966.t1 65.941
R9267 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t2 676.321
R9268 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t1 13.4532
R9269 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t0 10.7781
R9270 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.n0 4.72836
R9271 a_43026_2242.t0 a_43026_2242.t1 49.8467
R9272 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t2 672.722
R9273 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t1 10.7152
R9274 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.t0 10.6722
R9275 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20.n0 2.05317
R9276 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t3 593.396
R9277 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 231.554
R9278 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t1 140.53
R9279 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t0 26.5955
R9280 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.t2 26.5955
R9281 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 16.5652
R9282 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 9.03579
R9283 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n1 6.02403
R9284 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 1.72748
R9285 a_42609_17793.t0 a_42609_17793.t1 129.28
R9286 a_42609_17437.t0 a_42609_17437.t1 129.28
R9287 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.n0 663.232
R9288 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t1 10.6713
R9289 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v33.t2 10.5739
R9290 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.n0 668.13
R9291 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t1 12.1392
R9292 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v32.t2 12.0758
R9293 a_41529_18884.t0 a_41529_18884.t1 65.941
R9294 a_41787_18884.t0 a_41787_18884.t1 65.941
R9295 a_14728_6674.n0 a_14728_6674.t3 672.213
R9296 a_14728_6674.t0 a_14728_6674.n2 668.944
R9297 a_14728_6674.n2 a_14728_6674.t4 666.405
R9298 a_14728_6674.n0 a_14728_6674.t2 665.726
R9299 a_14728_6674.n1 a_14728_6674.t1 665.726
R9300 a_14728_6674.n1 a_14728_6674.n0 6.63383
R9301 a_14728_6674.n2 a_14728_6674.n1 3.73592
R9302 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t2 675.533
R9303 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t1 10.7625
R9304 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.t0 10.7161
R9305 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11.n0 2.72817
R9306 a_19370_19162.n2 a_19370_19162.t3 251.168
R9307 a_19370_19162.n0 a_19370_19162.t1 250.329
R9308 a_19370_19162.t0 a_19370_19162.n2 241.082
R9309 a_19370_19162.n1 a_19370_19162.t2 239.465
R9310 a_19370_19162.n0 a_19370_19162.t4 239.465
R9311 a_19370_19162.n1 a_19370_19162.n0 0.633833
R9312 a_19370_19162.n2 a_19370_19162.n1 0.20675
R9313 top_segment_2_0.rseg_2_v3_0.v32.t0 top_segment_2_0.rseg_2_v3_0.v32.n1 237.611
R9314 top_segment_2_0.rseg_2_v3_0.v32.n0 top_segment_2_0.rseg_2_v3_0.v32.t3 237.554
R9315 top_segment_2_0.rseg_2_v3_0.v32.n1 top_segment_2_0.rseg_2_v3_0.v32.t2 10.6569
R9316 top_segment_2_0.rseg_2_v3_0.v32.n0 top_segment_2_0.rseg_2_v3_0.v32.t1 10.6569
R9317 top_segment_2_0.rseg_2_v3_0.v32.n1 top_segment_2_0.rseg_2_v3_0.v32.n0 3.36262
R9318 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t2 675.533
R9319 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t1 10.7636
R9320 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.t0 10.7261
R9321 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59.n0 2.74248
R9322 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t1 677.236
R9323 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t2 10.7534
R9324 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t0 10.6226
R9325 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.n0 3.42573
R9326 top_segment_3_0.rseg_3_v3_0.v1.t0 top_segment_3_0.rseg_3_v3_0.v1.n0 663.775
R9327 top_segment_3_0.rseg_3_v3_0.v1.n0 top_segment_3_0.rseg_3_v3_0.v1.t1 10.6247
R9328 top_segment_3_0.rseg_3_v3_0.v1.n0 top_segment_3_0.rseg_3_v3_0.v1.t2 10.5285
R9329 a_15419_17684.t0 a_15419_17684.n0 670.976
R9330 a_15419_17684.n0 a_15419_17684.t1 666.78
R9331 a_15419_17684.n0 a_15419_17684.t2 665.487
R9332 VL3 VL3.t0 666.389
R9333 VL3.n0 VL3.t1 665.244
R9334 VL3.n0 VL3 0.063
R9335 VL3 VL3.n0 0.013
R9336 a_20750_19162.n1 a_20750_19162.t1 250.986
R9337 a_20750_19162.n0 a_20750_19162.t2 249.524
R9338 a_20750_19162.t0 a_20750_19162.n1 240.898
R9339 a_20750_19162.n0 a_20750_19162.t3 239.649
R9340 a_20750_19162.n1 a_20750_19162.n0 1.46092
R9341 a_41271_17460.t0 a_41271_17460.t1 65.941
R9342 a_17547_7938.n0 a_17547_7938.t1 670.336
R9343 a_17547_7938.n0 a_17547_7938.t2 670
R9344 a_17547_7938.t0 a_17547_7938.n0 666.258
R9345 a_42781_15250.t0 a_42781_15250.t1 114.052
R9346 top_segment_1_0.rseg_1_v3_1.v40 top_segment_1_0.rseg_1_v3_1.v40.t2 249.738
R9347 top_segment_1_0.rseg_1_v3_1.v40.n0 top_segment_1_0.rseg_1_v3_1.v40.t0 13.4756
R9348 top_segment_1_0.rseg_1_v3_1.v40.n0 top_segment_1_0.rseg_1_v3_1.v40.t1 10.7876
R9349 top_segment_1_0.rseg_1_v3_1.v40 top_segment_1_0.rseg_1_v3_1.v40.n0 4.72836
R9350 top_segment_2_0.rseg_2_v3_0.v38.n0 top_segment_2_0.rseg_2_v3_0.v38.t2 239.793
R9351 top_segment_2_0.rseg_2_v3_0.v38.t0 top_segment_2_0.rseg_2_v3_0.v38.n0 10.7638
R9352 top_segment_2_0.rseg_2_v3_0.v38.n0 top_segment_2_0.rseg_2_v3_0.v38.t1 10.7314
R9353 a_42781_6340.t0 a_42781_6340.t1 114.052
R9354 a_42245_5784.t0 a_42245_5784.n0 228.04
R9355 a_42245_5784.n0 a_42245_5784.t2 145.648
R9356 a_42245_5784.n0 a_42245_5784.t1 83.2159
R9357 top_segment_2_0.rseg_2_v3_0.v3.n0 top_segment_2_0.rseg_2_v3_0.v3.t1 241.31
R9358 top_segment_2_0.rseg_2_v3_0.v3.n0 top_segment_2_0.rseg_2_v3_0.v3.t2 10.5439
R9359 top_segment_2_0.rseg_2_v3_0.v3.t0 top_segment_2_0.rseg_2_v3_0.v3.n0 10.5295
R9360 a_37219_19465.t0 a_37219_19465.n0 233.361
R9361 a_37219_19465.n0 a_37219_19465.t2 229.339
R9362 a_37219_19465.n0 a_37219_19465.t1 227.399
R9363 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t1 668.13
R9364 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.n0 12.1235
R9365 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v16.t2 12.0758
R9366 a_42609_20285.t0 a_42609_20285.t1 129.28
R9367 a_41271_18884.t0 a_41271_18884.t1 65.941
R9368 a_32457_7938.n0 a_32457_7938.t2 244.909
R9369 a_32457_7938.t0 a_32457_7938.n0 243.178
R9370 a_32457_7938.n0 a_32457_7938.t1 239.489
R9371 a_21578_19162.n1 a_21578_19162.t3 250.069
R9372 a_21578_19162.n0 a_21578_19162.t2 249.745
R9373 a_21578_19162.n0 a_21578_19162.t1 240.565
R9374 a_21578_19162.t0 a_21578_19162.n1 239.982
R9375 a_21578_19162.n1 a_21578_19162.n0 0.323417
R9376 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t2 673.192
R9377 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t0 10.7578
R9378 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.t1 10.6535
R9379 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2.n0 0.67884
R9380 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.t0 10.7652
R9381 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.t1 10.6927
R9382 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61.n0 1.36672
R9383 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.n0 676.833
R9384 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t2 10.7929
R9385 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v62.t1 10.5285
R9386 a_43026_3158.t0 a_43026_3158.t1 49.8467
R9387 a_43026_3242.t0 a_43026_3242.t1 60.9236
R9388 a_42802_3518.t0 a_42802_3518.t1 49.8467
R9389 a_42802_3602.t0 a_42802_3602.t1 60.9236
R9390 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t2 672.309
R9391 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t1 10.791
R9392 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.t0 10.6937
R9393 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3.n0 1.35575
R9394 top_segment_3_0.rseg_3_v3_0.v3.t0 top_segment_3_0.rseg_3_v3_0.v3.n0 674.707
R9395 top_segment_3_0.rseg_3_v3_0.v3.n0 top_segment_3_0.rseg_3_v3_0.v3.t1 10.7549
R9396 top_segment_3_0.rseg_3_v3_0.v3.n0 top_segment_3_0.rseg_3_v3_0.v3.t2 10.6512
R9397 a_37853_19465.n0 a_37853_19465.t2 239.25
R9398 a_37853_19465.n0 a_37853_19465.t0 222.119
R9399 a_37853_19465.t1 a_37853_19465.n0 222.119
R9400 a_33127_7938.n0 a_33127_7938.t2 245.95
R9401 a_33127_7938.n0 a_33127_7938.t1 244.102
R9402 a_33127_7938.t0 a_33127_7938.n0 238.94
R9403 a_42781_6974.t0 a_42781_6974.t1 114.052
R9404 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t1 675.929
R9405 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t0 10.7912
R9406 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t2 10.6717
R9407 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.n0 4.09783
R9408 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t1 672.309
R9409 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t2 10.7751
R9410 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.t0 10.6965
R9411 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35.n0 1.35813
R9412 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t1 673.332
R9413 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t0 10.7393
R9414 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.t2 10.6478
R9415 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34.n0 0.682179
R9416 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 272.038
R9417 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t1 258.846
R9418 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t3 230.363
R9419 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n5 224.775
R9420 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t4 158.064
R9421 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n0 153.28
R9422 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t0 26.5955
R9423 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.t2 26.5955
R9424 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n1 19.4367
R9425 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 5.1205
R9426 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n4 3.76521
R9427 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n3 3.03935
R9428 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n2 1.56597
R9429 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.921363
R9430 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B.n2 0.737191
R9431 a_43570_17276.t0 a_43570_17276.t1 49.8467
R9432 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t3 743.342
R9433 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n7 586.745
R9434 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n6 289.24
R9435 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t5 230.576
R9436 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t4 158.275
R9437 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n2 152
R9438 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n0 94.1864
R9439 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n5 82.6525
R9440 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t1 26.5955
R9441 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t0 24.9236
R9442 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.t2 24.9236
R9443 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n5 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n4 21.3341
R9444 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n6 17.9639
R9445 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n3 9.3005
R9446 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_1.A 6.66717
R9447 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[1] 3.48572
R9448 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[1] 0.790679
R9449 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[1] 0.063
R9450 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.INB.n1 0.063
R9451 a_41394_3894.t0 a_41394_3894.t1 41.3705
R9452 top_segment_1_0.rseg_1_v3_1.v11 top_segment_1_0.rseg_1_v3_1.v11.t2 248.95
R9453 top_segment_1_0.rseg_1_v3_1.v11.n0 top_segment_1_0.rseg_1_v3_1.v11.t0 10.5761
R9454 top_segment_1_0.rseg_1_v3_1.v11.n0 top_segment_1_0.rseg_1_v3_1.v11.t1 10.5739
R9455 top_segment_1_0.rseg_1_v3_1.v11 top_segment_1_0.rseg_1_v3_1.v11.n0 2.84608
R9456 top_segment_1_0.rseg_1_v3_1.v12 top_segment_1_0.rseg_1_v3_1.v12.t2 249.594
R9457 top_segment_1_0.rseg_1_v3_1.v12.n0 top_segment_1_0.rseg_1_v3_1.v12.t1 10.5307
R9458 top_segment_1_0.rseg_1_v3_1.v12.n0 top_segment_1_0.rseg_1_v3_1.v12.t0 10.5295
R9459 top_segment_1_0.rseg_1_v3_1.v12 top_segment_1_0.rseg_1_v3_1.v12.n0 2.17402
R9460 a_12326_5238.n0 a_12326_5238.t1 672.093
R9461 a_12326_5238.n1 a_12326_5238.t4 671.721
R9462 a_12326_5238.t0 a_12326_5238.n2 671.35
R9463 a_12326_5238.n1 a_12326_5238.t3 665.299
R9464 a_12326_5238.n0 a_12326_5238.t2 665.299
R9465 a_12326_5238.n2 a_12326_5238.n0 4.60675
R9466 a_12326_5238.n2 a_12326_5238.n1 1.95467
R9467 a_41394_2698.t0 a_41394_2698.t1 41.3705
R9468 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[4] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t2 752.994
R9469 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t0 230.517
R9470 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t1 162.351
R9471 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[4] 26.8833
R9472 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y 11.6875
R9473 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y 7.23528
R9474 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 3.10353
R9475 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 1.93989
R9476 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[4] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[4] 0.790679
R9477 SH[1].n2 SH[1].n1 863.124
R9478 SH[1].n1 SH[1].n0 585
R9479 SH[1] SH[1].t1 495.469
R9480 SH[1].n3 SH[1].t0 141.189
R9481 SH[1].n1 SH[1].t1 140.738
R9482 SH[1] SH[1].n4 14.5776
R9483 SH[1].n2 SH[1] 11.6369
R9484 SH[1].n0 SH[1] 10.1408
R9485 SH[1].n4 SH[1] 8.14595
R9486 SH[1] SH[1].n3 7.94225
R9487 SH[1].n4 SH[1] 6.20656
R9488 SH[1].n3 SH[1] 6.14988
R9489 SH[1].n0 SH[1] 2.16154
R9490 SH[1] SH[1].n2 0.665435
R9491 a_42802_3434.t0 a_42802_3434.t1 49.8467
R9492 VS1 VS1.t0 239.155
R9493 VS1.n0 VS1.t1 238.716
R9494 VS1 VS1.n0 0.196333
R9495 VS1.n0 VS1 0.063
R9496 top_segment_1_0.rseg_1_v3_1.v15.n0 top_segment_1_0.rseg_1_v3_1.v15.t2 240.469
R9497 top_segment_1_0.rseg_1_v3_1.v15.t0 top_segment_1_0.rseg_1_v3_1.v15.n0 10.6713
R9498 top_segment_1_0.rseg_1_v3_1.v15.n0 top_segment_1_0.rseg_1_v3_1.v15.t1 10.5739
R9499 a_30417_6674.n2 a_30417_6674.t3 247.161
R9500 a_30417_6674.n0 a_30417_6674.t4 244.589
R9501 a_30417_6674.n0 a_30417_6674.t1 240.337
R9502 a_30417_6674.n1 a_30417_6674.t2 239.875
R9503 a_30417_6674.t0 a_30417_6674.n2 239.875
R9504 a_30417_6674.n2 a_30417_6674.n1 6.788
R9505 a_30417_6674.n1 a_30417_6674.n0 1.86925
R9506 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.n0 667.057
R9507 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t2 10.6819
R9508 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v47.t1 10.5739
R9509 top_segment_2_0.rseg_2_v3_0.v37.n0 top_segment_2_0.rseg_2_v3_0.v37.t2 239.32
R9510 top_segment_2_0.rseg_2_v3_0.v37.n0 top_segment_2_0.rseg_2_v3_0.v37.t1 10.716
R9511 top_segment_2_0.rseg_2_v3_0.v37.t0 top_segment_2_0.rseg_2_v3_0.v37.n0 10.6708
R9512 a_42609_18505.t0 a_42609_18505.t1 129.28
R9513 a_43570_17552.t0 a_43570_17552.t1 49.8467
R9514 top_segment_1_0.rseg_1_v3_1.v37 top_segment_1_0.rseg_1_v3_1.v37.t2 246.63
R9515 top_segment_1_0.rseg_1_v3_1.v37.n0 top_segment_1_0.rseg_1_v3_1.v37.t0 10.575
R9516 top_segment_1_0.rseg_1_v3_1.v37.n0 top_segment_1_0.rseg_1_v3_1.v37.t1 10.5739
R9517 top_segment_1_0.rseg_1_v3_1.v37 top_segment_1_0.rseg_1_v3_1.v37.n0 2.81913
R9518 a_42271_6380.t0 a_42271_6380.t1 55.3905
R9519 top_segment_2_0.rseg_2_v3_0.v27.t0 top_segment_2_0.rseg_2_v3_0.v27.n0 239.248
R9520 top_segment_2_0.rseg_2_v3_0.v27.n0 top_segment_2_0.rseg_2_v3_0.v27.t2 10.7181
R9521 top_segment_2_0.rseg_2_v3_0.v27.n0 top_segment_2_0.rseg_2_v3_0.v27.t1 10.6712
R9522 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t1 676.48
R9523 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t2 10.7826
R9524 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t0 10.6326
R9525 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.n0 3.43753
R9526 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t2 676.497
R9527 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t0 10.7173
R9528 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t1 10.675
R9529 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.n0 2.06176
R9530 a_41271_20650.t0 a_41271_20650.t1 65.941
R9531 SH[3].n2 SH[3].n1 863.124
R9532 SH[3].n1 SH[3].n0 585
R9533 SH[3] SH[3].t1 495.469
R9534 SH[3].n3 SH[3].t0 141.189
R9535 SH[3].n1 SH[3].t1 140.738
R9536 SH[3] SH[3].n4 14.5776
R9537 SH[3].n2 SH[3] 11.6369
R9538 SH[3].n0 SH[3] 10.1408
R9539 SH[3].n4 SH[3] 8.14595
R9540 SH[3] SH[3].n3 7.94225
R9541 SH[3].n4 SH[3] 6.20656
R9542 SH[3].n3 SH[3] 6.14988
R9543 SH[3].n0 SH[3] 2.16154
R9544 SH[3] SH[3].n2 0.665435
R9545 top_segment_1_0.rseg_1_v3_1.v30 top_segment_1_0.rseg_1_v3_1.v30.t0 249.358
R9546 top_segment_1_0.rseg_1_v3_1.v30.n0 top_segment_1_0.rseg_1_v3_1.v30.t1 10.5296
R9547 top_segment_1_0.rseg_1_v3_1.v30.n0 top_segment_1_0.rseg_1_v3_1.v30.t2 10.5285
R9548 top_segment_1_0.rseg_1_v3_1.v30 top_segment_1_0.rseg_1_v3_1.v30.n0 0.905521
R9549 top_segment_1_0.rseg_1_v3_1.v62 top_segment_1_0.rseg_1_v3_1.v62.t2 249.178
R9550 top_segment_1_0.rseg_1_v3_1.v62.n0 top_segment_1_0.rseg_1_v3_1.v62.t0 10.6257
R9551 top_segment_1_0.rseg_1_v3_1.v62.n0 top_segment_1_0.rseg_1_v3_1.v62.t1 10.5285
R9552 top_segment_1_0.rseg_1_v3_1.v62 top_segment_1_0.rseg_1_v3_1.v62.n0 0.872789
R9553 a_42271_8914.t0 a_42271_8914.t1 55.3905
R9554 a_42802_3066.t0 a_42802_3066.t1 49.8467
R9555 a_42802_3150.t0 a_42802_3150.t1 60.9236
R9556 top_segment_2_0.rseg_2_v3_0.v15.n0 top_segment_2_0.rseg_2_v3_0.v15.t1 237.542
R9557 top_segment_2_0.rseg_2_v3_0.v15.t0 top_segment_2_0.rseg_2_v3_0.v15.n0 10.5334
R9558 top_segment_2_0.rseg_2_v3_0.v15.n0 top_segment_2_0.rseg_2_v3_0.v15.t2 10.5312
R9559 a_22756_17121.n0 a_22756_17121.t1 241.857
R9560 a_22756_17121.n2 a_22756_17121.t2 241.815
R9561 a_22756_17121.n0 a_22756_17121.t3 238.881
R9562 a_22756_17121.n1 a_22756_17121.t4 238.881
R9563 a_22756_17121.t0 a_22756_17121.n2 238.881
R9564 a_22756_17121.n2 a_22756_17121.n1 2.93383
R9565 a_22756_17121.n1 a_22756_17121.n0 2.93383
R9566 a_21302_19162.n2 a_21302_19162.t2 250.435
R9567 a_21302_19162.n0 a_21302_19162.t3 249.549
R9568 a_21302_19162.t0 a_21302_19162.n2 240.347
R9569 a_21302_19162.n0 a_21302_19162.t4 240.2
R9570 a_21302_19162.n1 a_21302_19162.t1 240.2
R9571 a_21302_19162.n1 a_21302_19162.n0 0.633833
R9572 a_21302_19162.n2 a_21302_19162.n1 0.252583
R9573 a_42781_8954.t0 a_42781_8954.t1 114.052
R9574 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.n0 667.052
R9575 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t2 10.6713
R9576 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v31.t1 10.5739
R9577 top_segment_2_0.rseg_2_v3_0.v14.n0 top_segment_2_0.rseg_2_v3_0.v14.t1 238.232
R9578 top_segment_2_0.rseg_2_v3_0.v14.n0 top_segment_2_0.rseg_2_v3_0.v14.t2 10.5771
R9579 top_segment_2_0.rseg_2_v3_0.v14.t0 top_segment_2_0.rseg_2_v3_0.v14.n0 10.5739
R9580 a_14176_6674.n0 a_14176_6674.t3 671.846
R9581 a_14176_6674.t0 a_14176_6674.n2 667.794
R9582 a_14176_6674.n2 a_14176_6674.t4 667.572
R9583 a_14176_6674.n0 a_14176_6674.t2 665.36
R9584 a_14176_6674.n1 a_14176_6674.t1 665.36
R9585 a_14176_6674.n1 a_14176_6674.n0 6.63383
R9586 a_14176_6674.n2 a_14176_6674.n1 4.51925
R9587 a_41938_2782.t0 a_41938_2782.t1 49.8467
R9588 a_41938_2866.t0 a_41938_2866.t1 60.9236
R9589 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t1 668.13
R9590 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.n0 12.177
R9591 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v48.t2 12.0758
R9592 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t2 672.655
R9593 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t0 10.7134
R9594 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.t1 10.6712
R9595 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4.n0 2.05317
R9596 top_segment_2_0.rseg_2_v3_0.v28.t0 top_segment_2_0.rseg_2_v3_0.v28.n0 238.876
R9597 top_segment_2_0.rseg_2_v3_0.v28.n0 top_segment_2_0.rseg_2_v3_0.v28.t2 10.7601
R9598 top_segment_2_0.rseg_2_v3_0.v28.n0 top_segment_2_0.rseg_2_v3_0.v28.t1 10.719
R9599 a_41529_20992.t0 a_41529_20992.t1 65.941
R9600 a_41787_20992.t0 a_41787_20992.t1 65.941
R9601 a_42271_10340.t0 a_42271_10340.t1 55.3905
R9602 a_42245_9744.n0 a_42245_9744.t1 228.04
R9603 a_42245_9744.n0 a_42245_9744.t2 145.648
R9604 a_42245_9744.t0 a_42245_9744.n0 83.2159
R9605 a_43890_2882.t0 a_43890_2882.t1 49.8467
R9606 a_43890_2966.t0 a_43890_2966.t1 60.9236
R9607 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t1 274.793
R9608 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t5 231.017
R9609 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n3 205.28
R9610 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t4 158.716
R9611 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n0 153.347
R9612 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t2 130.49
R9613 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n4 67.4857
R9614 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n2 38.9629
R9615 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t3 26.5955
R9616 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.t0 26.5955
R9617 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n1 22.1046
R9618 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 3.81804
R9619 DIN2.n1 DIN2.t1 212.081
R9620 DIN2.n0 DIN2.t0 212.081
R9621 DIN2.n2 DIN2.n1 183.185
R9622 DIN2.n1 DIN2.t3 139.78
R9623 DIN2.n0 DIN2.t2 139.78
R9624 DIN2.n1 DIN2.n0 61.346
R9625 DIN2 DIN2.n2 14.2776
R9626 DIN2.n2 DIN2 5.8885
R9627 a_42781_8320.t0 a_42781_8320.t1 114.052
R9628 a_42781_15884.t0 a_42781_15884.t1 114.052
R9629 DIN5.n1 DIN5.t1 212.081
R9630 DIN5.n0 DIN5.t0 212.081
R9631 DIN5.n2 DIN5.n1 183.185
R9632 DIN5.n1 DIN5.t3 139.78
R9633 DIN5.n0 DIN5.t2 139.78
R9634 DIN5.n1 DIN5.n0 61.346
R9635 DIN5 DIN5.n2 14.2776
R9636 DIN5.n2 DIN5 5.8885
R9637 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t3 593.158
R9638 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 231.554
R9639 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t2 140.53
R9640 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t1 26.5955
R9641 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.t0 26.5955
R9642 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 16.5652
R9643 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 9.03579
R9644 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n1 6.02403
R9645 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y.n2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 1.72748
R9646 a_41271_20992.t0 a_41271_20992.t1 65.941
R9647 a_42781_12280.t0 a_42781_12280.t1 114.052
R9648 top_segment_1_0.rseg_1_v3_1.v28 top_segment_1_0.rseg_1_v3_1.v28.t0 249.328
R9649 top_segment_1_0.rseg_1_v3_1.v28.n0 top_segment_1_0.rseg_1_v3_1.v28.t2 10.5296
R9650 top_segment_1_0.rseg_1_v3_1.v28.n0 top_segment_1_0.rseg_1_v3_1.v28.t1 10.5285
R9651 top_segment_1_0.rseg_1_v3_1.v28 top_segment_1_0.rseg_1_v3_1.v28.n0 2.13671
R9652 a_19203_9019.n0 a_19203_9019.t2 667.841
R9653 a_19203_9019.n0 a_19203_9019.t1 667.491
R9654 a_19203_9019.t0 a_19203_9019.n0 665.484
R9655 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t1 675.929
R9656 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t0 10.8299
R9657 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t2 10.6741
R9658 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.n0 4.11253
R9659 top_segment_1_0.rseg_1_v3_1.v6 top_segment_1_0.rseg_1_v3_1.v6.t1 248.484
R9660 top_segment_1_0.rseg_1_v3_1.v6.n0 top_segment_1_0.rseg_1_v3_1.v6.t0 10.5338
R9661 top_segment_1_0.rseg_1_v3_1.v6.n0 top_segment_1_0.rseg_1_v3_1.v6.t2 10.5285
R9662 top_segment_1_0.rseg_1_v3_1.v6 top_segment_1_0.rseg_1_v3_1.v6.n0 3.63285
R9663 a_42271_5944.t0 a_42271_5944.t1 55.3905
R9664 a_42271_13864.t0 a_42271_13864.t1 55.3905
R9665 a_42781_12914.t0 a_42781_12914.t1 114.052
R9666 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t2 663.232
R9667 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t1 10.6701
R9668 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v49.n0 10.5739
R9669 DIN8.n1 DIN8.t3 212.081
R9670 DIN8.n0 DIN8.t2 212.081
R9671 DIN8.n2 DIN8.n1 183.185
R9672 DIN8.n1 DIN8.t1 139.78
R9673 DIN8.n0 DIN8.t0 139.78
R9674 DIN8.n1 DIN8.n0 61.346
R9675 DIN8 DIN8.n2 14.2776
R9676 DIN8.n2 DIN8 5.8885
R9677 top_segment_3_0.rseg_3_v3_0.v15.n0 top_segment_3_0.rseg_3_v3_0.v15.t2 666.722
R9678 top_segment_3_0.rseg_3_v3_0.v15.n0 top_segment_3_0.rseg_3_v3_0.v15.t1 10.6321
R9679 top_segment_3_0.rseg_3_v3_0.v15.t0 top_segment_3_0.rseg_3_v3_0.v15.n0 10.5295
R9680 a_13921_18854.t0 a_13921_18854.n0 671.848
R9681 a_13921_18854.n0 a_13921_18854.t2 666.814
R9682 a_13921_18854.n0 a_13921_18854.t1 665.327
R9683 top_segment_1_0.rseg_1_v3_1.v61 top_segment_1_0.rseg_1_v3_1.v61.t2 249.321
R9684 top_segment_1_0.rseg_1_v3_1.v61.n0 top_segment_1_0.rseg_1_v3_1.v61.t1 10.6701
R9685 top_segment_1_0.rseg_1_v3_1.v61.n0 top_segment_1_0.rseg_1_v3_1.v61.t0 10.5739
R9686 top_segment_1_0.rseg_1_v3_1.v61 top_segment_1_0.rseg_1_v3_1.v61.n0 1.53658
R9687 a_27705_5238.n2 a_27705_5238.t3 248.469
R9688 a_27705_5238.n0 a_27705_5238.t4 246.486
R9689 a_27705_5238.n1 a_27705_5238.t2 244.054
R9690 a_27705_5238.n0 a_27705_5238.t1 239.816
R9691 a_27705_5238.t0 a_27705_5238.n2 239.816
R9692 a_27705_5238.n2 a_27705_5238.n1 5.54425
R9693 a_27705_5238.n1 a_27705_5238.n0 1.47758
R9694 a_42271_14300.t0 a_42271_14300.t1 55.3905
R9695 a_22130_19162.n1 a_22130_19162.t3 249.335
R9696 a_22130_19162.n0 a_22130_19162.t1 247.23
R9697 a_22130_19162.n0 a_22130_19162.t2 241.299
R9698 a_22130_19162.t0 a_22130_19162.n1 239.248
R9699 a_22130_19162.n1 a_22130_19162.n0 2.10675
R9700 a_13219_17684.t0 a_13219_17684.n1 671.525
R9701 a_13219_17684.n0 a_13219_17684.t2 668.735
R9702 a_13219_17684.n1 a_13219_17684.t3 666.038
R9703 a_13219_17684.n0 a_13219_17684.t1 665.865
R9704 a_13219_17684.n1 a_13219_17684.n0 0.365083
R9705 top_segment_1_0.rseg_1_v3_1.v63.n0 top_segment_1_0.rseg_1_v3_1.v63.t2 240.469
R9706 top_segment_1_0.rseg_1_v3_1.v63.t0 top_segment_1_0.rseg_1_v3_1.v63.n0 10.6713
R9707 top_segment_1_0.rseg_1_v3_1.v63.n0 top_segment_1_0.rseg_1_v3_1.v63.t1 10.5739
R9708 a_43570_20676.t0 a_43570_20676.t1 49.8467
R9709 a_42609_19929.t0 a_42609_19929.t1 129.28
R9710 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t0 675.904
R9711 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t2 10.7799
R9712 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.t1 10.6965
R9713 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29.n0 1.35813
R9714 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t1 675.929
R9715 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t0 10.8167
R9716 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t2 10.6741
R9717 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.n0 4.10816
R9718 a_13337_17684.n0 a_13337_17684.t2 670.26
R9719 a_13337_17684.n0 a_13337_17684.t1 667.083
R9720 a_13337_17684.t0 a_13337_17684.n0 665.481
R9721 a_42245_6774.t0 a_42245_6774.n0 228.04
R9722 a_42245_6774.n0 a_42245_6774.t2 145.648
R9723 a_42245_6774.n0 a_42245_6774.t1 83.2159
R9724 a_42609_18149.t0 a_42609_18149.t1 129.28
R9725 a_43026_2518.t0 a_43026_2518.t1 49.8467
R9726 a_43026_2886.t0 a_43026_2886.t1 49.8467
R9727 a_41529_19226.t0 a_41529_19226.t1 65.941
R9728 a_41787_19226.t0 a_41787_19226.t1 65.941
R9729 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t1 675.975
R9730 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t2 10.7153
R9731 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t0 10.6746
R9732 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.n0 2.05556
R9733 top_segment_1_0.rseg_1_v3_1.v43 top_segment_1_0.rseg_1_v3_1.v43.t1 248.95
R9734 top_segment_1_0.rseg_1_v3_1.v43.n0 top_segment_1_0.rseg_1_v3_1.v43.t0 10.575
R9735 top_segment_1_0.rseg_1_v3_1.v43.n0 top_segment_1_0.rseg_1_v3_1.v43.t2 10.5739
R9736 top_segment_1_0.rseg_1_v3_1.v43 top_segment_1_0.rseg_1_v3_1.v43.n0 2.81389
R9737 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t1 663.232
R9738 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.n0 10.6701
R9739 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v1.t2 10.5739
R9740 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t2 674.658
R9741 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t0 10.7653
R9742 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t1 10.7376
R9743 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.n0 4.0963
R9744 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t2 676.321
R9745 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t0 13.5004
R9746 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t1 10.7723
R9747 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.n0 4.72836
R9748 a_43570_20952.t0 a_43570_20952.t1 49.8467
R9749 top_segment_1_0.rseg_1_v3_1.v13 top_segment_1_0.rseg_1_v3_1.v13.t2 249.321
R9750 top_segment_1_0.rseg_1_v3_1.v13.n0 top_segment_1_0.rseg_1_v3_1.v13.t1 10.575
R9751 top_segment_1_0.rseg_1_v3_1.v13.n0 top_segment_1_0.rseg_1_v3_1.v13.t0 10.5739
R9752 top_segment_1_0.rseg_1_v3_1.v13 top_segment_1_0.rseg_1_v3_1.v13.n0 1.60689
R9753 a_41714_3346.t0 a_41714_3346.t1 49.8467
R9754 top_segment_2_0.rseg_2_v3_0.v45.n0 top_segment_2_0.rseg_2_v3_0.v45.t2 238.496
R9755 top_segment_2_0.rseg_2_v3_0.v45.t0 top_segment_2_0.rseg_2_v3_0.v45.n0 10.7268
R9756 top_segment_2_0.rseg_2_v3_0.v45.n0 top_segment_2_0.rseg_2_v3_0.v45.t1 10.6617
R9757 a_42609_19217.t0 a_42609_19217.t1 129.28
R9758 a_42271_7370.t0 a_42271_7370.t1 55.3905
R9759 a_41529_18144.t0 a_41529_18144.t1 65.941
R9760 a_41787_18144.t0 a_41787_18144.t1 65.941
R9761 a_38483_21071.n0 a_38483_21071.t2 356.854
R9762 a_38483_21071.n0 a_38483_21071.t0 15.3866
R9763 a_38483_21071.t1 a_38483_21071.n0 15.3866
R9764 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t2 743.367
R9765 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t0 223.315
R9766 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.t1 152.889
R9767 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[1] 15.4066
R9768 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n0 12.2462
R9769 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_1.Y 2.22659
R9770 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/lvsf_0.IN.n1 1.55202
R9771 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[1] 0.84425
R9772 a_42802_2426.t0 a_42802_2426.t1 49.8467
R9773 a_42271_9904.t0 a_42271_9904.t1 55.3905
R9774 a_42271_10894.t0 a_42271_10894.t1 55.3905
R9775 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t0 675.533
R9776 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t2 10.7605
R9777 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.n0 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.t1 10.7175
R9778 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43.n0 2.73151
R9779 a_42271_11330.t0 a_42271_11330.t1 55.3905
R9780 top_segment_1_0.rseg_1_v3_1.v22 top_segment_1_0.rseg_1_v3_1.v22.t0 247.119
R9781 top_segment_1_0.rseg_1_v3_1.v22.n0 top_segment_1_0.rseg_1_v3_1.v22.t1 10.5296
R9782 top_segment_1_0.rseg_1_v3_1.v22.n0 top_segment_1_0.rseg_1_v3_1.v22.t2 10.5285
R9783 top_segment_1_0.rseg_1_v3_1.v22 top_segment_1_0.rseg_1_v3_1.v22.n0 3.54349
R9784 top_segment_2_0.rseg_2_v3_0.v31.t0 top_segment_2_0.rseg_2_v3_0.v31.n0 237.343
R9785 top_segment_2_0.rseg_2_v3_0.v31.n0 top_segment_2_0.rseg_2_v3_0.v31.t1 10.6247
R9786 top_segment_2_0.rseg_2_v3_0.v31.n0 top_segment_2_0.rseg_2_v3_0.v31.t2 10.5285
R9787 top_segment_1_0.rseg_1_v3_1.v14 top_segment_1_0.rseg_1_v3_1.v14.t2 249.623
R9788 top_segment_1_0.rseg_1_v3_1.v14.n0 top_segment_1_0.rseg_1_v3_1.v14.t1 10.5309
R9789 top_segment_1_0.rseg_1_v3_1.v14.n0 top_segment_1_0.rseg_1_v3_1.v14.t0 10.5295
R9790 top_segment_1_0.rseg_1_v3_1.v14 top_segment_1_0.rseg_1_v3_1.v14.n0 0.915451
R9791 a_41529_18542.t0 a_41529_18542.t1 65.941
R9792 a_43890_2242.t0 a_43890_2242.t1 49.8467
R9793 top_segment_1_0.rseg_1_v3_1.v23 top_segment_1_0.rseg_1_v3_1.v23.t0 248.075
R9794 top_segment_1_0.rseg_1_v3_1.v23.n0 top_segment_1_0.rseg_1_v3_1.v23.t1 10.6701
R9795 top_segment_1_0.rseg_1_v3_1.v23.n0 top_segment_1_0.rseg_1_v3_1.v23.t2 10.5739
R9796 top_segment_1_0.rseg_1_v3_1.v23 top_segment_1_0.rseg_1_v3_1.v23.n0 4.17455
R9797 a_41938_2698.t0 a_41938_2698.t1 49.8467
R9798 a_42781_13904.t0 a_42781_13904.t1 114.052
R9799 top_segment_1_0.rseg_1_v3_1.v41 top_segment_1_0.rseg_1_v3_1.v41.t2 249.345
R9800 top_segment_1_0.rseg_1_v3_1.v41.n0 top_segment_1_0.rseg_1_v3_1.v41.t1 10.575
R9801 top_segment_1_0.rseg_1_v3_1.v41.n0 top_segment_1_0.rseg_1_v3_1.v41.t0 10.5739
R9802 top_segment_1_0.rseg_1_v3_1.v41 top_segment_1_0.rseg_1_v3_1.v41.n0 4.20348
R9803 a_42781_16240.t0 a_42781_16240.t1 114.052
R9804 a_41529_17460.t0 a_41529_17460.t1 65.941
R9805 a_43570_19528.t0 a_43570_19528.t1 49.8467
R9806 ROUT.n1 ROUT.t3 134.847
R9807 ROUT.n2 ROUT.t1 134.246
R9808 ROUT.n3 ROUT 13.0108
R9809 ROUT.n1 ROUT.n0 8.36161
R9810 ROUT.t5 ROUT.t4 5.8809
R9811 ROUT.t2 ROUT.t5 5.0615
R9812 ROUT.n0 ROUT.t0 2.9407
R9813 ROUT.n0 ROUT.t2 2.9407
R9814 ROUT.n2 ROUT.n1 0.601043
R9815 ROUT.n3 ROUT.n2 0.271587
R9816 ROUT ROUT.n3 0.023
R9817 a_42541_21510.n0 a_42541_21510.t3 135.572
R9818 a_42541_21510.n1 a_42541_21510.t0 135.572
R9819 a_42541_21510.n0 a_42541_21510.t2 134.246
R9820 a_42541_21510.t1 a_42541_21510.n1 134.246
R9821 a_42541_21510.n1 a_42541_21510.n0 1.1418
R9822 a_13889_17684.n0 a_13889_17684.t2 670.384
R9823 a_13889_17684.n0 a_13889_17684.t1 668.327
R9824 a_13889_17684.t0 a_13889_17684.n0 665.848
R9825 a_42271_6934.t0 a_42271_6934.t1 55.3905
R9826 a_41529_20650.t0 a_41529_20650.t1 65.941
C0 SH[2] SH[1] 19.066f
C1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.0386f
C2 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v14 0.02042f
C3 VL3 top_segment_4_1.b3 0.32205f
C4 SH[2] top_segment_2_0.DEC2[0] 0.04929f
C5 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.18677f
C6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.07012f
C7 a_36142_18450# a_36284_18467# 0.04234f
C8 a_38408_21045# VDDH 0.2924f
C9 VDDH top_segment_3_0.b[5] 1.54847f
C10 top_segment_3_0.b[6] top_segment_4_1.DEC2 0.09f
C11 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 1.95031f
C12 top_segment_2_0.DEC0[2] top_segment_3_0.bb[5] 0.0436f
C13 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC2[2] 0.02204f
C14 top_segment_2_0.DEC0[1] VDDH 0.89706f
C15 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.05882f
C16 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_4_1.DEC3 0.01611f
C17 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.14262f
C18 VH3 top_segment_4_1.bb3 0.31565f
C19 top_segment_2_0.DEC0[2] top_segment_4_1.bb3 0.04843f
C20 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04786f
C21 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.02165f
C22 a_43890_3816# top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.01719f
C23 SH[2] top_segment_4_1.bb1 0.09502f
C24 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_4_1.DEC1 0.04402f
C25 DIN1 DIN2 0.33f
C26 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 1.33533f
C27 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.16197f
C28 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.26736f
C29 top_segment_2_0.DEC0[0] top_segment_3_0.bb[5] 0.0436f
C30 top_segment_3_0.bb[4] top_segment_2_0.DEC2[2] 0.09591f
C31 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 1.3467f
C32 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 0.10095f
C33 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.04529f
C34 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v39 0.23003f
C35 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC1[0] 0.43649f
C36 top_segment_2_0.DEC0[0] top_segment_4_1.bb3 0.04843f
C37 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.24261f
C38 top_segment_1_0.rseg_1_v3_1.v24 top_segment_1_0.rseg_1_v3_1.v39 0.04787f
C39 VDD DIN3 0.67007f
C40 top_segment_1_0.rseg_1_v3_1.v28 top_segment_1_0.rseg_1_v3_1.v35 0.03392f
C41 top_segment_1_0.rseg_1_v3_1.v26 top_segment_1_0.rseg_1_v3_1.v37 0.02766f
C42 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.10926f
C43 top_segment_4_1.bb3 top_segment_4_1.bb2 0.10465f
C44 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.10472f
C45 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.13238f
C46 top_segment_2_0.DEC1[2] top_segment_2_0.DEC1[3] 17.3168f
C47 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_35569_19283# 0.01181f
C48 SH[3] top_segment_4_1.b2 0.09762f
C49 top_segment_2_0.DEC1[2] top_segment_2_0.DEC2[0] 0.04931f
C50 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.05884f
C51 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.04684f
C52 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC0[1] 0.15469f
C53 top_segment_4_1.DEC3 top_segment_4_1.bb2 0.05186f
C54 VDDH top_segment_2_0.DEC2[2] 1.30585f
C55 top_segment_4_1.DEC1 top_segment_4_1.bb2 0.04792f
C56 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v38 0.0857f
C57 top_segment_1_0.rseg_1_v3_1.v61 top_segment_1_0.rseg_1_v3_1.v62 1.25122f
C58 a_38315_19653# a_38315_19377# 0.02286f
C59 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_37164_18842# 0.01035f
C60 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.11542f
C61 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.0151f
C62 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV SH[2] 0.01125f
C63 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.41311f
C64 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.0583f
C65 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 VDDH 3.10831f
C66 DIN8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.01582f
C67 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_38408_20445# 0.06598f
C68 top_segment_3_0.bb[5] top_segment_3_0.b[5] 17.3348f
C69 SH[1] top_segment_4_1.b2 0.12742f
C70 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B VDD 0.25878f
C71 VH2 top_segment_2_0.DEC2[2] 0.31312f
C72 top_segment_2_0.DEC0[1] top_segment_3_0.bb[5] 0.04362f
C73 top_segment_2_0.DEC2[0] top_segment_4_1.b2 0.04942f
C74 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 1.32352f
C75 top_segment_1_0.rseg_1_v3_1.v13 top_segment_1_0.rseg_1_v3_1.v14 1.16723f
C76 top_segment_3_0.b[5] top_segment_4_1.bb3 0.05224f
C77 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC2[2] 0.07846f
C78 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v37 0.20454f
C79 top_segment_1_0.rseg_1_v3_1.v60 top_segment_1_0.rseg_1_v3_1.v62 1.15664f
C80 top_segment_2_0.DEC0[1] top_segment_4_1.bb3 0.04843f
C81 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.21766f
C82 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 0.10974f
C83 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 2.97868f
C84 top_segment_3_0.b[6] top_segment_2_0.DEC1[3] 0.03535f
C85 top_segment_4_1.DEC3 top_segment_3_0.b[5] 0.09294f
C86 top_segment_2_0.DEC1[1] top_segment_2_0.DEC1[3] 0.50988f
C87 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.60657f
C88 top_segment_3_0.b[6] top_segment_2_0.DEC2[0] 0.09013f
C89 top_segment_2_0.DEC1[1] top_segment_2_0.DEC2[0] 0.10018f
C90 top_segment_4_1.b2 top_segment_4_1.bb1 0.09973f
C91 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.21449f
C92 top_segment_4_1.bb2 top_segment_4_1.b1 14.2376f
C93 top_segment_3_0.b[5] top_segment_4_1.DEC1 0.08819f
C94 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 VDDH 6.21616f
C95 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC2[3] 0.18654f
C96 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 3.68198f
C97 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.04651f
C98 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.29277f
C99 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v10 0.01136f
C100 VDDH SH[2] 0.58996f
C101 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC1[2] 0.02122f
C102 top_segment_1_0.rseg_1_v3_1.v12 top_segment_1_0.rseg_1_v3_1.v14 1.15763f
C103 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y VDD 0.49613f
C104 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC2[1] 0.26638f
C105 top_segment_1_0.rseg_1_v3_1.v60 top_segment_1_0.rseg_1_v3_1.v61 1.24381f
C106 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v36 0.14746f
C107 top_segment_1_0.rseg_1_v3_1.v59 top_segment_1_0.rseg_1_v3_1.v62 0.0119f
C108 a_38408_20445# VDDH 0.40618f
C109 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.01833f
C110 top_segment_3_0.bb[5] top_segment_2_0.DEC2[2] 0.09114f
C111 VDDH top_segment_1_0.rseg_1_v3_1.v40 0.09915f
C112 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.01844f
C113 top_segment_3_0.bb[6] top_segment_4_1.DEC2 0.10492f
C114 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC a_38315_19653# 0.01079f
C115 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B 0.18203f
C116 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.20535f
C117 top_segment_2_0.DEC1[2] top_segment_3_0.bb[4] 0.04845f
C118 top_segment_4_1.bb3 top_segment_2_0.DEC2[2] 0.09612f
C119 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.58839f
C120 SH[2] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.01383f
C121 VDDH DIN2 0.42749f
C122 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 1.27501f
C123 top_segment_4_1.b3 top_segment_4_1.DEC2 0.10421f
C124 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.04477f
C125 top_segment_1_0.rseg_1_v3_1.v12 top_segment_1_0.rseg_1_v3_1.v13 1.15809f
C126 top_segment_1_0.rseg_1_v3_1.v11 top_segment_1_0.rseg_1_v3_1.v14 0.0119f
C127 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v35 0.20093f
C128 top_segment_2_0.DEC2[3] top_segment_4_1.DEC2 0.05383f
C129 top_segment_1_0.rseg_1_v3_1.v59 top_segment_1_0.rseg_1_v3_1.v61 1.73155f
C130 top_segment_4_1.DEC3 top_segment_2_0.DEC2[2] 0.35307f
C131 top_segment_1_0.rseg_1_v3_1.v58 top_segment_1_0.rseg_1_v3_1.v62 0.31595f
C132 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.05396f
C133 top_segment_2_0.V0 top_segment_4_1.DEC2 0.11409f
C134 top_segment_1_0.rseg_1_v3_1.v29 top_segment_1_0.rseg_1_v3_1.v22 0.02015f
C135 top_segment_4_1.DEC2 top_segment_2_0.DEC2[1] 0.26895f
C136 top_segment_2_0.DEC2[2] top_segment_4_1.DEC1 0.05025f
C137 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C138 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.12526f
C139 top_segment_2_0.DEC1[0] top_segment_2_0.DEC1[3] 0.53884f
C140 top_segment_1_0.rseg_1_v3_1.v38 top_segment_1_0.rseg_1_v3_1.v39 0.62948f
C141 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.05552f
C142 top_segment_2_0.DEC1[2] VDDH 0.88394f
C143 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_36284_18467# 0.02737f
C144 top_segment_2_0.DEC1[0] top_segment_2_0.DEC2[0] 0.15968f
C145 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.01132f
C146 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.18941f
C147 top_segment_1_0.rseg_1_v3_1.v10 top_segment_1_0.rseg_1_v3_1.v14 0.43907f
C148 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC1[1] 0.02121f
C149 top_segment_1_0.rseg_1_v3_1.v11 top_segment_1_0.rseg_1_v3_1.v13 1.72759f
C150 top_segment_3_0.b[4] top_segment_4_1.DEC2 0.09522f
C151 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_3_0.b[6] 0.11135f
C152 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.04526f
C153 top_segment_3_0.bb[4] top_segment_4_1.b2 0.01389f
C154 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 1.28515f
C155 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 0.0953f
C156 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v34 0.30567f
C157 top_segment_1_0.rseg_1_v3_1.v59 top_segment_1_0.rseg_1_v3_1.v60 1.37492f
C158 top_segment_1_0.rseg_1_v3_1.v58 top_segment_1_0.rseg_1_v3_1.v61 0.0961f
C159 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.33687f
C160 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.09522f
C161 DIN7 DIN8 0.33719f
C162 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 1.13576f
C163 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.7893f
C164 top_segment_1_0.rseg_1_v3_1.v37 top_segment_1_0.rseg_1_v3_1.v39 1.97694f
C165 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.02834f
C166 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.09544f
C167 top_segment_3_0.b[6] top_segment_3_0.bb[4] 0.04882f
C168 top_segment_2_0.DEC1[1] top_segment_3_0.bb[4] 0.04846f
C169 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.6218f
C170 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 0.20568f
C171 SH[2] top_segment_4_1.bb3 0.09759f
C172 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC1[2] 0.11523f
C173 SH[3] top_segment_4_1.b3 0.0966f
C174 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 1.27523f
C175 VDDH top_segment_4_1.b2 1.41293f
C176 top_segment_2_0.DEC2[2] top_segment_4_1.b1 0.04747f
C177 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.05972f
C178 SH[3] top_segment_2_0.DEC2[3] 0.05359f
C179 top_segment_2_0.V0 SH[3] 0.11409f
C180 top_segment_1_0.rseg_1_v3_1.v10 top_segment_1_0.rseg_1_v3_1.v13 0.09535f
C181 top_segment_1_0.rseg_1_v3_1.v11 top_segment_1_0.rseg_1_v3_1.v12 1.2875f
C182 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.02821f
C183 SH[3] top_segment_2_0.DEC2[1] 0.04851f
C184 top_segment_1_0.rseg_1_v3_1.v57 top_segment_1_0.rseg_1_v3_1.v61 0.08493f
C185 top_segment_1_0.rseg_1_v3_1.v58 top_segment_1_0.rseg_1_v3_1.v60 1.89956f
C186 VL2 top_segment_2_0.DEC2[0] 0.18852f
C187 top_segment_1_0.rseg_1_v3_1.v27 top_segment_1_0.rseg_1_v3_1.v22 0.05302f
C188 top_segment_1_0.rseg_1_v3_1.v29 top_segment_1_0.rseg_1_v3_1.v20 0.02197f
C189 SH[2] top_segment_4_1.DEC3 0.05175f
C190 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 0.65201f
C191 SH[2] top_segment_4_1.DEC1 0.04779f
C192 top_segment_1_0.rseg_1_v3_1.v36 top_segment_1_0.rseg_1_v3_1.v39 0.06132f
C193 top_segment_1_0.rseg_1_v3_1.v37 top_segment_1_0.rseg_1_v3_1.v38 0.4572f
C194 top_segment_3_0.b[6] VDDH 2.1953f
C195 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.09312f
C196 top_segment_2_0.DEC1[1] VDDH 0.85743f
C197 VDD DIN7 0.71581f
C198 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.08251f
C199 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.21631f
C200 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_37131_19653# 0.01092f
C201 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] ROUT 0.06337f
C202 top_segment_3_0.bb[6] top_segment_2_0.DEC1[3] 0.05174f
C203 top_segment_3_0.bb[6] top_segment_2_0.DEC2[0] 0.1029f
C204 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC a_38315_19377# 0.02668f
C205 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.21415f
C206 top_segment_1_0.rseg_1_v3_1.v10 top_segment_1_0.rseg_1_v3_1.v12 2.0142f
C207 top_segment_1_0.rseg_1_v3_1.v9 top_segment_1_0.rseg_1_v3_1.v13 0.08427f
C208 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.05244f
C209 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC1[0] 0.02121f
C210 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 1.83395f
C211 top_segment_2_0.DEC1[2] top_segment_3_0.bb[5] 0.04363f
C212 SH[1] top_segment_4_1.b3 0.12916f
C213 VDD DIN8 0.72319f
C214 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.09546f
C215 top_segment_1_0.rseg_1_v3_1.v57 top_segment_1_0.rseg_1_v3_1.v60 0.02715f
C216 top_segment_1_0.rseg_1_v3_1.v56 top_segment_1_0.rseg_1_v3_1.v61 0.21492f
C217 top_segment_1_0.rseg_1_v3_1.v58 top_segment_1_0.rseg_1_v3_1.v59 1.36638f
C218 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 1.32046f
C219 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.06256f
C220 top_segment_2_0.DEC1[3] top_segment_4_1.b3 0.04805f
C221 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.02737f
C222 SH[1] top_segment_2_0.DEC2[3] 0.06598f
C223 top_segment_2_0.DEC1[2] top_segment_4_1.bb3 0.0485f
C224 top_segment_4_1.b3 top_segment_2_0.DEC2[0] 0.09746f
C225 top_segment_2_0.V0 SH[1] 0.18545f
C226 top_segment_2_0.DEC1[3] top_segment_2_0.DEC2[3] 0.12584f
C227 top_segment_2_0.V0 top_segment_2_0.DEC1[3] 0.11848f
C228 SH[1] top_segment_2_0.DEC2[1] 0.06343f
C229 top_segment_2_0.DEC2[3] top_segment_2_0.DEC2[0] 0.48051f
C230 top_segment_1_0.rseg_1_v3_1.v35 top_segment_1_0.rseg_1_v3_1.v39 0.05244f
C231 top_segment_2_0.V0 top_segment_2_0.DEC2[0] 0.11409f
C232 top_segment_1_0.rseg_1_v3_1.v36 top_segment_1_0.rseg_1_v3_1.v38 1.64648f
C233 top_segment_2_0.DEC1[3] top_segment_2_0.DEC2[1] 0.04856f
C234 top_segment_2_0.DEC2[1] top_segment_2_0.DEC2[0] 17.3231f
C235 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.20664f
C236 top_segment_2_0.DEC1[0] top_segment_3_0.bb[4] 0.04847f
C237 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.04626f
C238 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.02163f
C239 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.1866f
C240 DIN6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.03492f
C241 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.02139f
C242 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.0921f
C243 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC1[1] 0.09505f
C244 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.29779f
C245 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.64353f
C246 VDD DIN0 0.71624f
C247 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 1.27264f
C248 top_segment_4_1.b3 top_segment_4_1.bb1 0.11032f
C249 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.02873f
C250 top_segment_1_0.rseg_1_v3_1.v10 top_segment_1_0.rseg_1_v3_1.v11 1.27692f
C251 top_segment_1_0.rseg_1_v3_1.v8 top_segment_1_0.rseg_1_v3_1.v13 0.2143f
C252 top_segment_1_0.rseg_1_v3_1.v9 top_segment_1_0.rseg_1_v3_1.v12 0.02715f
C253 top_segment_2_0.DEC2[3] top_segment_4_1.bb1 0.05175f
C254 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.28898f
C255 SH[2] top_segment_4_1.b1 0.09468f
C256 top_segment_1_0.rseg_1_v3_1.v57 top_segment_1_0.rseg_1_v3_1.v59 1.79255f
C257 top_segment_2_0.V0 top_segment_4_1.bb1 0.61294f
C258 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v23 0.15222f
C259 top_segment_2_0.DEC1[3] top_segment_3_0.b[4] 0.04329f
C260 top_segment_2_0.DEC2[1] top_segment_4_1.bb1 0.04858f
C261 top_segment_1_0.rseg_1_v3_1.v24 top_segment_1_0.rseg_1_v3_1.v23 0.10072f
C262 top_segment_1_0.rseg_1_v3_1.v25 top_segment_1_0.rseg_1_v3_1.v22 0.04732f
C263 top_segment_1_0.rseg_1_v3_1.v29 top_segment_1_0.rseg_1_v3_1.v18 0.02163f
C264 top_segment_1_0.rseg_1_v3_1.v27 top_segment_1_0.rseg_1_v3_1.v20 0.02198f
C265 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 0.47118f
C266 top_segment_3_0.b[4] top_segment_2_0.DEC2[0] 0.09272f
C267 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 1.9819f
C268 top_segment_1_0.rseg_1_v3_1.v36 top_segment_1_0.rseg_1_v3_1.v37 0.57403f
C269 top_segment_1_0.rseg_1_v3_1.v34 top_segment_1_0.rseg_1_v3_1.v39 0.05777f
C270 top_segment_2_0.DEC1[0] VDDH 0.88599f
C271 top_segment_4_1.bb3 top_segment_4_1.b2 14.2467f
C272 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.0259f
C273 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.29614f
C274 VDD ROUT 0.6068f
C275 top_segment_1_0.rseg_1_v3_1.v9 top_segment_1_0.rseg_1_v3_1.v11 1.78725f
C276 top_segment_3_0.b[6] top_segment_3_0.bb[5] 0.20876f
C277 top_segment_2_0.DEC1[1] top_segment_3_0.bb[5] 0.04366f
C278 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C279 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.05244f
C280 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 1.81409f
C281 top_segment_4_1.DEC3 top_segment_4_1.b2 0.05188f
C282 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.21631f
C283 top_segment_1_0.rseg_1_v3_1.v57 top_segment_1_0.rseg_1_v3_1.v58 1.34945f
C284 top_segment_1_0.rseg_1_v3_1.v56 top_segment_1_0.rseg_1_v3_1.v59 0.09809f
C285 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 1.34913f
C286 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.09546f
C287 a_43890_3816# top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.01335f
C288 top_segment_1_0.rseg_1_v3_1.v24 top_segment_1_0.rseg_1_v3_1.v22 1.73509f
C289 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v22 0.1278f
C290 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_3_0.bb[6] 0.07088f
C291 VDDH top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.90617f
C292 top_segment_2_0.DEC1[1] top_segment_4_1.bb3 0.04851f
C293 top_segment_4_1.DEC1 top_segment_4_1.b2 0.04795f
C294 top_segment_2_0.DEC0[2] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 17.0519f
C295 top_segment_3_0.b[6] top_segment_4_1.bb3 0.05544f
C296 top_segment_1_0.rseg_1_v3_1.v35 top_segment_1_0.rseg_1_v3_1.v37 1.45085f
C297 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v14 0.15587f
C298 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.14089f
C299 top_segment_3_0.b[6] top_segment_4_1.DEC3 0.08857f
C300 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC1[0] 0.09358f
C301 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.02163f
C302 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.13214f
C303 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.02218f
C304 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.04735f
C305 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC2[3] 0.02136f
C306 SH[4] top_segment_4_1.bb2 0.09808f
C307 top_segment_2_0.DEC0[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.93455f
C308 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.66863f
C309 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.2656f
C310 top_segment_3_0.b[6] top_segment_4_1.DEC1 0.09146f
C311 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC2[1] 0.02207f
C312 top_segment_3_0.bb[6] top_segment_3_0.bb[4] 0.073f
C313 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C314 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C315 top_segment_1_0.rseg_1_v3_1.v9 top_segment_1_0.rseg_1_v3_1.v10 1.25806f
C316 top_segment_1_0.rseg_1_v3_1.v8 top_segment_1_0.rseg_1_v3_1.v11 0.0981f
C317 VDDH DIN6 0.42765f
C318 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.0203f
C319 top_segment_1_0.rseg_1_v3_1.v56 top_segment_1_0.rseg_1_v3_1.v58 0.55355f
C320 VS4 top_segment_4_1.b3 0.04487f
C321 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v21 0.06072f
C322 top_segment_1_0.rseg_1_v3_1.v14 top_segment_1_0.rseg_1_v3_1.v23 0.01643f
C323 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.15973f
C324 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.05823f
C325 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.04809f
C326 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.5508f
C327 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.11272f
C328 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.01028f
C329 top_segment_3_0.bb[4] top_segment_4_1.b3 14.4527f
C330 DIN2 DIN3 0.33146f
C331 VDDH top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.01032f
C332 top_segment_1_0.rseg_1_v3_1.v35 top_segment_1_0.rseg_1_v3_1.v36 0.57986f
C333 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 1.97214f
C334 top_segment_2_0.DEC2[3] top_segment_3_0.bb[4] 0.10026f
C335 top_segment_1_0.rseg_1_v3_1.v34 top_segment_1_0.rseg_1_v3_1.v37 0.04811f
C336 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v13 0.17825f
C337 top_segment_2_0.V0 top_segment_3_0.bb[4] 0.11409f
C338 top_segment_3_0.bb[4] top_segment_2_0.DEC2[1] 0.09785f
C339 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] VDD 1.24016f
C340 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 11.41f
C341 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_3_0.b[4] 0.01148f
C342 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.10009f
C343 top_segment_3_0.bb[6] VDDH 2.618f
C344 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.03366f
C345 VS1 top_segment_4_1.bb3 0.02487f
C346 VDD DIN5 0.67364f
C347 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.04942f
C348 top_segment_4_1.b2 top_segment_4_1.b1 0.31778f
C349 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.18751f
C350 top_segment_1_0.rseg_1_v3_1.v8 top_segment_1_0.rseg_1_v3_1.v10 0.54398f
C351 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 VDDH 2.32429f
C352 top_segment_2_0.DEC1[0] top_segment_3_0.bb[5] 0.04368f
C353 top_segment_1_0.rseg_1_v3_1.v56 top_segment_1_0.rseg_1_v3_1.v57 3.83937f
C354 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.05253f
C355 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.04039f
C356 VH2 VL2 1.05021f
C357 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 1.81035f
C358 a_35360_18748# a_35360_18450# 0.015f
C359 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v20 0.03142f
C360 VDDH top_segment_4_1.b3 2.54466f
C361 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 0.09544f
C362 top_segment_2_0.DEC1[0] top_segment_4_1.bb3 0.04852f
C363 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 1.37192f
C364 VDDH top_segment_2_0.DEC2[3] 1.39235f
C365 top_segment_3_0.b[4] top_segment_3_0.bb[4] 15.8859f
C366 top_segment_2_0.V0 VDDH 0.0402f
C367 VDDH top_segment_2_0.DEC2[1] 1.26896f
C368 top_segment_1_0.rseg_1_v3_1.v34 top_segment_1_0.rseg_1_v3_1.v36 1.22987f
C369 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 0.09468f
C370 VDDH top_segment_1_0.rseg_1_v3_1.v24 0.10118f
C371 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 1.16961f
C372 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v12 0.09116f
C373 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.09623f
C374 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A VDD 1.0555f
C375 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 4.16288f
C376 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_3_0.b[5] 0.05551f
C377 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.16418f
C378 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.0249f
C379 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.02218f
C380 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.04751f
C381 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.02156f
C382 top_segment_2_0.DEC0[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.72578f
C383 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.05999f
C384 top_segment_1_0.rseg_1_v3_1.v8 top_segment_1_0.rseg_1_v3_1.v9 3.76093f
C385 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 1.04282f
C386 top_segment_2_0.DEC0[2] ROUT 0.02421f
C387 VDDH top_segment_3_0.b[4] 2.06537f
C388 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v19 0.03135f
C389 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.07818f
C390 VH2 top_segment_2_0.DEC2[3] 0.37249f
C391 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.578f
C392 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.04811f
C393 top_segment_1_0.rseg_1_v3_1.v34 top_segment_1_0.rseg_1_v3_1.v35 0.66352f
C394 VH2 top_segment_2_0.DEC2[1] 0.47342f
C395 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 1.97317f
C396 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.30168f
C397 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC2[3] 0.12411f
C398 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v11 0.09117f
C399 top_segment_2_0.DEC0[0] ROUT 0.01445f
C400 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC2[1] 0.06721f
C401 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.04638f
C402 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.09624f
C403 VDDH top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.01046f
C404 SH[4] top_segment_2_0.DEC2[2] 0.04736f
C405 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v18 0.06065f
C406 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 1.79741f
C407 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.05244f
C408 top_segment_1_0.rseg_1_v3_1.v24 top_segment_1_0.rseg_1_v3_1.v18 0.0119f
C409 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_38315_19653# 0.03153f
C410 top_segment_3_0.bb[6] top_segment_3_0.bb[5] 0.04811f
C411 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_2_0.DEC2[2] 0.06295f
C412 SH[3] top_segment_4_1.DEC2 0.05177f
C413 top_segment_3_0.bb[6] top_segment_4_1.bb3 0.1782f
C414 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v10 0.17828f
C415 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC1[3] 0.55413f
C416 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.05843f
C417 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 0.33228f
C418 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.09942f
C419 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC2[0] 0.42123f
C420 top_segment_3_0.bb[5] top_segment_4_1.b3 0.31045f
C421 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05095f
C422 a_43562_3816# VDD 0.03791f
C423 VDDH VL3 0.10866f
C424 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.0152f
C425 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 4.12073f
C426 top_segment_2_0.DEC2[3] top_segment_3_0.bb[5] 0.09548f
C427 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.01429f
C428 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.02254f
C429 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.04788f
C430 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 0.02199f
C431 top_segment_2_0.V0 top_segment_3_0.bb[5] 0.11409f
C432 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.19295f
C433 top_segment_4_1.b3 top_segment_4_1.bb3 15.6923f
C434 top_segment_3_0.bb[6] top_segment_4_1.DEC3 0.10426f
C435 top_segment_3_0.bb[5] top_segment_2_0.DEC2[1] 0.09312f
C436 VDDH top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.90804f
C437 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.10646f
C438 a_43284_3816# top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.02083f
C439 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.03386f
C440 top_segment_2_0.DEC2[3] top_segment_4_1.bb3 0.10029f
C441 top_segment_2_0.V0 top_segment_4_1.bb3 0.13343f
C442 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 9.03926f
C443 top_segment_3_0.bb[6] top_segment_4_1.DEC1 0.10201f
C444 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.10246f
C445 top_segment_1_0.rseg_1_v3_1.v10 top_segment_1_0.rseg_1_v3_1.v23 1.34685f
C446 top_segment_1_0.rseg_1_v3_1.v12 top_segment_1_0.rseg_1_v3_1.v21 0.0266f
C447 top_segment_1_0.rseg_1_v3_1.v14 top_segment_1_0.rseg_1_v3_1.v19 0.02541f
C448 top_segment_4_1.bb3 top_segment_2_0.DEC2[1] 0.4374f
C449 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC0[2] 0.01854f
C450 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.02665f
C451 VDDH DIN4 0.42749f
C452 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.02537f
C453 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 1.48f
C454 VDDH top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.01064f
C455 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.01148f
C456 top_segment_4_1.DEC3 top_segment_4_1.b3 0.09992f
C457 a_36142_18748# a_36142_18450# 0.015f
C458 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.60845f
C459 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.04843f
C460 top_segment_2_0.DEC2[3] top_segment_4_1.DEC3 0.64599f
C461 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v9 0.15598f
C462 top_segment_4_1.b3 top_segment_4_1.DEC1 0.4087f
C463 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 1.05222f
C464 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 1.96808f
C465 top_segment_2_0.V0 top_segment_4_1.DEC3 0.11409f
C466 top_segment_4_1.DEC3 top_segment_2_0.DEC2[1] 0.20774f
C467 SH[1] top_segment_4_1.DEC2 0.06246f
C468 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.08664f
C469 top_segment_2_0.DEC2[3] top_segment_4_1.DEC1 0.05329f
C470 top_segment_2_0.DEC0[1] ROUT 0.0162f
C471 top_segment_2_0.V0 top_segment_4_1.DEC1 0.11409f
C472 top_segment_3_0.bb[5] top_segment_3_0.b[4] 14.0478f
C473 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 0.18469f
C474 top_segment_2_0.DEC2[1] top_segment_4_1.DEC1 0.58792f
C475 top_segment_4_1.DEC2 top_segment_2_0.DEC2[0] 0.11771f
C476 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC0[0] 0.01806f
C477 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.15933f
C478 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B VDD 0.4727f
C479 top_segment_3_0.b[4] top_segment_4_1.bb3 0.20364f
C480 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04695f
C481 top_segment_1_0.rseg_1_v3_1.v54 top_segment_1_0.rseg_1_v3_1.v61 0.02015f
C482 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.06718f
C483 top_segment_2_0.DEC0[2] top_segment_2_0.DEC0[0] 0.69498f
C484 top_segment_4_1.DEC3 top_segment_3_0.b[4] 0.09515f
C485 top_segment_4_1.DEC2 top_segment_4_1.bb1 0.05602f
C486 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v8 0.1529f
C487 top_segment_3_0.b[4] top_segment_4_1.DEC1 0.17416f
C488 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05297f
C489 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 4.13148f
C490 a_43284_3816# top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.04364f
C491 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.38958f
C492 top_segment_1_0.rseg_1_v3_1.v10 top_segment_1_0.rseg_1_v3_1.v21 0.02839f
C493 top_segment_1_0.rseg_1_v3_1.v12 top_segment_1_0.rseg_1_v3_1.v19 0.03446f
C494 top_segment_1_0.rseg_1_v3_1.v8 top_segment_1_0.rseg_1_v3_1.v23 0.05173f
C495 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 1.04528f
C496 top_segment_4_1.b3 top_segment_4_1.b1 0.10741f
C497 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.02948f
C498 top_segment_2_0.DEC2[3] top_segment_4_1.b1 0.05183f
C499 top_segment_2_0.V0 top_segment_4_1.b1 0.17102f
C500 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 1.47954f
C501 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.02493f
C502 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.02615f
C503 a_37131_19653# a_37131_19377# 0.02286f
C504 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.04809f
C505 VL3 top_segment_4_1.bb3 0.22736f
C506 top_segment_2_0.DEC2[1] top_segment_4_1.b1 0.04859f
C507 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.64115f
C508 SH[3] top_segment_2_0.DEC2[0] 0.04929f
C509 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.02113f
C510 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC0[1] 0.01814f
C511 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_2_0.DEC1[2] 0.73909f
C512 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C513 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 0.16077f
C514 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.01148f
C515 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 0.31985f
C516 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.38434f
C517 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A VDD 0.35622f
C518 top_segment_1_0.rseg_1_v3_1.v45 top_segment_1_0.rseg_1_v3_1.v46 1.22792f
C519 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.21618f
C520 top_segment_2_0.DEC0[2] top_segment_3_0.b[5] 0.04064f
C521 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y VDD 0.23023f
C522 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_4_1.DEC2 0.02214f
C523 top_segment_1_0.rseg_1_v3_1.v54 top_segment_1_0.rseg_1_v3_1.v59 0.05305f
C524 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.23151f
C525 top_segment_1_0.rseg_1_v3_1.v52 top_segment_1_0.rseg_1_v3_1.v61 0.02197f
C526 SH[3] top_segment_4_1.bb1 0.09558f
C527 top_segment_2_0.DEC0[2] top_segment_2_0.DEC0[1] 18.3073f
C528 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_37164_18842# 0.02826f
C529 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.23151f
C530 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.06984f
C531 DIN7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.0349f
C532 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC VDDH 4.26993f
C533 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.22399f
C534 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B VDD 0.36582f
C535 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.04842f
C536 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.14095f
C537 top_segment_2_0.DEC0[0] top_segment_3_0.b[5] 0.04064f
C538 SH[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.16758f
C539 a_38408_21484# VDDH 1.43189f
C540 top_segment_3_0.bb[4] top_segment_4_1.DEC2 0.10038f
C541 top_segment_2_0.DEC0[1] top_segment_2_0.DEC0[0] 17.6537f
C542 SH[1] top_segment_2_0.DEC2[0] 0.06421f
C543 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 4.14551f
C544 top_segment_2_0.DEC1[3] top_segment_2_0.DEC2[0] 0.04903f
C545 SH[4] top_segment_4_1.b2 0.09767f
C546 top_segment_1_0.rseg_1_v3_1.v44 top_segment_1_0.rseg_1_v3_1.v46 1.15703f
C547 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.15149f
C548 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.15063f
C549 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC2[2] 0.03788f
C550 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 1.19314f
C551 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 9.22813f
C552 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 1.47977f
C553 VDD DIN2 0.66783f
C554 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.02615f
C555 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.02523f
C556 SH[1] top_segment_4_1.bb1 0.12456f
C557 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.09248f
C558 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.01687f
C559 top_segment_2_0.DEC2[0] top_segment_4_1.bb1 0.04937f
C560 VDDH top_segment_4_1.DEC2 3.49035f
C561 top_segment_2_0.DEC0[2] top_segment_2_0.DEC2[2] 0.19079f
C562 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 3.73465f
C563 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_2_0.DEC1[1] 0.06525f
C564 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.01514f
C565 top_segment_3_0.b[6] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.04595f
C566 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.02015f
C567 top_segment_1_0.rseg_1_v3_1.v43 top_segment_1_0.rseg_1_v3_1.v46 0.0119f
C568 top_segment_1_0.rseg_1_v3_1.v44 top_segment_1_0.rseg_1_v3_1.v45 1.21986f
C569 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.06438f
C570 top_segment_1_0.rseg_1_v3_1.v50 top_segment_1_0.rseg_1_v3_1.v61 0.02147f
C571 top_segment_1_0.rseg_1_v3_1.v52 top_segment_1_0.rseg_1_v3_1.v59 0.02201f
C572 top_segment_1_0.rseg_1_v3_1.v55 top_segment_1_0.rseg_1_v3_1.v56 0.17104f
C573 top_segment_1_0.rseg_1_v3_1.v54 top_segment_1_0.rseg_1_v3_1.v57 0.04735f
C574 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.21864f
C575 top_segment_2_0.DEC0[0] top_segment_2_0.DEC2[2] 0.049f
C576 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.18005f
C577 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v46 0.15602f
C578 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] 0.28496f
C579 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 1.73139f
C580 VDDH top_segment_1_0.rseg_1_v3_1.v8 0.11672f
C581 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.10024f
C582 top_segment_2_0.DEC2[2] top_segment_4_1.bb2 0.19372f
C583 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.0707f
C584 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 1.8611f
C585 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 3.28115f
C586 top_segment_2_0.DEC0[1] top_segment_3_0.b[5] 0.04066f
C587 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.0239f
C588 top_segment_1_0.rseg_1_v3_1.v43 top_segment_1_0.rseg_1_v3_1.v45 1.73307f
C589 top_segment_1_0.rseg_1_v3_1.v42 top_segment_1_0.rseg_1_v3_1.v46 0.33336f
C590 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.08581f
C591 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.13238f
C592 top_segment_1_0.rseg_1_v3_1.v13 top_segment_1_0.rseg_1_v3_1.v6 0.02015f
C593 top_segment_1_0.rseg_1_v3_1.v54 top_segment_1_0.rseg_1_v3_1.v56 1.73519f
C594 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 VDDH 2.20196f
C595 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 0.15179f
C596 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.01212f
C597 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.0979f
C598 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV SH[1] 0.01068f
C599 top_segment_1_0.rseg_1_v3_1.v22 top_segment_1_0.rseg_1_v3_1.v23 0.59336f
C600 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.29339f
C601 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC1[3] 0.03108f
C602 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 1.22509f
C603 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v45 0.17853f
C604 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC2[0] 0.02595f
C605 VDDH SH[3] 0.58919f
C606 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.07006f
C607 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05095f
C608 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_2_0.DEC1[0] 0.06658f
C609 DIN3 DIN4 0.3362f
C610 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 0.61284f
C611 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.02015f
C612 VDDH top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.18887f
C613 top_segment_1_0.rseg_1_v3_1.v43 top_segment_1_0.rseg_1_v3_1.v44 1.34563f
C614 top_segment_1_0.rseg_1_v3_1.v42 top_segment_1_0.rseg_1_v3_1.v45 0.09544f
C615 top_segment_2_0.DEC1[3] top_segment_3_0.bb[4] 0.04845f
C616 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.02024f
C617 a_42614_21484# VDDH 1.22217f
C618 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.04287f
C619 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_4_1.bb1 0.01812f
C620 top_segment_3_0.bb[4] top_segment_2_0.DEC2[0] 0.09789f
C621 VDDH DIN9 0.40422f
C622 top_segment_3_0.b[5] top_segment_2_0.DEC2[2] 0.08824f
C623 SH[3] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.1675f
C624 top_segment_3_0.bb[5] top_segment_4_1.DEC2 0.09596f
C625 top_segment_1_0.rseg_1_v3_1.v55 top_segment_1_0.rseg_1_v3_1.v46 0.01649f
C626 top_segment_2_0.DEC0[1] top_segment_2_0.DEC2[2] 0.04875f
C627 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.01131f
C628 top_segment_1_0.rseg_1_v3_1.v21 top_segment_1_0.rseg_1_v3_1.v23 1.97444f
C629 SH[4] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.1675f
C630 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v44 0.09162f
C631 top_segment_4_1.bb3 top_segment_4_1.DEC2 0.10472f
C632 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.10324f
C633 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.4235f
C634 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A VDD 0.32055f
C635 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.06152f
C636 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.3835f
C637 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.12875f
C638 SH[2] top_segment_4_1.bb2 0.09784f
C639 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.01807f
C640 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 1.85532f
C641 top_segment_2_0.DEC2[3] top_segment_1_0.rseg_1_v3_1.v62 0.15788f
C642 VDDH SH[1] 1.7748f
C643 VDDH top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.82663f
C644 VDDH top_segment_2_0.DEC1[3] 0.98177f
C645 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC1[2] 0.01718f
C646 top_segment_4_1.DEC3 top_segment_4_1.DEC2 16.2094f
C647 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v62 0.87032f
C648 VDDH DIN1 0.42749f
C649 VDDH top_segment_2_0.DEC2[0] 1.28968f
C650 top_segment_4_1.DEC2 top_segment_4_1.DEC1 15.5261f
C651 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.14904f
C652 top_segment_1_0.rseg_1_v3_1.v42 top_segment_1_0.rseg_1_v3_1.v44 1.916f
C653 top_segment_1_0.rseg_1_v3_1.v41 top_segment_1_0.rseg_1_v3_1.v45 0.08427f
C654 top_segment_1_0.rseg_1_v3_1.v13 top_segment_1_0.rseg_1_v3_1.v4 0.01848f
C655 top_segment_1_0.rseg_1_v3_1.v11 top_segment_1_0.rseg_1_v3_1.v6 0.04904f
C656 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.07123f
C657 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.22976f
C658 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.15972f
C659 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.22293f
C660 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_36351_19701# 0.0211f
C661 top_segment_2_0.DEC0[2] top_segment_2_0.DEC1[2] 0.94034f
C662 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v43 0.09478f
C663 top_segment_1_0.rseg_1_v3_1.v21 top_segment_1_0.rseg_1_v3_1.v22 0.42912f
C664 top_segment_1_0.rseg_1_v3_1.v20 top_segment_1_0.rseg_1_v3_1.v23 0.06177f
C665 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 1.2479f
C666 VDDH top_segment_4_1.bb1 1.16908f
C667 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.05296f
C668 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 0.56552f
C669 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.05308f
C670 DIN6 DIN7 0.33364f
C671 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 0.0686f
C672 top_segment_2_0.DEC2[3] top_segment_1_0.rseg_1_v3_1.v61 0.17902f
C673 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 1.27914f
C674 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 0.02715f
C675 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 0.21461f
C676 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B VDD 0.25715f
C677 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v61 0.07524f
C678 top_segment_2_0.DEC0[0] top_segment_2_0.DEC1[2] 0.16544f
C679 top_segment_1_0.rseg_1_v3_1.v40 top_segment_1_0.rseg_1_v3_1.v45 0.21426f
C680 top_segment_1_0.rseg_1_v3_1.v41 top_segment_1_0.rseg_1_v3_1.v44 0.02715f
C681 VH2 top_segment_2_0.DEC2[0] 0.20764f
C682 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.30979f
C683 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.02015f
C684 top_segment_1_0.rseg_1_v3_1.v42 top_segment_1_0.rseg_1_v3_1.v43 1.34308f
C685 top_segment_3_0.bb[6] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.06259f
C686 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC1[3] 0.57206f
C687 DIN7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.01582f
C688 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC2[0] 0.06788f
C689 SH[3] top_segment_4_1.bb3 0.09763f
C690 SH[4] top_segment_4_1.b3 0.09664f
C691 top_segment_1_0.rseg_1_v3_1.v19 top_segment_1_0.rseg_1_v3_1.v23 0.05244f
C692 top_segment_1_0.rseg_1_v3_1.v20 top_segment_1_0.rseg_1_v3_1.v22 1.68068f
C693 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v42 0.17921f
C694 SH[4] top_segment_2_0.DEC2[3] 0.05175f
C695 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_40454_21045# 0.02974f
C696 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_4_1.b3 0.06291f
C697 top_segment_2_0.V0 SH[4] 0.11409f
C698 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.4555f
C699 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_3_0.bb[4] 0.02167f
C700 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 0.01142f
C701 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.06121f
C702 VDDH top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.01105f
C703 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 11.5953f
C704 SH[4] top_segment_2_0.DEC2[1] 0.04851f
C705 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_2_0.DEC2[3] 0.0642f
C706 top_segment_4_1.DEC2 top_segment_4_1.b1 0.06377f
C707 top_segment_2_0.V0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.18985f
C708 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.33918f
C709 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 1.85343f
C710 SH[3] top_segment_4_1.DEC3 0.05175f
C711 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_2_0.DEC2[1] 0.06276f
C712 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 3.83598f
C713 DIN8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.17935f
C714 top_segment_2_0.DEC2[3] top_segment_1_0.rseg_1_v3_1.v60 0.09357f
C715 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_3_0.b[6] 0.01397f
C716 SH[3] top_segment_4_1.DEC1 0.04957f
C717 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC1[1] 0.01814f
C718 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v60 0.25566f
C719 top_segment_1_0.rseg_1_v3_1.v41 top_segment_1_0.rseg_1_v3_1.v43 1.7882f
C720 top_segment_1_0.rseg_1_v3_1.v8 top_segment_1_0.rseg_1_v3_1.v7 0.04824f
C721 top_segment_1_0.rseg_1_v3_1.v9 top_segment_1_0.rseg_1_v3_1.v6 0.04313f
C722 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.14505f
C723 top_segment_1_0.rseg_1_v3_1.v11 top_segment_1_0.rseg_1_v3_1.v4 0.01835f
C724 top_segment_1_0.rseg_1_v3_1.v13 top_segment_1_0.rseg_1_v3_1.v2 0.01887f
C725 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y VDD 0.28031f
C726 top_segment_1_0.rseg_1_v3_1.v50 top_segment_1_0.rseg_1_v3_1.v56 0.0119f
C727 top_segment_1_0.rseg_1_v3_1.v20 top_segment_1_0.rseg_1_v3_1.v21 0.54188f
C728 top_segment_3_0.b[6] top_segment_2_0.DEC0[2] 0.03532f
C729 top_segment_2_0.DEC0[2] top_segment_2_0.DEC1[1] 0.10242f
C730 top_segment_1_0.rseg_1_v3_1.v18 top_segment_1_0.rseg_1_v3_1.v23 0.05838f
C731 top_segment_2_0.DEC1[3] top_segment_3_0.bb[5] 0.04361f
C732 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v41 0.16476f
C733 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV VDDH 17.253f
C734 top_segment_3_0.bb[5] top_segment_2_0.DEC2[0] 0.09325f
C735 top_segment_4_1.b2 top_segment_4_1.bb2 15.3143f
C736 SH[1] top_segment_4_1.bb3 0.12741f
C737 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_3_0.b[4] 0.05817f
C738 VDD DIN6 0.70858f
C739 top_segment_2_0.DEC1[3] top_segment_4_1.bb3 0.04843f
C740 top_segment_4_1.bb3 top_segment_2_0.DEC2[0] 0.09787f
C741 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.11006f
C742 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.0942f
C743 top_segment_2_0.DEC1[2] top_segment_3_0.b[5] 0.04068f
C744 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 1.5609f
C745 top_segment_2_0.DEC2[3] top_segment_1_0.rseg_1_v3_1.v59 0.09964f
C746 VDDH VS4 0.16195f
C747 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.02308f
C748 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v59 0.05743f
C749 SH[2] top_segment_2_0.DEC2[2] 0.04736f
C750 top_segment_2_0.DEC0[1] top_segment_2_0.DEC1[2] 0.33598f
C751 top_segment_3_0.b[6] top_segment_2_0.DEC0[0] 0.03532f
C752 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 1.3157f
C753 top_segment_2_0.DEC0[0] top_segment_2_0.DEC1[1] 0.48656f
C754 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.06014f
C755 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.02715f
C756 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.21475f
C757 a_40454_21045# VDDH 0.31401f
C758 VDDH top_segment_3_0.bb[4] 1.54537f
C759 SH[1] top_segment_4_1.DEC3 0.06246f
C760 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 1.96314f
C761 top_segment_1_0.rseg_1_v3_1.v40 top_segment_1_0.rseg_1_v3_1.v43 0.09811f
C762 top_segment_1_0.rseg_1_v3_1.v41 top_segment_1_0.rseg_1_v3_1.v42 1.32022f
C763 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.02001f
C764 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.30168f
C765 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.02015f
C766 top_segment_1_0.rseg_1_v3_1.v8 top_segment_1_0.rseg_1_v3_1.v6 1.73087f
C767 top_segment_4_1.DEC3 top_segment_2_0.DEC2[0] 15.7968f
C768 SH[1] top_segment_4_1.DEC1 0.0627f
C769 top_segment_1_0.rseg_1_v3_1.v53 top_segment_1_0.rseg_1_v3_1.v44 0.02615f
C770 top_segment_1_0.rseg_1_v3_1.v55 top_segment_1_0.rseg_1_v3_1.v42 1.33973f
C771 top_segment_1_0.rseg_1_v3_1.v51 top_segment_1_0.rseg_1_v3_1.v46 0.02493f
C772 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.02163f
C773 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.14754f
C774 top_segment_4_1.DEC1 top_segment_2_0.DEC2[0] 0.30645f
C775 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.08462f
C776 top_segment_1_0.rseg_1_v3_1.v19 top_segment_1_0.rseg_1_v3_1.v21 1.44458f
C777 top_segment_4_1.bb3 top_segment_4_1.bb1 0.09934f
C778 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v40 0.26016f
C779 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 0.80349f
C780 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.0977f
C781 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.01646f
C782 SH[3] top_segment_4_1.b1 0.09498f
C783 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y VDD 0.41365f
C784 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.06107f
C785 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.48603f
C786 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.48595f
C787 DIN7 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.17937f
C788 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.31886f
C789 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 1.85017f
C790 top_segment_2_0.DEC2[3] top_segment_1_0.rseg_1_v3_1.v58 0.17986f
C791 top_segment_4_1.DEC3 top_segment_4_1.bb1 0.05183f
C792 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC1[0] 0.01617f
C793 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v58 0.18788f
C794 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 0.09454f
C795 top_segment_1_0.rseg_1_v3_1.v40 top_segment_1_0.rseg_1_v3_1.v42 0.55369f
C796 top_segment_4_1.DEC1 top_segment_4_1.bb1 0.04788f
C797 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.06214f
C798 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 0.49734f
C799 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 0.54952f
C800 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B 0.01088f
C801 top_segment_1_0.rseg_1_v3_1.v18 top_segment_1_0.rseg_1_v3_1.v21 0.04809f
C802 top_segment_2_0.DEC0[2] top_segment_2_0.DEC1[0] 0.05224f
C803 top_segment_1_0.rseg_1_v3_1.v19 top_segment_1_0.rseg_1_v3_1.v20 0.54711f
C804 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.21387f
C805 top_segment_2_0.DEC1[2] top_segment_2_0.DEC2[2] 0.05675f
C806 VDDH top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.90751f
C807 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C808 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v7 0.1499f
C809 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C VDD 0.33516f
C810 SH[1] top_segment_4_1.b1 0.12436f
C811 top_segment_2_0.DEC2[3] top_segment_1_0.rseg_1_v3_1.v57 0.16919f
C812 top_segment_2_0.DEC1[1] top_segment_3_0.b[5] 0.04071f
C813 top_segment_3_0.b[6] top_segment_3_0.b[5] 0.21021f
C814 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV a_39072_20445# 0.0755f
C815 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 1.57341f
C816 top_segment_2_0.DEC0[0] top_segment_2_0.DEC1[0] 0.85676f
C817 top_segment_3_0.b[6] top_segment_2_0.DEC0[1] 0.03534f
C818 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v57 0.05667f
C819 top_segment_2_0.DEC0[1] top_segment_2_0.DEC1[1] 0.8597f
C820 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_3_0.bb[5] 0.02352f
C821 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.21451f
C822 top_segment_1_0.rseg_1_v3_1.v40 top_segment_1_0.rseg_1_v3_1.v41 3.81788f
C823 top_segment_2_0.DEC2[0] top_segment_4_1.b1 0.04939f
C824 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 1.34745f
C825 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.02715f
C826 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_4_1.bb3 0.01826f
C827 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.0203f
C828 DIN5 DIN6 0.36448f
C829 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC VDDH 1.19654f
C830 top_segment_1_0.rseg_1_v3_1.v55 top_segment_1_0.rseg_1_v3_1.v40 0.0484f
C831 top_segment_1_0.rseg_1_v3_1.v51 top_segment_1_0.rseg_1_v3_1.v44 0.03397f
C832 top_segment_1_0.rseg_1_v3_1.v53 top_segment_1_0.rseg_1_v3_1.v42 0.02726f
C833 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.22605f
C834 top_segment_1_0.rseg_1_v3_1.v18 top_segment_1_0.rseg_1_v3_1.v20 1.26125f
C835 top_segment_1_0.rseg_1_v3_1.v54 top_segment_1_0.rseg_1_v3_1.v55 0.65418f
C836 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v30 0.02106f
C837 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.04651f
C838 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.14826f
C839 top_segment_3_0.bb[5] top_segment_3_0.bb[4] 0.05167f
C840 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.05001f
C841 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.01649f
C842 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_4_1.DEC3 0.02121f
C843 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 2.59466f
C844 top_segment_4_1.b1 top_segment_4_1.bb1 15.9617f
C845 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.5188f
C846 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.06095f
C847 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v6 0.11835f
C848 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_4_1.DEC1 0.12689f
C849 top_segment_2_0.DEC2[2] top_segment_4_1.b2 0.05451f
C850 DIN8 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.0349f
C851 top_segment_2_0.DEC2[3] top_segment_1_0.rseg_1_v3_1.v56 0.29715f
C852 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.54094f
C853 top_segment_3_0.bb[4] top_segment_4_1.bb3 0.17417f
C854 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v56 0.0944f
C855 top_segment_2_0.DEC0[2] VL2 0.0806f
C856 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.09855f
C857 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 0.20563f
C858 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.02047f
C859 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.02948f
C860 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 0.09239f
C861 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.63972f
C862 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.06351f
C863 top_segment_4_1.DEC3 top_segment_3_0.bb[4] 0.10032f
C864 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 0.5556f
C865 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.01904f
C866 a_39072_20445# VDDH 0.35437f
C867 top_segment_1_0.rseg_1_v3_1.v18 top_segment_1_0.rseg_1_v3_1.v19 0.63647f
C868 top_segment_3_0.b[6] top_segment_2_0.DEC2[2] 0.09106f
C869 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.07187f
C870 top_segment_2_0.DEC1[1] top_segment_2_0.DEC2[2] 0.05322f
C871 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.03773f
C872 top_segment_1_0.rseg_1_v3_1.v53 top_segment_1_0.rseg_1_v3_1.v55 1.97838f
C873 VDDH top_segment_3_0.bb[5] 1.98171f
C874 top_segment_3_0.bb[4] top_segment_4_1.DEC1 0.15269f
C875 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.03404f
C876 top_segment_3_0.bb[6] VH3 0.05139f
C877 top_segment_3_0.bb[6] top_segment_2_0.DEC0[2] 0.05177f
C878 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v5 0.06052f
C879 VDDH top_segment_4_1.bb3 2.86721f
C880 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC2[3] 0.03409f
C881 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC2[1] 0.03991f
C882 top_segment_2_0.DEC1[0] top_segment_3_0.b[5] 0.04075f
C883 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.0119f
C884 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.28212f
C885 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 1.57642f
C886 top_segment_2_0.DEC0[1] top_segment_2_0.DEC1[0] 0.10571f
C887 VDD DIN4 0.67214f
C888 top_segment_2_0.DEC0[2] top_segment_4_1.b3 0.04799f
C889 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 1.60464f
C890 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 1.3734f
C891 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 0.21361f
C892 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 0.02715f
C893 VH3 top_segment_4_1.b3 0.16841f
C894 top_segment_1_0.rseg_1_v3_1.v8 top_segment_1_0.rseg_1_v3_1.v2 0.0119f
C895 VDDH top_segment_4_1.DEC3 3.72487f
C896 top_segment_2_0.DEC0[2] top_segment_2_0.DEC2[3] 0.06841f
C897 top_segment_2_0.V0 top_segment_2_0.DEC0[2] 0.11848f
C898 top_segment_3_0.bb[6] top_segment_2_0.DEC0[0] 0.05177f
C899 VDDH top_segment_4_1.DEC1 3.65941f
C900 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 0.16825f
C901 top_segment_2_0.DEC0[2] top_segment_2_0.DEC2[1] 0.10148f
C902 top_segment_1_0.rseg_1_v3_1.v53 top_segment_1_0.rseg_1_v3_1.v54 0.48841f
C903 top_segment_1_0.rseg_1_v3_1.v52 top_segment_1_0.rseg_1_v3_1.v55 0.06115f
C904 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.21507f
C905 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.56698f
C906 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 VDDH 2.01261f
C907 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.04706f
C908 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y 0.15447f
C909 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_38430_18467# 0.02736f
C910 top_segment_2_0.DEC0[0] top_segment_4_1.b3 0.04799f
C911 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.01651f
C912 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v4 0.03958f
C913 top_segment_2_0.DEC0[0] top_segment_2_0.DEC2[3] 0.05159f
C914 top_segment_4_1.b3 top_segment_4_1.bb2 0.11077f
C915 top_segment_2_0.DEC2[3] top_segment_1_0.rseg_1_v3_1.v46 0.02186f
C916 top_segment_2_0.V0 top_segment_2_0.DEC0[0] 0.25426f
C917 top_segment_2_0.DEC0[0] top_segment_2_0.DEC2[1] 0.04839f
C918 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.19158f
C919 top_segment_2_0.DEC2[3] top_segment_4_1.bb2 0.05183f
C920 SH[2] top_segment_4_1.b2 0.09759f
C921 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v46 0.10302f
C922 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.50346f
C923 top_segment_2_0.V0 top_segment_4_1.bb2 0.15088f
C924 top_segment_2_0.DEC0[2] top_segment_3_0.b[4] 0.04324f
C925 top_segment_2_0.DEC2[1] top_segment_4_1.bb2 0.0486f
C926 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.01808f
C927 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.6765f
C928 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.02906f
C929 top_segment_2_0.DEC1[0] top_segment_2_0.DEC2[2] 0.05891f
C930 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.5557f
C931 top_segment_1_0.rseg_1_v3_1.v51 top_segment_1_0.rseg_1_v3_1.v55 0.05244f
C932 top_segment_1_0.rseg_1_v3_1.v52 top_segment_1_0.rseg_1_v3_1.v54 1.63811f
C933 a_43562_3816# top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.02963f
C934 DIN9 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.17935f
C935 VDDH top_segment_1_0.rseg_1_v3_1.v7 0.02285f
C936 top_segment_2_0.DEC0[0] top_segment_3_0.b[4] 0.04328f
C937 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v3 0.03915f
C938 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC 0.12736f
C939 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.03009f
C940 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A VDD 0.59039f
C941 VDDH top_segment_4_1.b1 1.08229f
C942 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v45 0.0759f
C943 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 0.0119f
C944 SH[4] top_segment_4_1.DEC2 0.05178f
C945 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 1.57251f
C946 a_43562_3816# top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y 0.02202f
C947 top_segment_3_0.bb[6] top_segment_3_0.b[5] 15.2414f
C948 top_segment_3_0.bb[5] top_segment_4_1.bb3 0.05478f
C949 top_segment_3_0.bb[6] top_segment_2_0.DEC0[1] 0.05179f
C950 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.2354f
C951 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v26 0.01144f
C952 top_segment_1_0.rseg_1_v3_1.v50 top_segment_1_0.rseg_1_v3_1.v55 0.05769f
C953 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C954 top_segment_1_0.rseg_1_v3_1.v52 top_segment_1_0.rseg_1_v3_1.v53 0.60003f
C955 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.22406f
C956 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 0.16949f
C957 top_segment_3_0.b[5] top_segment_4_1.b3 0.05424f
C958 DIN4 DIN5 0.34355f
C959 top_segment_2_0.DEC2[3] top_segment_3_0.b[5] 0.09256f
C960 top_segment_2_0.DEC0[1] top_segment_4_1.b3 0.04799f
C961 VL3 VH3 0.25091f
C962 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B 0.77374f
C963 top_segment_4_1.DEC3 top_segment_3_0.bb[5] 0.09577f
C964 top_segment_2_0.V0 top_segment_3_0.b[5] 0.11409f
C965 top_segment_2_0.DEC2[0] top_segment_1_0.rseg_1_v3_1.v2 0.06158f
C966 top_segment_3_0.b[5] top_segment_2_0.DEC2[1] 0.09024f
C967 top_segment_2_0.DEC0[1] top_segment_2_0.DEC2[3] 0.0505f
C968 top_segment_2_0.V0 top_segment_2_0.DEC0[1] 0.11848f
C969 top_segment_3_0.bb[5] top_segment_4_1.DEC1 0.09063f
C970 top_segment_4_1.DEC3 top_segment_4_1.bb3 0.24407f
C971 top_segment_2_0.DEC0[1] top_segment_2_0.DEC2[1] 0.0483f
C972 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v44 0.07383f
C973 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.05086f
C974 VL2 top_segment_2_0.DEC2[2] 0.23574f
C975 top_segment_3_0.b[6] top_segment_2_0.DEC1[2] 0.03539f
C976 top_segment_2_0.DEC1[1] top_segment_2_0.DEC1[2] 17.521f
C977 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.14301f
C978 top_segment_4_1.bb3 top_segment_4_1.DEC1 0.09642f
C979 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.02775f
C980 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 0.03397f
C981 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.0672f
C982 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.69667f
C983 top_segment_1_0.rseg_1_v3_1.v51 top_segment_1_0.rseg_1_v3_1.v53 1.45197f
C984 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.13531f
C985 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 0.55111f
C986 top_segment_4_1.DEC3 top_segment_4_1.DEC1 0.06201f
C987 VDDH DIN3 0.42749f
C988 top_segment_3_0.b[5] top_segment_3_0.b[4] 1.24741f
C989 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.15687f
C990 top_segment_2_0.DEC0[1] top_segment_3_0.b[4] 0.0433f
C991 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.02077f
C992 top_segment_3_0.bb[6] top_segment_2_0.DEC2[2] 0.10104f
C993 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.11246f
C994 SH[4] SH[3] 17.4953f
C995 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC ROUT 0.01108f
C996 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.20262f
C997 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v43 0.05973f
C998 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.11989f
C999 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.0119f
C1000 top_segment_1_0.rseg_1_v3_1.v29 top_segment_1_0.rseg_1_v3_1.v30 1.19856f
C1001 a_38408_21484# ROUT 0.13835f
C1002 top_segment_4_1.b3 top_segment_2_0.DEC2[2] 0.09997f
C1003 top_segment_2_0.DEC2[3] top_segment_2_0.DEC2[2] 17.2409f
C1004 top_segment_2_0.V0 top_segment_2_0.DEC2[2] 1.88678f
C1005 top_segment_2_0.DEC2[2] top_segment_2_0.DEC2[1] 17.4112f
C1006 top_segment_1_0.rseg_1_v3_1.v51 top_segment_1_0.rseg_1_v3_1.v52 0.60342f
C1007 top_segment_1_0.rseg_1_v3_1.v50 top_segment_1_0.rseg_1_v3_1.v53 0.04864f
C1008 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 0.13705f
C1009 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 1.57937f
C1010 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 3.55677f
C1011 top_segment_4_1.bb3 top_segment_4_1.b1 0.10583f
C1012 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.18669f
C1013 top_segment_2_0.DEC2[3] top_segment_1_0.rseg_1_v3_1.v42 0.01149f
C1014 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.06435f
C1015 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v42 0.04946f
C1016 top_segment_1_0.rseg_1_v3_1.v28 top_segment_1_0.rseg_1_v3_1.v30 1.1572f
C1017 top_segment_2_0.DEC1[0] top_segment_2_0.DEC1[2] 0.68733f
C1018 top_segment_3_0.b[6] top_segment_2_0.DEC1[1] 0.03545f
C1019 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.01469f
C1020 top_segment_3_0.b[4] top_segment_2_0.DEC2[2] 0.09076f
C1021 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.14057f
C1022 top_segment_4_1.DEC3 top_segment_4_1.b1 0.05185f
C1023 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 1.15198f
C1024 SH[4] top_segment_2_0.DEC2[0] 0.04929f
C1025 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.3076f
C1026 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.03419f
C1027 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.06886f
C1028 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.02748f
C1029 top_segment_4_1.DEC1 top_segment_4_1.b1 0.04789f
C1030 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_2_0.DEC1[3] 0.70899f
C1031 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_2_0.DEC2[0] 0.06345f
C1032 top_segment_1_0.rseg_1_v3_1.v50 top_segment_1_0.rseg_1_v3_1.v52 1.21429f
C1033 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 0.71512f
C1034 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.05086f
C1035 DIN8 DIN9 0.33674f
C1036 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 1.24591f
C1037 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 0.11236f
C1038 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.02181f
C1039 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C VDD 0.26024f
C1040 SH[4] top_segment_4_1.bb1 0.09685f
C1041 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v41 0.06043f
C1042 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.82681f
C1043 top_segment_1_0.rseg_1_v3_1.v55 top_segment_2_0.DEC2[3] 0.15103f
C1044 top_segment_1_0.rseg_1_v3_1.v28 top_segment_1_0.rseg_1_v3_1.v29 1.19056f
C1045 top_segment_1_0.rseg_1_v3_1.v27 top_segment_1_0.rseg_1_v3_1.v30 0.0119f
C1046 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 0.0119f
C1047 top_segment_1_0.rseg_1_v3_1.v55 top_segment_2_0.V0 0.03652f
C1048 SH[2] top_segment_4_1.b3 0.09657f
C1049 VDDH top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.01029f
C1050 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.2275f
C1051 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.15123f
C1052 top_segment_1_0.rseg_1_v3_1.v45 top_segment_1_0.rseg_1_v3_1.v38 0.02015f
C1053 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 0.04651f
C1054 SH[2] top_segment_2_0.DEC2[3] 0.05186f
C1055 top_segment_2_0.V0 SH[2] 0.11409f
C1056 top_segment_1_0.rseg_1_v3_1.v50 top_segment_1_0.rseg_1_v3_1.v51 0.69962f
C1057 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC0[2] 0.24881f
C1058 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.11902f
C1059 SH[2] top_segment_2_0.DEC2[1] 0.04851f
C1060 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.01138f
C1061 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 ROUT 0.01358f
C1062 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.01056f
C1063 a_43284_3816# VDD 0.02571f
C1064 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.0191f
C1065 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.48049f
C1066 VDD DIN9 0.75623f
C1067 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v40 0.09994f
C1068 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.26572f
C1069 top_segment_3_0.b[6] top_segment_2_0.DEC1[0] 0.03552f
C1070 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.09312f
C1071 top_segment_1_0.rseg_1_v3_1.v27 top_segment_1_0.rseg_1_v3_1.v29 1.72824f
C1072 top_segment_2_0.DEC1[0] top_segment_2_0.DEC1[1] 17.3149f
C1073 top_segment_1_0.rseg_1_v3_1.v26 top_segment_1_0.rseg_1_v3_1.v30 0.36625f
C1074 top_segment_1_0.rseg_1_v3_1.v54 top_segment_2_0.DEC2[3] 0.09709f
C1075 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC0[0] 0.44826f
C1076 top_segment_1_0.rseg_1_v3_1.v54 top_segment_2_0.V0 0.05551f
C1077 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 2.1375f
C1078 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 0.33162f
C1079 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_4_1.DEC2 0.02213f
C1080 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C 0.2455f
C1081 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 11.8244f
C1082 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 0.0119f
C1083 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 1.18866f
C1084 DIN0 DIN1 0.32901f
C1085 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 0.03375f
C1086 top_segment_3_0.bb[6] top_segment_2_0.DEC1[2] 0.05169f
C1087 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.02726f
C1088 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.06862f
C1089 top_segment_1_0.rseg_1_v3_1.v6 top_segment_1_0.rseg_1_v3_1.v7 0.55841f
C1090 a_42614_21484# ROUT 0.08397f
C1091 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.03966f
C1092 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.06435f
C1093 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v39 0.15057f
C1094 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.21864f
C1095 VDD DIN1 0.66672f
C1096 top_segment_2_0.DEC1[2] top_segment_4_1.b3 0.04806f
C1097 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 0.05213f
C1098 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 0.02116f
C1099 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.06069f
C1100 top_segment_2_0.DEC1[2] top_segment_2_0.DEC2[3] 0.1111f
C1101 top_segment_2_0.V0 top_segment_2_0.DEC1[2] 0.11848f
C1102 top_segment_2_0.DEC1[2] top_segment_2_0.DEC2[1] 0.09914f
C1103 top_segment_1_0.rseg_1_v3_1.v27 top_segment_1_0.rseg_1_v3_1.v28 1.31906f
C1104 top_segment_1_0.rseg_1_v3_1.v53 top_segment_2_0.DEC2[3] 0.06038f
C1105 top_segment_1_0.rseg_1_v3_1.v26 top_segment_1_0.rseg_1_v3_1.v29 0.0954f
C1106 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.24855f
C1107 top_segment_1_0.rseg_1_v3_1.v53 top_segment_2_0.V0 0.04346f
C1108 top_segment_1_0.rseg_1_v3_1.v45 top_segment_1_0.rseg_1_v3_1.v36 0.02194f
C1109 top_segment_1_0.rseg_1_v3_1.v43 top_segment_1_0.rseg_1_v3_1.v38 0.05318f
C1110 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 1.31557f
C1111 top_segment_4_1.DEC2 top_segment_4_1.bb2 0.07184f
C1112 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B VDD 0.29366f
C1113 top_segment_1_0.rseg_1_v3_1.v5 top_segment_1_0.rseg_1_v3_1.v7 1.9603f
C1114 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 0.04533f
C1115 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B 0.28615f
C1116 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 2.29207f
C1117 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 0.0847f
C1118 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_3_0.bb[4] 0.06334f
C1119 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v38 0.09809f
C1120 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 0.0921f
C1121 top_segment_2_0.DEC1[2] top_segment_3_0.b[4] 0.04329f
C1122 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.08478f
C1123 a_43018_3816# top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.01759f
C1124 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.21776f
C1125 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v30 0.15598f
C1126 top_segment_1_0.rseg_1_v3_1.v52 top_segment_2_0.DEC2[3] 0.03202f
C1127 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC0[1] 0.30079f
C1128 top_segment_1_0.rseg_1_v3_1.v25 top_segment_1_0.rseg_1_v3_1.v29 0.08427f
C1129 SH[2] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A 0.1676f
C1130 top_segment_1_0.rseg_1_v3_1.v26 top_segment_1_0.rseg_1_v3_1.v28 1.94958f
C1131 top_segment_4_1.b3 top_segment_4_1.b2 0.22613f
C1132 top_segment_1_0.rseg_1_v3_1.v52 top_segment_2_0.V0 0.07007f
C1133 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 2.15445f
C1134 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 0.36689f
C1135 VDDH SH[4] 0.68463f
C1136 top_segment_2_0.DEC2[3] top_segment_4_1.b2 0.0532f
C1137 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 0.0119f
C1138 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 1.21733f
C1139 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 1.81308f
C1140 top_segment_3_0.bb[6] top_segment_2_0.DEC1[1] 0.0517f
C1141 top_segment_1_0.rseg_1_v3_1.v5 top_segment_1_0.rseg_1_v3_1.v6 0.39192f
C1142 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.13356f
C1143 top_segment_3_0.b[6] top_segment_3_0.bb[6] 16.6023f
C1144 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] VDDH 2.1111f
C1145 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC a_37131_19377# 0.02882f
C1146 top_segment_1_0.rseg_1_v3_1.v4 top_segment_1_0.rseg_1_v3_1.v7 0.05585f
C1147 top_segment_2_0.V0 top_segment_4_1.b2 0.11409f
C1148 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.48636f
C1149 top_segment_2_0.DEC2[1] top_segment_4_1.b2 0.04862f
C1150 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.13195f
C1151 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v37 0.06065f
C1152 top_segment_2_0.DEC1[1] top_segment_4_1.b3 0.04807f
C1153 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 10.3939f
C1154 top_segment_3_0.b[6] top_segment_4_1.b3 0.04999f
C1155 VDDH DIN7 0.42767f
C1156 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.02213f
C1157 top_segment_3_0.b[6] top_segment_2_0.DEC2[3] 0.09163f
C1158 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 0.05322f
C1159 top_segment_2_0.DEC1[1] top_segment_2_0.DEC2[3] 0.11775f
C1160 top_segment_2_0.V0 top_segment_2_0.DEC1[1] 0.11848f
C1161 top_segment_2_0.V0 top_segment_3_0.b[6] 0.11409f
C1162 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B 0.13753f
C1163 top_segment_3_0.b[6] top_segment_2_0.DEC2[1] 0.09344f
C1164 top_segment_2_0.DEC1[1] top_segment_2_0.DEC2[1] 0.05719f
C1165 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v29 0.17836f
C1166 top_segment_1_0.rseg_1_v3_1.v26 top_segment_1_0.rseg_1_v3_1.v27 1.31057f
C1167 top_segment_1_0.rseg_1_v3_1.v51 top_segment_2_0.DEC2[3] 0.03135f
C1168 top_segment_1_0.rseg_1_v3_1.v25 top_segment_1_0.rseg_1_v3_1.v28 0.02715f
C1169 top_segment_1_0.rseg_1_v3_1.v24 top_segment_1_0.rseg_1_v3_1.v29 0.21425f
C1170 top_segment_3_0.b[5] top_segment_4_1.DEC2 0.09326f
C1171 top_segment_1_0.rseg_1_v3_1.v51 top_segment_2_0.V0 0.0658f
C1172 SH[3] top_segment_4_1.bb2 0.09789f
C1173 top_segment_1_0.rseg_1_v3_1.v45 top_segment_1_0.rseg_1_v3_1.v34 0.02179f
C1174 top_segment_1_0.rseg_1_v3_1.v43 top_segment_1_0.rseg_1_v3_1.v36 0.02214f
C1175 top_segment_1_0.rseg_1_v3_1.v40 top_segment_1_0.rseg_1_v3_1.v39 0.14454f
C1176 top_segment_1_0.rseg_1_v3_1.v41 top_segment_1_0.rseg_1_v3_1.v38 0.04748f
C1177 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A 0.10895f
C1178 top_segment_1_0.rseg_1_v3_1.v4 top_segment_1_0.rseg_1_v3_1.v6 1.8445f
C1179 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC1[3] 0.01796f
C1180 top_segment_1_0.rseg_1_v3_1.v3 top_segment_1_0.rseg_1_v3_1.v7 0.05245f
C1181 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.16165f
C1182 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.1481f
C1183 VDDH DIN8 0.4277f
C1184 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 0.05787f
C1185 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_segment_2_0.DEC2[0] 0.04948f
C1186 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.53572f
C1187 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC2[2] 0.19276f
C1188 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] 0.21309f
C1189 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 2.14311f
C1190 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 0.08427f
C1191 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v36 0.03176f
C1192 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.02488f
C1193 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV ROUT 0.25958f
C1194 top_segment_3_0.b[6] top_segment_3_0.b[4] 0.08389f
C1195 top_segment_2_0.DEC1[1] top_segment_3_0.b[4] 0.0433f
C1196 top_segment_2_0.DEC0[2] top_segment_2_0.DEC1[3] 0.26998f
C1197 top_segment_2_0.DEC0[2] top_segment_2_0.DEC2[0] 0.05872f
C1198 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.07378f
C1199 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v28 0.09131f
C1200 top_segment_1_0.rseg_1_v3_1.v50 top_segment_2_0.DEC2[3] 0.06054f
C1201 top_segment_1_0.rseg_1_v3_1.v25 top_segment_1_0.rseg_1_v3_1.v27 1.789f
C1202 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y VDD 0.33964f
C1203 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 0.09271f
C1204 top_segment_1_0.rseg_1_v3_1.v50 top_segment_2_0.V0 0.158f
C1205 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.10418f
C1206 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 1.93547f
C1207 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 2.90337f
C1208 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 2.15145f
C1209 VDDH DIN0 0.4291f
C1210 top_segment_1_0.rseg_1_v3_1.v40 top_segment_1_0.rseg_1_v3_1.v38 1.73225f
C1211 top_segment_3_0.bb[6] top_segment_2_0.DEC1[0] 0.05174f
C1212 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 0.0119f
C1213 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 1.24994f
C1214 top_segment_1_0.rseg_1_v3_1.v4 top_segment_1_0.rseg_1_v3_1.v5 0.50407f
C1215 top_segment_1_0.rseg_1_v3_1.v2 top_segment_1_0.rseg_1_v3_1.v7 0.0555f
C1216 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.0483f
C1217 top_segment_2_0.DEC0[0] top_segment_2_0.DEC1[3] 16.1091f
C1218 SH[1] top_segment_4_1.bb2 0.12766f
C1219 top_segment_2_0.DEC0[0] top_segment_2_0.DEC2[0] 0.04891f
C1220 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 0.1869f
C1221 VDDH top_segment_1_0.rseg_1_v3_1.v58 0.15493f
C1222 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.13341f
C1223 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.09312f
C1224 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v35 0.03135f
C1225 VDDH VDD 5.2366f
C1226 top_segment_2_0.DEC2[0] top_segment_4_1.bb2 0.0494f
C1227 top_segment_2_0.DEC2[2] top_segment_4_1.DEC2 0.55748f
C1228 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 0.41945f
C1229 top_segment_2_0.DEC1[0] top_segment_4_1.b3 0.04809f
C1230 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 1.26639f
C1231 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 0.10213f
C1232 top_segment_2_0.DEC1[0] top_segment_2_0.DEC2[3] 16.2949f
C1233 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_3_0.bb[5] 0.05842f
C1234 SH[4] top_segment_4_1.bb3 0.09769f
C1235 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 0.05305f
C1236 top_segment_2_0.V0 top_segment_2_0.DEC1[0] 0.11848f
C1237 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 0.02197f
C1238 top_segment_1_0.rseg_1_v3_1.v25 top_segment_1_0.rseg_1_v3_1.v26 1.29067f
C1239 top_segment_1_0.rseg_1_v3_1.v24 top_segment_1_0.rseg_1_v3_1.v27 0.09809f
C1240 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v27 0.09136f
C1241 top_segment_2_0.DEC1[0] top_segment_2_0.DEC2[1] 0.05223f
C1242 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] top_segment_4_1.bb3 0.06335f
C1243 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] a_43890_3816# 0.01631f
C1244 VDDH ROUT 9.92565f
C1245 top_segment_1_0.rseg_1_v3_1.v30 top_segment_1_0.rseg_1_v3_1.v39 0.01647f
C1246 top_segment_4_1.bb2 top_segment_4_1.bb1 0.31324f
C1247 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC 0.35106f
C1248 top_segment_1_0.rseg_1_v3_1.v3 top_segment_1_0.rseg_1_v3_1.v5 1.41253f
C1249 SH[4] top_segment_4_1.DEC3 0.05177f
C1250 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 0.05772f
C1251 SH[4] top_segment_4_1.DEC1 0.0478f
C1252 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 0.57187f
C1253 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y 0.10297f
C1254 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] 2.8803f
C1255 top_segment_2_0.DEC2[2] top_segment_1_0.rseg_1_v3_1.v34 0.06082f
C1256 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 2.09546f
C1257 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.08427f
C1258 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] 0.0421f
C1259 top_segment_2_0.DEC1[0] top_segment_3_0.b[4] 0.04333f
C1260 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 2.73645f
C1261 top_segment_2_0.V0 top_segment_1_0.rseg_1_v3_1.v26 0.01034f
C1262 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] 0.19767f
C1263 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v26 0.17853f
C1264 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.07f
C1265 top_segment_1_0.rseg_1_v3_1.v24 top_segment_1_0.rseg_1_v3_1.v26 0.55643f
C1266 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 1.94253f
C1267 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.06751f
C1268 top_segment_2_0.DEC1[3] top_segment_3_0.b[5] 0.04066f
C1269 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.01119f
C1270 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y 0.08193f
C1271 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 2.15109f
C1272 top_segment_1_0.rseg_1_v3_1.v3 top_segment_1_0.rseg_1_v3_1.v4 0.51079f
C1273 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC0[2] 0.02388f
C1274 top_segment_1_0.rseg_1_v3_1.v2 top_segment_1_0.rseg_1_v3_1.v5 0.0481f
C1275 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 0.20641f
C1276 top_segment_3_0.b[5] top_segment_2_0.DEC2[0] 0.09038f
C1277 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.2275f
C1278 top_segment_2_0.DEC0[1] top_segment_2_0.DEC1[3] 0.33061f
C1279 VL2 top_segment_2_0.DEC2[3] 0.14343f
C1280 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.01753f
C1281 top_segment_2_0.DEC0[1] top_segment_2_0.DEC2[0] 0.04883f
C1282 SH[3] top_segment_2_0.DEC2[2] 0.04736f
C1283 VDDH top_segment_1_0.rseg_1_v3_1.v56 0.10984f
C1284 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV a_38430_18842# 0.02806f
C1285 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y 0.0673f
C1286 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.17953f
C1287 VL2 top_segment_2_0.DEC2[1] 0.12679f
C1288 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.05433f
C1289 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 0.15152f
C1290 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 0.03011f
C1291 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 1.36438f
C1292 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 0.18775f
C1293 SH[2] top_segment_4_1.DEC2 0.05175f
C1294 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 0.10119f
C1295 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 1.3027f
C1296 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.05434f
C1297 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC0[0] 0.02124f
C1298 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 0.02197f
C1299 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 0.05322f
C1300 top_segment_3_0.bb[6] top_segment_4_1.b3 0.1857f
C1301 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v25 0.15742f
C1302 top_segment_2_0.DEC0[2] top_segment_3_0.bb[4] 0.04841f
C1303 top_segment_1_0.rseg_1_v3_1.v24 top_segment_1_0.rseg_1_v3_1.v25 3.7974f
C1304 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] 0.21283f
C1305 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.17741f
C1306 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_4_1.bb2 0.01812f
C1307 top_segment_3_0.bb[6] top_segment_2_0.DEC2[3] 0.10422f
C1308 VDDH DIN5 0.42749f
C1309 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.01851f
C1310 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC1[2] 0.30111f
C1311 top_segment_2_0.V0 top_segment_3_0.bb[6] 0.11409f
C1312 SH[4] top_segment_4_1.b1 0.09554f
C1313 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 0.05833f
C1314 top_segment_3_0.bb[6] top_segment_2_0.DEC2[1] 0.10358f
C1315 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 0.11563f
C1316 top_segment_1_0.rseg_1_v3_1.v2 top_segment_1_0.rseg_1_v3_1.v4 1.40088f
C1317 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV VDDH 1.06415f
C1318 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.24146f
C1319 top_segment_4_1.DEC2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 0.17101f
C1320 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.36098f
C1321 top_segment_2_0.DEC2[3] top_segment_4_1.b3 0.20079f
C1322 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 0.05765f
C1323 top_segment_2_0.DEC0[0] top_segment_3_0.bb[4] 0.04845f
C1324 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C 0.01642f
C1325 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.59731f
C1326 top_segment_2_0.V0 top_segment_4_1.b3 0.11409f
C1327 top_segment_4_1.b3 top_segment_2_0.DEC2[1] 0.09743f
C1328 top_segment_2_0.V0 top_segment_2_0.DEC2[3] 0.13293f
C1329 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 2.07729f
C1330 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 0.08427f
C1331 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 0.01346f
C1332 top_segment_2_0.DEC2[3] top_segment_2_0.DEC2[1] 0.56233f
C1333 SH[1] top_segment_2_0.DEC2[2] 0.05806f
C1334 top_segment_2_0.DEC0[2] VDDH 0.99488f
C1335 top_segment_2_0.V0 top_segment_2_0.DEC2[1] 0.13739f
C1336 top_segment_2_0.DEC1[3] top_segment_2_0.DEC2[2] 0.09461f
C1337 VDDH VH3 0.16466f
C1338 top_segment_4_1.DEC3 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 0.1877f
C1339 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC a_37131_19653# 0.02697f
C1340 top_segment_2_0.DEC2[2] top_segment_2_0.DEC2[0] 0.73748f
C1341 DIN6 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.01584f
C1342 top_segment_2_0.DEC2[1] top_segment_1_0.rseg_1_v3_1.v24 0.20729f
C1343 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 0.80785f
C1344 top_segment_3_0.bb[6] top_segment_3_0.b[4] 0.05996f
C1345 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A 0.10925f
C1346 top_segment_1_0.rseg_1_v3_1.v40 top_segment_1_0.rseg_1_v3_1.v34 0.0119f
C1347 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 1.95068f
C1348 top_segment_1_0.rseg_1_v3_1.v2 top_segment_1_0.rseg_1_v3_1.v3 0.59845f
C1349 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.12526f
C1350 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] 3.15778f
C1351 top_segment_2_0.DEC0[0] VDDH 1.07221f
C1352 top_segment_3_0.b[4] top_segment_4_1.b3 0.15163f
C1353 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] 0.1906f
C1354 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.20918f
C1355 top_segment_2_0.DEC2[3] top_segment_3_0.b[4] 0.09513f
C1356 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV 2.49981f
C1357 VDDH top_segment_4_1.bb2 1.55711f
C1358 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.04783f
C1359 SH[3] SH[2] 18.6008f
C1360 VDD top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y 0.2275f
C1361 top_segment_2_0.V0 top_segment_3_0.b[4] 0.11409f
C1362 top_segment_2_0.DEC2[2] top_segment_4_1.bb1 0.05983f
C1363 top_segment_3_0.b[4] top_segment_2_0.DEC2[1] 0.09271f
C1364 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] 0.0184f
C1365 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.05681f
C1366 a_38408_21045# top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV 0.03219f
C1367 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.04792f
C1368 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 ROUT 0.0484f
C1369 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_3_0.b[5] 0.01172f
C1370 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 1.3376f
C1371 top_segment_2_0.DEC0[2] VH2 0.07283f
C1372 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV top_segment_2_0.DEC0[1] 0.02339f
C1373 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 0.10107f
C1374 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] 0.18515f
C1375 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 1.33058f
C1376 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC0[2] 0.16626f
C1377 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC top_segment_2_0.DEC1[1] 0.28795f
C1378 top_segment_1_0.rseg_1_v3_1.v28 top_segment_1_0.rseg_1_v3_1.v37 0.02611f
C1379 top_segment_1_0.rseg_1_v3_1.v30 top_segment_1_0.rseg_1_v3_1.v35 0.02537f
C1380 top_segment_1_0.rseg_1_v3_1.v26 top_segment_1_0.rseg_1_v3_1.v39 1.34056f
C1381 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 top_segment_1_0.rseg_1_v3_1.v7 0.20097f
C1382 VDDH top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 0.0706f
C1383 top_segment_4_1.DEC1 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 0.05995f
C1384 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y 0.07189f
C1385 top_segment_3_0.b[5] top_segment_3_0.bb[4] 0.0497f
C1386 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A VDD 0.33616f
C1387 top_segment_3_0.bb[6] VL3 0.04899f
C1388 top_segment_2_0.DEC0[1] top_segment_3_0.bb[4] 0.04841f
C1389 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC top_segment_2_0.DEC0[0] 0.19453f
C1390 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 0.05759f
C1391 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 0.61579f
C1392 top_segment_4_1.DEC2 top_segment_4_1.b2 0.22616f
C1393 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y 0.06351f
C1394 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] 10.4407f
C1395 SH[1] GND 26.75718f
C1396 SH[2] GND 39.47077f
C1397 DIN9 GND 2.58682f
C1398 DIN8 GND 2.24158f
C1399 SH[3] GND 37.52045f
C1400 DIN7 GND 2.21448f
C1401 DIN6 GND 2.18502f
C1402 SH[4] GND 34.58608f
C1403 VS1 GND 0.29156f
C1404 VS4 GND 0.10631f
C1405 DIN5 GND 2.16664f
C1406 DIN4 GND 2.15816f
C1407 DIN3 GND 2.13965f
C1408 DIN2 GND 2.11716f
C1409 DIN1 GND 2.1019f
C1410 DIN0 GND 2.34399f
C1411 VL2 GND 0.45135f
C1412 VH2 GND 0.6129f
C1413 VH3 GND 0.11819f
C1414 VL3 GND 0.05336f
C1415 ROUT GND 14.28184f
C1416 VDD GND 0.15655p
C1417 VDDH GND 0.35579p
C1418 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.B GND 0.39231f
C1419 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.Y GND 0.3768f
C1420 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.A GND 0.68099f
C1421 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x6.Y GND 0.70838f
C1422 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.C GND 0.3332f
C1423 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.B GND 0.32574f
C1424 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.B GND 0.31137f
C1425 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.A GND 0.25769f
C1426 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x4.A GND 0.32968f
C1427 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.Y GND 0.45293f
C1428 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.C GND 0.41678f
C1429 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.B GND 0.42992f
C1430 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.Y GND 0.33977f
C1431 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x4.A GND 0.73456f
C1432 a_43890_3816# GND 0.02142f $ **FLOATING
C1433 a_43018_3816# GND 0.02172f $ **FLOATING
C1434 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.B GND 0.44413f
C1435 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x3.A GND 0.49956f
C1436 top_segment_1_0.rseg_1_v3_1.v55 GND 1.58565f
C1437 top_segment_1_0.rseg_1_v3_1.v54 GND 1.01698f
C1438 top_segment_1_0.rseg_1_v3_1.v53 GND 0.83396f
C1439 top_segment_1_0.rseg_1_v3_1.v52 GND 0.84338f
C1440 top_segment_1_0.rseg_1_v3_1.v51 GND 0.72928f
C1441 top_segment_1_0.rseg_1_v3_1.v50 GND 0.81839f
C1442 top_segment_1_0.rseg_1_v3_1.v39 GND 1.60815f
C1443 top_segment_1_0.rseg_1_v3_1.v38 GND 1.05072f
C1444 top_segment_1_0.rseg_1_v3_1.v37 GND 0.85279f
C1445 top_segment_1_0.rseg_1_v3_1.v36 GND 0.85992f
C1446 top_segment_1_0.rseg_1_v3_1.v35 GND 0.74171f
C1447 top_segment_1_0.rseg_1_v3_1.v34 GND 0.83636f
C1448 top_segment_1_0.rseg_1_v3_1.v23 GND 1.64361f
C1449 top_segment_1_0.rseg_1_v3_1.v22 GND 1.10159f
C1450 top_segment_1_0.rseg_1_v3_1.v21 GND 0.88377f
C1451 top_segment_1_0.rseg_1_v3_1.v20 GND 0.74063f
C1452 top_segment_1_0.rseg_1_v3_1.v19 GND 0.77336f
C1453 top_segment_1_0.rseg_1_v3_1.v18 GND 0.88264f
C1454 top_segment_1_0.rseg_1_v3_1.v7 GND 2.61761f
C1455 top_segment_1_0.rseg_1_v3_1.v6 GND 1.84052f
C1456 top_segment_1_0.rseg_1_v3_1.v5 GND 1.36319f
C1457 top_segment_1_0.rseg_1_v3_1.v4 GND 1.54449f
C1458 top_segment_1_0.rseg_1_v3_1.v3 GND 1.34744f
C1459 top_segment_1_0.rseg_1_v3_1.v2 GND 2.56072f
C1460 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55 GND 1.89955f
C1461 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v54 GND 0.92879f
C1462 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53 GND 1.14314f
C1463 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v52 GND 0.8323f
C1464 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v51 GND 0.71956f
C1465 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v50 GND 0.79316f
C1466 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39 GND 1.88785f
C1467 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v38 GND 0.87481f
C1468 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37 GND 1.12833f
C1469 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v36 GND 0.79452f
C1470 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v35 GND 0.69232f
C1471 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v34 GND 0.75887f
C1472 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23 GND 1.8686f
C1473 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v22 GND 0.85431f
C1474 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21 GND 1.11076f
C1475 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v20 GND 0.77008f
C1476 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v19 GND 0.66926f
C1477 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v18 GND 0.73878f
C1478 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7 GND 2.26064f
C1479 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v6 GND 0.84054f
C1480 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5 GND 1.1469f
C1481 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v4 GND 0.77243f
C1482 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v3 GND 0.70301f
C1483 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v2 GND 0.72818f
C1484 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_0/sky130_fd_sc_hvl__inv_1_1.A GND 0.9729f
C1485 top_segment_1_0.rseg_1_v3_1.v62 GND 1.00383f
C1486 top_segment_1_0.rseg_1_v3_1.v61 GND 0.94283f
C1487 top_segment_1_0.rseg_1_v3_1.v60 GND 0.92717f
C1488 top_segment_1_0.rseg_1_v3_1.v59 GND 0.86196f
C1489 top_segment_1_0.rseg_1_v3_1.v58 GND 1.47451f
C1490 top_segment_1_0.rseg_1_v3_1.v57 GND 2.4135f
C1491 top_segment_1_0.rseg_1_v3_1.v56 GND 3.29904f
C1492 top_segment_1_0.rseg_1_v3_1.v46 GND 0.999f
C1493 top_segment_1_0.rseg_1_v3_1.v45 GND 0.9622f
C1494 top_segment_1_0.rseg_1_v3_1.v44 GND 0.95203f
C1495 top_segment_1_0.rseg_1_v3_1.v43 GND 0.93445f
C1496 top_segment_1_0.rseg_1_v3_1.v42 GND 1.12363f
C1497 top_segment_1_0.rseg_1_v3_1.v41 GND 2.48462f
C1498 top_segment_1_0.rseg_1_v3_1.v40 GND 3.37108f
C1499 top_segment_1_0.rseg_1_v3_1.v30 GND 1.03387f
C1500 top_segment_1_0.rseg_1_v3_1.v29 GND 0.98141f
C1501 top_segment_1_0.rseg_1_v3_1.v28 GND 0.97038f
C1502 top_segment_1_0.rseg_1_v3_1.v27 GND 0.95434f
C1503 top_segment_1_0.rseg_1_v3_1.v26 GND 1.13854f
C1504 top_segment_1_0.rseg_1_v3_1.v25 GND 2.48866f
C1505 top_segment_1_0.rseg_1_v3_1.v24 GND 3.44747f
C1506 top_segment_1_0.rseg_1_v3_1.v14 GND 1.10941f
C1507 top_segment_1_0.rseg_1_v3_1.v13 GND 1.06449f
C1508 top_segment_1_0.rseg_1_v3_1.v12 GND 1.50227f
C1509 top_segment_1_0.rseg_1_v3_1.v11 GND 1.05333f
C1510 top_segment_1_0.rseg_1_v3_1.v10 GND 1.44211f
C1511 top_segment_1_0.rseg_1_v3_1.v9 GND 2.61871f
C1512 top_segment_1_0.rseg_1_v3_1.v8 GND 4.12386f
C1513 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v61 GND 0.98593f
C1514 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60 GND 1.48196f
C1515 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v59 GND 0.92766f
C1516 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58 GND 2.04138f
C1517 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57 GND 2.40878f
C1518 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56 GND 3.28652f
C1519 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v46 GND 0.83546f
C1520 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v45 GND 0.83142f
C1521 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44 GND 1.31433f
C1522 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v43 GND 0.8334f
C1523 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42 GND 1.49005f
C1524 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41 GND 2.32599f
C1525 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40 GND 3.09657f
C1526 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v30 GND 0.79398f
C1527 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v29 GND 0.79447f
C1528 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28 GND 1.27612f
C1529 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v27 GND 0.80491f
C1530 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26 GND 1.44901f
C1531 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25 GND 2.29709f
C1532 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24 GND 3.04183f
C1533 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v14 GND 0.76536f
C1534 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v13 GND 0.79117f
C1535 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12 GND 1.26691f
C1536 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v11 GND 0.79436f
C1537 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10 GND 1.44302f
C1538 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9 GND 2.29524f
C1539 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8 GND 3.03441f
C1540 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_1/sky130_fd_sc_hvl__inv_1_1.A GND 0.77271f
C1541 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9] GND 4.20597f
C1542 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9] GND 8.05747f
C1543 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8] GND 4.29275f
C1544 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8] GND 3.2508f
C1545 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/sky130_fd_sc_hvl__inv_1_1.A GND 0.76913f
C1546 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/sky130_fd_sc_hvl__inv_1_1.A GND 0.77224f
C1547 top_segment_4_1.bb1 GND 8.29676f
C1548 top_segment_4_1.b1 GND 8.059f
C1549 top_segment_4_1.bb2 GND 8.39631f
C1550 top_segment_4_1.b2 GND 7.53453f
C1551 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.79418f
C1552 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.67704f
C1553 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.643f
C1554 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.61395f
C1555 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.65617f
C1556 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1] GND 10.40641f
C1557 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.67288f
C1558 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.64256f
C1559 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1] GND 9.02532f
C1560 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.61568f
C1561 top_segment_2_0.DEC2[0] GND 18.48324f
C1562 top_segment_4_1.DEC1 GND 6.67564f
C1563 top_segment_2_0.DEC2[1] GND 15.81785f
C1564 top_segment_4_1.DEC2 GND 17.83715f
C1565 top_segment_2_0.DEC2[2] GND 15.65918f
C1566 top_segment_4_1.bb3 GND 13.44233f
C1567 top_segment_4_1.b3 GND 11.34697f
C1568 top_segment_3_0.bb[4] GND 17.38965f
C1569 top_segment_3_0.b[4] GND 17.10753f
C1570 top_segment_3_0.b[5] GND 18.54467f
C1571 top_segment_3_0.bb[5] GND 19.28971f
C1572 top_segment_4_1.DEC3 GND 18.01239f
C1573 top_segment_2_0.DEC2[3] GND 16.77999f
C1574 top_segment_2_0.DEC1[3] GND 15.58448f
C1575 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.Y GND 0.61845f
C1576 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1] GND 7.27954f
C1577 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.Y GND 0.66383f
C1578 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0] GND 7.07277f
C1579 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.Y GND 0.63305f
C1580 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1] GND 7.21126f
C1581 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0] GND 8.73283f
C1582 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.Y GND 0.75299f
C1583 top_segment_2_0.DEC1[2] GND 15.57756f
C1584 top_segment_2_0.DEC1[1] GND 15.53398f
C1585 top_segment_2_0.DEC1[0] GND 15.68788f
C1586 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3] GND 50.81347f
C1587 a_38430_18086# GND 0.21843f $ **FLOATING
C1588 a_35824_18086# GND 0.24267f $ **FLOATING
C1589 a_38430_18467# GND 0.20382f $ **FLOATING
C1590 a_36284_18467# GND 0.18912f $ **FLOATING
C1591 a_38430_18842# GND 0.20634f $ **FLOATING
C1592 a_37164_18842# GND 0.21532f $ **FLOATING
C1593 a_36142_18450# GND 0.15668f $ **FLOATING
C1594 a_35360_18450# GND 0.19962f $ **FLOATING
C1595 a_36142_18748# GND 0.19172f $ **FLOATING
C1596 a_35360_18748# GND 0.19708f $ **FLOATING
C1597 a_38315_19377# GND 0.17117f $ **FLOATING
C1598 a_37131_19377# GND 0.17006f $ **FLOATING
C1599 a_38315_19653# GND 0.17317f $ **FLOATING
C1600 a_37131_19653# GND 0.17331f $ **FLOATING
C1601 a_36351_19283# GND 0.18145f $ **FLOATING
C1602 a_35569_19283# GND 0.17721f $ **FLOATING
C1603 a_36351_19701# GND 0.18276f $ **FLOATING
C1604 a_35569_19701# GND 0.17864f $ **FLOATING
C1605 top_segment_2_0.DEC0[0] GND 17.68075f
C1606 top_segment_2_0.DEC0[1] GND 17.46284f
C1607 top_segment_2_0.DEC0[2] GND 18.90041f
C1608 top_segment_3_0.bb[6] GND 17.33524f
C1609 top_segment_3_0.b[6] GND 17.90471f
C1610 a_39072_20445# GND 0.05335f $ **FLOATING
C1611 a_38408_20445# GND 0.01074f $ **FLOATING
C1612 a_40454_21045# GND 0.01121f $ **FLOATING
C1613 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV GND 11.21902f
C1614 a_42614_21484# GND 0.18164f $ **FLOATING
C1615 a_38408_21484# GND 0.0387f $ **FLOATING
C1616 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV GND 19.55606f
C1617 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC GND 4.69893f
C1618 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC GND 11.75439f
C1619 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3 GND 0.2652f
C1620 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1 GND 0.28781f
C1621 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2 GND 2.93597f
C1622 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4 GND 3.21084f
C1623 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0 GND 2.10079f
C1624 top_segment_2_0.V0 GND 9.79343f
C1625 ROUT.t3 GND 0.02488f
C1626 ROUT.t0 GND 1.41742f
C1627 ROUT.t4 GND 2.04267f
C1628 ROUT.t5 GND 2.33027f
C1629 ROUT.t2 GND 1.70501f
C1630 ROUT.n0 GND 1.47089f
C1631 ROUT.n1 GND 0.21478f
C1632 ROUT.t1 GND 0.02473f
C1633 ROUT.n2 GND 0.02835f
C1634 ROUT.n3 GND 0.09357f
C1635 top_segment_1_0.rseg_1_v3_1.v41.t2 GND 0.04657f
C1636 top_segment_1_0.rseg_1_v3_1.v41.t1 GND 0.13984f
C1637 top_segment_1_0.rseg_1_v3_1.v41.t0 GND 0.13973f
C1638 top_segment_1_0.rseg_1_v3_1.v41.n0 GND 2.57846f
C1639 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t2 GND 0.02245f
C1640 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t1 GND 0.13085f
C1641 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.t0 GND 0.40072f
C1642 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v40.n0 GND 2.7728f
C1643 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t2 GND 0.0125f
C1644 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t1 GND 0.08878f
C1645 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.t0 GND 0.0907f
C1646 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v39.n0 GND 1.58019f
C1647 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t1 GND 0.01506f
C1648 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t2 GND 0.09069f
C1649 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.t0 GND 0.08797f
C1650 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v44.n0 GND 1.45497f
C1651 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t1 GND 0.02728f
C1652 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t2 GND 0.1501f
C1653 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.t0 GND 0.16768f
C1654 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v41.n0 GND 2.84284f
C1655 a_13219_17684.t2 GND 0.03023f
C1656 a_13219_17684.t1 GND 0.02819f
C1657 a_13219_17684.n0 GND 0.98182f
C1658 a_13219_17684.t3 GND 0.02853f
C1659 a_13219_17684.n1 GND 1.49664f
C1660 a_13219_17684.t0 GND 0.0346f
C1661 a_22130_19162.t1 GND 0.13926f
C1662 a_22130_19162.t2 GND 0.0925f
C1663 a_22130_19162.n0 GND 5.29359f
C1664 a_22130_19162.t3 GND 0.17307f
C1665 a_22130_19162.n1 GND 5.33077f
C1666 a_22130_19162.t0 GND 0.07081f
C1667 a_27705_5238.t4 GND 0.14531f
C1668 a_27705_5238.t1 GND 0.08367f
C1669 a_27705_5238.n0 GND 4.77562f
C1670 a_27705_5238.t2 GND 0.14572f
C1671 a_27705_5238.n1 GND 4.0453f
C1672 a_27705_5238.t3 GND 0.17762f
C1673 a_27705_5238.n2 GND 6.44309f
C1674 a_27705_5238.t0 GND 0.08367f
C1675 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t1 GND 0.02752f
C1676 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t2 GND 0.15141f
C1677 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.t0 GND 0.17047f
C1678 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v9.n0 GND 2.83038f
C1679 top_segment_2_0.rseg_2_v3_0.v28.t2 GND 0.10104f
C1680 top_segment_2_0.rseg_2_v3_0.v28.t1 GND 0.09807f
C1681 top_segment_2_0.rseg_2_v3_0.v28.n0 GND 1.8875f
C1682 top_segment_2_0.rseg_2_v3_0.v28.t0 GND 0.01339f
C1683 a_14176_6674.t3 GND 0.0947f
C1684 a_14176_6674.t2 GND 0.07612f
C1685 a_14176_6674.n0 GND 5.33217f
C1686 a_14176_6674.t1 GND 0.07612f
C1687 a_14176_6674.n1 GND 2.97065f
C1688 a_14176_6674.t4 GND 0.08576f
C1689 a_14176_6674.n2 GND 3.98477f
C1690 a_14176_6674.t0 GND 0.07971f
C1691 a_21302_19162.t2 GND 0.16937f
C1692 a_21302_19162.t3 GND 0.15559f
C1693 a_21302_19162.t4 GND 0.06731f
C1694 a_21302_19162.n0 GND 4.60037f
C1695 a_21302_19162.t1 GND 0.06731f
C1696 a_21302_19162.n1 GND 0.88718f
C1697 a_21302_19162.n2 GND 4.88352f
C1698 a_21302_19162.t0 GND 0.06934f
C1699 a_22756_17121.t2 GND 0.04042f
C1700 a_22756_17121.t1 GND 0.03955f
C1701 a_22756_17121.t3 GND 0.03423f
C1702 a_22756_17121.n0 GND 1.24539f
C1703 a_22756_17121.t4 GND 0.03423f
C1704 a_22756_17121.n1 GND 0.78371f
C1705 a_22756_17121.n2 GND 1.28824f
C1706 a_22756_17121.t0 GND 0.03423f
C1707 SH[3].t1 GND 0.12078f
C1708 SH[3].n0 GND 0.04952f
C1709 SH[3].n1 GND 0.10661f
C1710 SH[3].n2 GND 0.07078f
C1711 SH[3].t0 GND 0.11571f
C1712 SH[3].n3 GND 0.01462f
C1713 SH[3].n4 GND 0.08197f
C1714 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t2 GND 0.01662f
C1715 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t1 GND 0.09404f
C1716 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.t0 GND 0.09697f
C1717 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v60.n0 GND 1.57947f
C1718 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t1 GND 0.01438f
C1719 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t2 GND 0.08736f
C1720 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.t0 GND 0.07781f
C1721 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v10.n0 GND 1.43709f
C1722 top_segment_2_0.rseg_2_v3_0.v27.t2 GND 0.10482f
C1723 top_segment_2_0.rseg_2_v3_0.v27.t1 GND 0.10131f
C1724 top_segment_2_0.rseg_2_v3_0.v27.n0 GND 1.97943f
C1725 top_segment_2_0.rseg_2_v3_0.v27.t0 GND 0.01445f
C1726 top_segment_2_0.rseg_2_v3_0.v37.t1 GND 0.11065f
C1727 top_segment_2_0.rseg_2_v3_0.v37.t2 GND 0.0154f
C1728 top_segment_2_0.rseg_2_v3_0.v37.n0 GND 2.06691f
C1729 top_segment_2_0.rseg_2_v3_0.v37.t0 GND 0.10705f
C1730 a_30417_6674.t4 GND 0.05828f
C1731 a_30417_6674.t1 GND 0.04276f
C1732 a_30417_6674.n0 GND 2.03892f
C1733 a_30417_6674.t2 GND 0.04087f
C1734 a_30417_6674.n1 GND 1.29976f
C1735 a_30417_6674.t3 GND 0.07543f
C1736 a_30417_6674.n2 GND 3.00311f
C1737 a_30417_6674.t0 GND 0.04087f
C1738 SH[1].t1 GND 0.0605f
C1739 SH[1].n0 GND 0.02481f
C1740 SH[1].n1 GND 0.0534f
C1741 SH[1].n2 GND 0.03545f
C1742 SH[1].t0 GND 0.05796f
C1743 SH[1].n4 GND 0.04106f
C1744 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t1 GND 0.09569f
C1745 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_2.Y GND 0.31167f
C1746 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n0 GND 0.02473f
C1747 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t2 GND 0.30126f
C1748 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[4] GND 5.44042f
C1749 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[4] GND 0.68417f
C1750 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.n1 GND 0.21176f
C1751 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.INB.t0 GND 0.13031f
C1752 a_12326_5238.t1 GND 0.04948f
C1753 a_12326_5238.t2 GND 0.039f
C1754 a_12326_5238.n0 GND 2.59143f
C1755 a_12326_5238.t4 GND 0.04849f
C1756 a_12326_5238.t3 GND 0.039f
C1757 a_12326_5238.n1 GND 2.19006f
C1758 a_12326_5238.n2 GND 2.38608f
C1759 a_12326_5238.t0 GND 0.05645f
C1760 top_segment_1_0.rseg_1_v3_1.v12.t2 GND 0.02587f
C1761 top_segment_1_0.rseg_1_v3_1.v12.t1 GND 0.07997f
C1762 top_segment_1_0.rseg_1_v3_1.v12.t0 GND 0.07985f
C1763 top_segment_1_0.rseg_1_v3_1.v12.n0 GND 1.3573f
C1764 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t1 GND 0.02716f
C1765 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t2 GND 0.1492f
C1766 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.t0 GND 0.16449f
C1767 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v57.n0 GND 2.95161f
C1768 a_33127_7938.t1 GND 0.10677f
C1769 a_33127_7938.t2 GND 0.12828f
C1770 a_33127_7938.n0 GND 6.09613f
C1771 a_33127_7938.t0 GND 0.06882f
C1772 a_21578_19162.t2 GND 0.15567f
C1773 a_21578_19162.t1 GND 0.07037f
C1774 a_21578_19162.n0 GND 4.70467f
C1775 a_21578_19162.t3 GND 0.16064f
C1776 a_21578_19162.n1 GND 4.64301f
C1777 a_21578_19162.t0 GND 0.06564f
C1778 a_32457_7938.t2 GND 0.10902f
C1779 a_32457_7938.t1 GND 0.0723f
C1780 a_32457_7938.n0 GND 5.42682f
C1781 a_32457_7938.t0 GND 0.09187f
C1782 top_segment_2_0.rseg_2_v3_0.v3.t1 GND 0.03836f
C1783 top_segment_2_0.rseg_2_v3_0.v3.t2 GND 0.19594f
C1784 top_segment_2_0.rseg_2_v3_0.v3.n0 GND 4.27168f
C1785 top_segment_2_0.rseg_2_v3_0.v3.t0 GND 0.19402f
C1786 top_segment_2_0.rseg_2_v3_0.v38.t1 GND 0.19941f
C1787 top_segment_2_0.rseg_2_v3_0.v38.t2 GND 0.02987f
C1788 top_segment_2_0.rseg_2_v3_0.v38.n0 GND 4.06638f
C1789 top_segment_2_0.rseg_2_v3_0.v38.t0 GND 0.20435f
C1790 top_segment_1_0.rseg_1_v3_1.v40.t2 GND 0.03678f
C1791 top_segment_1_0.rseg_1_v3_1.v40.t1 GND 0.12307f
C1792 top_segment_1_0.rseg_1_v3_1.v40.t0 GND 0.36728f
C1793 top_segment_1_0.rseg_1_v3_1.v40.n0 GND 2.56971f
C1794 a_17547_7938.t2 GND 0.07342f
C1795 a_17547_7938.t1 GND 0.07455f
C1796 a_17547_7938.n0 GND 5.18539f
C1797 a_17547_7938.t0 GND 0.06664f
C1798 a_20750_19162.t1 GND 0.17024f
C1799 a_20750_19162.t2 GND 0.14851f
C1800 a_20750_19162.t3 GND 0.05862f
C1801 a_20750_19162.n0 GND 4.26715f
C1802 a_20750_19162.n1 GND 5.08543f
C1803 a_20750_19162.t0 GND 0.07006f
C1804 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t1 GND 0.01583f
C1805 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t2 GND 0.09012f
C1806 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.t0 GND 0.08109f
C1807 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v58.n0 GND 1.56677f
C1808 a_19370_19162.t1 GND 0.15734f
C1809 a_19370_19162.t4 GND 0.05584f
C1810 a_19370_19162.n0 GND 4.21706f
C1811 a_19370_19162.t2 GND 0.05584f
C1812 a_19370_19162.n1 GND 0.59217f
C1813 a_19370_19162.t3 GND 0.16998f
C1814 a_19370_19162.n2 GND 4.88166f
C1815 a_19370_19162.t0 GND 0.07011f
C1816 a_14728_6674.t3 GND 0.09319f
C1817 a_14728_6674.t2 GND 0.07394f
C1818 a_14728_6674.n0 GND 5.40641f
C1819 a_14728_6674.t1 GND 0.07394f
C1820 a_14728_6674.n1 GND 2.82116f
C1821 a_14728_6674.t4 GND 0.07704f
C1822 a_14728_6674.n2 GND 3.67426f
C1823 a_14728_6674.t0 GND 0.08006f
C1824 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t2 GND 0.02279f
C1825 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t0 GND 0.13331f
C1826 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.t1 GND 0.39585f
C1827 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v8.n0 GND 2.76318f
C1828 a_12602_5238.t1 GND 0.09741f
C1829 a_12602_5238.t2 GND 0.07626f
C1830 a_12602_5238.n0 GND 5.27749f
C1831 a_12602_5238.t4 GND 0.09544f
C1832 a_12602_5238.t3 GND 0.07626f
C1833 a_12602_5238.n1 GND 4.32003f
C1834 a_12602_5238.n2 GND 4.74566f
C1835 a_12602_5238.t0 GND 0.11145f
C1836 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t0 GND 0.01441f
C1837 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t2 GND 0.07654f
C1838 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.t1 GND 0.08569f
C1839 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v42.n0 GND 1.43498f
C1840 top_segment_2_0.DEC1[2].t6 GND 0.17266f
C1841 top_segment_2_0.DEC1[2].t4 GND 0.17211f
C1842 top_segment_2_0.DEC1[2].n0 GND 0.24239f
C1843 top_segment_2_0.DEC1[2].t9 GND 0.17306f
C1844 top_segment_2_0.DEC1[2].t2 GND 0.17211f
C1845 top_segment_2_0.DEC1[2].n1 GND 0.60536f
C1846 top_segment_2_0.DEC1[2].n2 GND 0.18843f
C1847 top_segment_2_0.DEC1[2].t7 GND 0.16963f
C1848 top_segment_2_0.DEC1[2].n3 GND 16.2245f
C1849 top_segment_2_0.DEC1[2].t5 GND 0.5519f
C1850 top_segment_2_0.DEC1[2].t1 GND 0.12067f
C1851 top_segment_2_0.DEC1[2].t0 GND 0.14179f
C1852 top_segment_2_0.DEC1[2].n4 GND 0.78071f
C1853 top_segment_2_0.DEC1[2].n5 GND 0.62147f
C1854 top_segment_2_0.DEC1[2].t8 GND 0.56361f
C1855 top_segment_2_0.DEC1[2].t3 GND 0.56124f
C1856 top_segment_2_0.DEC1[2].n6 GND 1.24769f
C1857 top_segment_2_0.DEC1[2].n7 GND 0.92779f
C1858 top_segment_3_0.rseg_3_v3_0.v8.t2 GND 0.16796f
C1859 top_segment_3_0.rseg_3_v3_0.v8.t1 GND 0.63095f
C1860 top_segment_3_0.rseg_3_v3_0.v8.n0 GND 4.13463f
C1861 top_segment_3_0.rseg_3_v3_0.v8.t3 GND 0.02217f
C1862 top_segment_3_0.rseg_3_v3_0.v8.n1 GND 1.41681f
C1863 top_segment_3_0.rseg_3_v3_0.v8.t0 GND 0.02748f
C1864 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.Y GND 0.58917f
C1865 top_segment_4_1.b0.t1 GND 0.1033f
C1866 top_segment_4_1.b0.n0 GND 0.04235f
C1867 top_segment_4_1.b0.n1 GND 0.09117f
C1868 top_segment_4_1.b0.n2 GND 0.06053f
C1869 top_segment_4_1.b0.t3 GND 1.65873f
C1870 top_segment_1_0.b[0] GND 0.20711f
C1871 top_segment_4_1.b0.t2 GND 0.19215f
C1872 top_segment_4_1.b0.n3 GND 2.02603f
C1873 top_segment_4_1.b0.n4 GND 22.6437f
C1874 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.b[0] GND 3.71602f
C1875 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUT GND 0.35439f
C1876 top_segment_4_1.b0.n5 GND 0.06516f
C1877 top_segment_4_1.b0.t0 GND 0.09896f
C1878 top_segment_4_1.b0.n6 GND 0.05119f
C1879 top_segment_3_0.rseg_3_v3_0.v7.t2 GND 0.08527f
C1880 top_segment_3_0.rseg_3_v3_0.v7.t1 GND 0.08305f
C1881 top_segment_3_0.rseg_3_v3_0.v7.n0 GND 1.91518f
C1882 top_segment_3_0.rseg_3_v3_0.v7.t0 GND 0.01651f
C1883 top_segment_3_0.rseg_3_v3_0.v6.t1 GND 0.11479f
C1884 top_segment_3_0.rseg_3_v3_0.v6.t2 GND 0.11222f
C1885 top_segment_3_0.rseg_3_v3_0.v6.n0 GND 2.55165f
C1886 top_segment_3_0.rseg_3_v3_0.v6.t0 GND 0.02134f
C1887 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t2 GND 0.01294f
C1888 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t1 GND 0.10145f
C1889 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.t0 GND 0.09797f
C1890 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v5.n0 GND 1.62712f
C1891 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t3 GND 0.1968f
C1892 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t0 GND 0.20388f
C1893 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t1 GND 0.19134f
C1894 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n0 GND 1.5154f
C1895 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.n1 GND 0.75134f
C1896 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S2.t2 GND 0.39307f
C1897 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t2 GND 0.02762f
C1898 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t3 GND 0.02762f
C1899 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n0 GND 0.06586f
C1900 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.Y GND 0.21353f
C1901 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n1 GND 0.12938f
C1902 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t4 GND 0.72401f
C1903 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n2 GND 15.9934f
C1904 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n3 GND 0.04026f
C1905 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t1 GND 0.04249f
C1906 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.t0 GND 0.04249f
C1907 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.IN.n4 GND 0.09332f
C1908 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t1 GND 0.04053f
C1909 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t2 GND 0.04053f
C1910 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n0 GND 0.089f
C1911 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x1.Y GND 0.20365f
C1912 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n1 GND 0.03839f
C1913 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t7 GND 0.06304f
C1914 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t4 GND 0.03715f
C1915 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t6 GND 0.06304f
C1916 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t8 GND 0.03715f
C1917 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n2 GND 0.10577f
C1918 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n3 GND 0.15692f
C1919 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_4.x2.A GND 0.01051f
C1920 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n4 GND 0.04732f
C1921 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t5 GND 0.51546f
C1922 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n5 GND 15.6837f
C1923 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n6 GND 0.02899f
C1924 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t3 GND 0.02634f
C1925 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.t0 GND 0.02634f
C1926 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n7 GND 0.06281f
C1927 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_3/lvsf_0.INB.n8 GND 0.1234f
C1928 a_30141_6674.t4 GND 0.11133f
C1929 a_30141_6674.t1 GND 0.08541f
C1930 a_30141_6674.n0 GND 3.94271f
C1931 a_30141_6674.t2 GND 0.08147f
C1932 a_30141_6674.n1 GND 2.66272f
C1933 a_30141_6674.t3 GND 0.14987f
C1934 a_30141_6674.n2 GND 5.98504f
C1935 a_30141_6674.t0 GND 0.08147f
C1936 a_20198_19162.t1 GND 0.21223f
C1937 a_20198_19162.t3 GND 0.15786f
C1938 a_20198_19162.t2 GND 0.0607f
C1939 a_20198_19162.n0 GND 4.57762f
C1940 a_20198_19162.n1 GND 6.60332f
C1941 a_20198_19162.t0 GND 0.08827f
C1942 a_22958_19162.t1 GND 0.17057f
C1943 a_22958_19162.t3 GND 0.16728f
C1944 a_22958_19162.t2 GND 0.0867f
C1945 a_22958_19162.n0 GND 5.40937f
C1946 a_22958_19162.n1 GND 4.89637f
C1947 a_22958_19162.t0 GND 0.06972f
C1948 a_21016_17121.t3 GND 0.07551f
C1949 a_21016_17121.t2 GND 0.06407f
C1950 a_21016_17121.t1 GND 0.06237f
C1951 a_21016_17121.n0 GND 1.93846f
C1952 a_21016_17121.t4 GND 0.0628f
C1953 a_21016_17121.n1 GND 1.70138f
C1954 a_21016_17121.t5 GND 0.0628f
C1955 a_21016_17121.n2 GND 1.51601f
C1956 a_21016_17121.n3 GND 2.55379f
C1957 a_21016_17121.t0 GND 0.0628f
C1958 a_13771_17684.t1 GND 0.02918f
C1959 a_13771_17684.t2 GND 0.03032f
C1960 a_13771_17684.n0 GND 2.00335f
C1961 a_13771_17684.t0 GND 0.03715f
C1962 top_segment_2_0.rseg_2_v3_0.v21.t2 GND 0.10089f
C1963 top_segment_2_0.rseg_2_v3_0.v21.t1 GND 0.01431f
C1964 top_segment_2_0.rseg_2_v3_0.v21.n0 GND 1.89096f
C1965 top_segment_2_0.rseg_2_v3_0.v21.t0 GND 0.09384f
C1966 a_23234_19162.t1 GND 0.16517f
C1967 a_23234_19162.t3 GND 0.12791f
C1968 a_23234_19162.t2 GND 0.07601f
C1969 a_23234_19162.n0 GND 4.60987f
C1970 a_23234_19162.n1 GND 5.15358f
C1971 a_23234_19162.t0 GND 0.06747f
C1972 a_32733_7938.t2 GND 0.11818f
C1973 a_32733_7938.t1 GND 0.07481f
C1974 a_32733_7938.n0 GND 5.80655f
C1975 a_32733_7938.t0 GND 0.10046f
C1976 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t1 GND -0.50828f
C1977 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t0 GND -3.67942f
C1978 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t4 GND -2.37382f
C1979 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t3 GND -2.36382f
C1980 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n0 GND -3.97308f
C1981 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].t2 GND -2.36382f
C1982 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n1 GND -3.49244f
C1983 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec0[3].n2 GND -5.38322f
C1984 top_segment_3_0.rseg_3_v3_0.v11.t1 GND 0.07822f
C1985 top_segment_3_0.rseg_3_v3_0.v11.t2 GND 0.01384f
C1986 top_segment_3_0.rseg_3_v3_0.v11.n0 GND 1.81943f
C1987 top_segment_3_0.rseg_3_v3_0.v11.t0 GND 0.08852f
C1988 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t1 GND 0.01248f
C1989 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t2 GND 0.08856f
C1990 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.t0 GND 0.09062f
C1991 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v7.n0 GND 1.58095f
C1992 top_segment_1_0.rseg_1_v3_1.v57.t1 GND 0.04652f
C1993 top_segment_1_0.rseg_1_v3_1.v57.t0 GND 0.13968f
C1994 top_segment_1_0.rseg_1_v3_1.v57.t2 GND 0.13957f
C1995 top_segment_1_0.rseg_1_v3_1.v57.n0 GND 2.57959f
C1996 a_12878_5238.t1 GND 0.0968f
C1997 a_12878_5238.t2 GND 0.07529f
C1998 a_12878_5238.n0 GND 5.41272f
C1999 a_12878_5238.t4 GND 0.09483f
C2000 a_12878_5238.t3 GND 0.07529f
C2001 a_12878_5238.n1 GND 4.30036f
C2002 a_12878_5238.n2 GND 4.73412f
C2003 a_12878_5238.t0 GND 0.1106f
C2004 a_25891_5238.t4 GND 0.06897f
C2005 a_25891_5238.t1 GND 0.04091f
C2006 a_25891_5238.n0 GND 2.62657f
C2007 a_25891_5238.t2 GND 0.08929f
C2008 a_25891_5238.n1 GND 2.43648f
C2009 a_25891_5238.t3 GND 0.08534f
C2010 a_25891_5238.n2 GND 2.71152f
C2011 a_25891_5238.t0 GND 0.04091f
C2012 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t3 GND 0.02769f
C2013 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t2 GND 0.02769f
C2014 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n0 GND 0.06602f
C2015 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x1.Y GND 0.21405f
C2016 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n1 GND 0.1297f
C2017 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t5 GND 0.06626f
C2018 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t8 GND 0.03905f
C2019 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t4 GND 0.06626f
C2020 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t7 GND 0.03905f
C2021 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n2 GND 0.11117f
C2022 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n3 GND 0.16493f
C2023 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.A GND 0.01104f
C2024 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n4 GND 0.04974f
C2025 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t6 GND 0.51398f
C2026 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n5 GND 16.3238f
C2027 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n6 GND 0.03047f
C2028 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n7 GND 0.04035f
C2029 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t0 GND 0.04259f
C2030 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.t1 GND 0.04259f
C2031 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.INB.n8 GND 0.09355f
C2032 top_segment_2_0.rseg_2_v3_0.v24.t2 GND 0.16286f
C2033 top_segment_2_0.rseg_2_v3_0.v24.t1 GND 0.59039f
C2034 top_segment_2_0.rseg_2_v3_0.v24.n0 GND 4.42116f
C2035 top_segment_2_0.rseg_2_v3_0.v24.t0 GND 0.0256f
C2036 a_15990_6674.t3 GND 0.04624f
C2037 a_15990_6674.t2 GND 0.03583f
C2038 a_15990_6674.n0 GND 2.81877f
C2039 a_15990_6674.t1 GND 0.03583f
C2040 a_15990_6674.n1 GND 1.26954f
C2041 a_15990_6674.t4 GND 0.0365f
C2042 a_15990_6674.n2 GND 2.11432f
C2043 a_15990_6674.t0 GND 0.04297f
C2044 SH[4].t1 GND 0.11131f
C2045 SH[4].n0 GND 0.04564f
C2046 SH[4].n1 GND 0.09824f
C2047 SH[4].n2 GND 0.06522f
C2048 SH[4].t0 GND 0.10663f
C2049 SH[4].n3 GND 0.01347f
C2050 SH[4].n4 GND 0.07554f
C2051 a_22682_19162.t1 GND 0.15093f
C2052 a_22682_19162.t2 GND 0.0995f
C2053 a_22682_19162.n0 GND 5.6647f
C2054 a_22682_19162.t3 GND 0.17697f
C2055 a_22682_19162.n1 GND 5.33538f
C2056 a_22682_19162.t0 GND 0.07252f
C2057 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t2 GND 0.01499f
C2058 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t1 GND 0.08877f
C2059 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.t0 GND 0.09145f
C2060 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v12.n0 GND 1.46182f
C2061 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t3 GND 0.0247f
C2062 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t2 GND 0.0247f
C2063 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n0 GND 0.05889f
C2064 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.Y GND 0.19095f
C2065 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n1 GND 0.1157f
C2066 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t4 GND 0.70975f
C2067 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n2 GND 14.2799f
C2068 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n3 GND 0.036f
C2069 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t1 GND 0.038f
C2070 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.t0 GND 0.038f
C2071 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.IN.n4 GND 0.08345f
C2072 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t1 GND 0.01209f
C2073 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t2 GND 0.08547f
C2074 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.t0 GND 0.08753f
C2075 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v55.n0 GND 1.50136f
C2076 top_segment_2_0.rseg_2_v3_0.v11.t2 GND 0.01522f
C2077 top_segment_2_0.rseg_2_v3_0.v11.t1 GND 0.09422f
C2078 top_segment_2_0.rseg_2_v3_0.v11.n0 GND 1.89603f
C2079 top_segment_2_0.rseg_2_v3_0.v11.t0 GND 0.09453f
C2080 top_segment_1_0.rseg_1_v3_1.v24.t0 GND 0.03636f
C2081 top_segment_1_0.rseg_1_v3_1.v24.t1 GND 0.12209f
C2082 top_segment_1_0.rseg_1_v3_1.v24.t2 GND 0.36895f
C2083 top_segment_1_0.rseg_1_v3_1.v24.n0 GND 2.57743f
C2084 a_27981_5238.t4 GND 0.07592f
C2085 a_27981_5238.t1 GND 0.04358f
C2086 a_27981_5238.n0 GND 2.54446f
C2087 a_27981_5238.t2 GND 0.06837f
C2088 a_27981_5238.n1 GND 1.92423f
C2089 a_27981_5238.t3 GND 0.09262f
C2090 a_27981_5238.n2 GND 3.30724f
C2091 a_27981_5238.t0 GND 0.04358f
C2092 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_0.Y GND 0.52659f
C2093 top_segment_4_1.bb0.t1 GND 0.09973f
C2094 top_segment_4_1.bb0.n0 GND 0.04089f
C2095 top_segment_4_1.bb0.n1 GND 0.08803f
C2096 top_segment_4_1.bb0.n2 GND 0.05844f
C2097 top_segment_4_1.bb0.t2 GND 1.63719f
C2098 top_segment_1_0.bb[0] GND 0.20459f
C2099 top_segment_4_1.bb0.t5 GND 0.18552f
C2100 top_segment_4_1.bb0.n3 GND 1.90581f
C2101 top_segment_4_1.bb0.n4 GND 21.8065f
C2102 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.bb[0] GND 3.50091f
C2103 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.OUTB GND 0.35162f
C2104 top_segment_4_1.bb0.t3 GND 0.3488f
C2105 top_segment_4_1.bb0.t4 GND 0.19349f
C2106 top_segment_4_1.bb0.n5 GND 0.30394f
C2107 top_segment_4_1.bb0.n6 GND 0.06047f
C2108 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/buff_hvl_0.sky130_fd_sc_hvl__inv_1_1.A GND 0.15587f
C2109 top_segment_4_1.bb0.n7 GND 0.0867f
C2110 top_segment_4_1.bb0.n8 GND 0.04942f
C2111 top_segment_4_1.bb0.t0 GND 0.09555f
C2112 a_27153_5238.t4 GND 0.12539f
C2113 a_27153_5238.t1 GND 0.07275f
C2114 a_27153_5238.n0 GND 3.93804f
C2115 a_27153_5238.t2 GND 0.15297f
C2116 a_27153_5238.n1 GND 4.11942f
C2117 a_27153_5238.t3 GND 0.15386f
C2118 a_27153_5238.n2 GND 5.76483f
C2119 a_27153_5238.t0 GND 0.07275f
C2120 a_21854_19162.t1 GND 0.12979f
C2121 a_21854_19162.t3 GND 0.07321f
C2122 a_21854_19162.n0 GND 4.33997f
C2123 a_21854_19162.t2 GND 0.07321f
C2124 a_21854_19162.n1 GND 1.20642f
C2125 a_21854_19162.t4 GND 0.1514f
C2126 a_21854_19162.n2 GND 4.46413f
C2127 a_21854_19162.t0 GND 0.06185f
C2128 a_20740_17121.t2 GND 0.04172f
C2129 a_20740_17121.t1 GND 0.04844f
C2130 a_20740_17121.t3 GND 0.03452f
C2131 a_20740_17121.n0 GND 1.72763f
C2132 a_20740_17121.t4 GND 0.03452f
C2133 a_20740_17121.n1 GND 0.84517f
C2134 a_20740_17121.n2 GND 1.43346f
C2135 a_20740_17121.t0 GND 0.03452f
C2136 a_13864_5238.t1 GND 0.09555f
C2137 a_13864_5238.t2 GND 0.07299f
C2138 a_13864_5238.n0 GND 4.6643f
C2139 a_13864_5238.t4 GND 0.09358f
C2140 a_13864_5238.t3 GND 0.07299f
C2141 a_13864_5238.n1 GND 5.4004f
C2142 a_13864_5238.n2 GND 4.00369f
C2143 a_13864_5238.t0 GND 0.0965f
C2144 SH[2].t1 GND 0.12244f
C2145 SH[2].n0 GND 0.0502f
C2146 SH[2].n1 GND 0.10807f
C2147 SH[2].n2 GND 0.07175f
C2148 SH[2].t0 GND 0.1173f
C2149 SH[2].n3 GND 0.01482f
C2150 SH[2].n4 GND 0.08309f
C2151 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t3 GND 0.0261f
C2152 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t2 GND 0.0261f
C2153 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n0 GND 0.06224f
C2154 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x1.Y GND 0.20181f
C2155 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n1 GND 0.12228f
C2156 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t5 GND 0.06247f
C2157 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t8 GND 0.03681f
C2158 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t4 GND 0.06247f
C2159 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t6 GND 0.03681f
C2160 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n2 GND 0.10482f
C2161 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n3 GND 0.1555f
C2162 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_11.x2.A GND 0.01041f
C2163 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n4 GND 0.04689f
C2164 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t7 GND 0.57365f
C2165 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n5 GND 15.4363f
C2166 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n6 GND 0.02873f
C2167 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n7 GND 0.03805f
C2168 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t1 GND 0.04016f
C2169 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.t0 GND 0.04016f
C2170 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_0/lvsf_0.INB.n8 GND 0.0882f
C2171 a_13495_17684.t1 GND 0.06282f
C2172 a_13495_17684.t2 GND 0.0622f
C2173 a_13495_17684.n0 GND 4.49915f
C2174 a_13495_17684.t0 GND 0.07583f
C2175 top_segment_2_0.DEC1[1].t6 GND 0.17284f
C2176 top_segment_2_0.DEC1[1].t4 GND 0.17234f
C2177 top_segment_2_0.DEC1[1].n0 GND 0.21906f
C2178 top_segment_2_0.DEC1[1].t3 GND 0.17321f
C2179 top_segment_2_0.DEC1[1].t5 GND 0.17234f
C2180 top_segment_2_0.DEC1[1].n1 GND 0.56133f
C2181 top_segment_2_0.DEC1[1].n2 GND 0.18922f
C2182 top_segment_2_0.DEC1[1].t9 GND 0.17035f
C2183 top_segment_2_0.DEC1[1].n3 GND 16.4341f
C2184 top_segment_2_0.DEC1[1].t0 GND 0.1425f
C2185 top_segment_2_0.DEC1[1].t1 GND 0.12117f
C2186 top_segment_2_0.DEC1[1].n4 GND 0.97482f
C2187 top_segment_2_0.DEC1[1].t2 GND 0.56576f
C2188 top_segment_2_0.DEC1[1].t7 GND 0.56342f
C2189 top_segment_2_0.DEC1[1].n5 GND 0.89432f
C2190 top_segment_2_0.DEC1[1].n6 GND 0.57694f
C2191 top_segment_2_0.DEC1[1].t8 GND 0.595f
C2192 top_segment_2_0.DEC1[1].n7 GND 1.24415f
C2193 a_14140_5238.t1 GND 0.09595f
C2194 a_14140_5238.t2 GND 0.07288f
C2195 a_14140_5238.n0 GND 4.84371f
C2196 a_14140_5238.t4 GND 0.09395f
C2197 a_14140_5238.t3 GND 0.07288f
C2198 a_14140_5238.n1 GND 5.40773f
C2199 a_14140_5238.n2 GND 3.72117f
C2200 a_14140_5238.t0 GND 0.09172f
C2201 a_20474_19162.t1 GND 0.18645f
C2202 a_20474_19162.t3 GND 0.14562f
C2203 a_20474_19162.t2 GND 0.05846f
C2204 a_20474_19162.n0 GND 4.28874f
C2205 a_20474_19162.n1 GND 5.74363f
C2206 a_20474_19162.t0 GND 0.0771f
C2207 a_29865_6674.t4 GND 0.10563f
C2208 a_29865_6674.t1 GND 0.08474f
C2209 a_29865_6674.n0 GND 3.77304f
C2210 a_29865_6674.t2 GND 0.08064f
C2211 a_29865_6674.n1 GND 2.70857f
C2212 a_29865_6674.t3 GND 0.14779f
C2213 a_29865_6674.n2 GND 5.91896f
C2214 a_29865_6674.t0 GND 0.08064f
C2215 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t3 GND 0.0257f
C2216 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t2 GND 0.0257f
C2217 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n0 GND 0.06128f
C2218 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x2.Y GND 0.19868f
C2219 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n1 GND 0.12038f
C2220 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t4 GND 0.06536f
C2221 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t5 GND 0.04079f
C2222 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n2 GND 0.12995f
C2223 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.B GND 0.05637f
C2224 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.A GND 0.02254f
C2225 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t7 GND 0.06545f
C2226 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t8 GND 0.04086f
C2227 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n3 GND 0.12458f
C2228 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n4 GND 0.02451f
C2229 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n5 GND 0.06185f
C2230 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[1] GND 2.34134f
C2231 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t6 GND 0.24665f
C2232 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n6 GND 11.5282f
C2233 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n7 GND 2.61648f
C2234 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n8 GND 0.03746f
C2235 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t1 GND 0.03954f
C2236 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.t0 GND 0.03954f
C2237 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.IN.n9 GND 0.08683f
C2238 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t1 GND 0.02477f
C2239 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t2 GND 0.02477f
C2240 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n0 GND 0.05907f
C2241 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_6.x1.Y GND 0.19154f
C2242 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n1 GND 0.11606f
C2243 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t12 GND 0.05929f
C2244 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t7 GND 0.03494f
C2245 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t11 GND 0.05929f
C2246 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t4 GND 0.03494f
C2247 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n2 GND 0.09948f
C2248 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n3 GND 0.14758f
C2249 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n4 GND 0.04451f
C2250 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t9 GND 0.06301f
C2251 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t10 GND 0.03932f
C2252 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n5 GND 0.12528f
C2253 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.A GND 0.02173f
C2254 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t5 GND 0.06309f
C2255 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t8 GND 0.03939f
C2256 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n6 GND 0.1201f
C2257 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n7 GND 0.03507f
C2258 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.B GND 0.1019f
C2259 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[1] GND 2.24751f
C2260 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t6 GND 0.23705f
C2261 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n8 GND 9.91961f
C2262 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n9 GND 3.7575f
C2263 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n10 GND 0.02727f
C2264 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n11 GND 0.03611f
C2265 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t3 GND 0.03811f
C2266 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.t0 GND 0.03811f
C2267 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_4/lvsf_0.INB.n12 GND 0.08371f
C2268 top_segment_2_0.rseg_2_v3_0.v9.t1 GND 0.0362f
C2269 top_segment_2_0.rseg_2_v3_0.v9.t2 GND 0.20214f
C2270 top_segment_2_0.rseg_2_v3_0.v9.n0 GND 4.25884f
C2271 top_segment_2_0.rseg_2_v3_0.v9.t0 GND 0.20281f
C2272 a_21026_19162.t1 GND 0.1868f
C2273 a_21026_19162.t2 GND 0.17175f
C2274 a_21026_19162.t3 GND 0.07075f
C2275 a_21026_19162.n0 GND 4.99847f
C2276 a_21026_19162.n1 GND 5.49565f
C2277 a_21026_19162.t0 GND 0.07658f
C2278 top_segment_4_1.bb1.t1 GND 0.09482f
C2279 top_segment_4_1.bb1.n0 GND 0.03888f
C2280 top_segment_4_1.bb1.n1 GND 0.08369f
C2281 top_segment_4_1.bb1.n2 GND 0.05556f
C2282 top_segment_4_1.bb1.t2 GND 0.18746f
C2283 top_segment_4_1.bb1.n3 GND 0.39156f
C2284 top_segment_4_1.bb1.t3 GND 0.18537f
C2285 top_segment_4_1.bb1.n4 GND 8.96447f
C2286 top_segment_4_1.bb1.t6 GND 0.17903f
C2287 top_segment_4_1.bb1.t5 GND 0.17637f
C2288 top_segment_4_1.bb1.n5 GND 1.89914f
C2289 top_segment_4_1.bb1.n6 GND 13.6142f
C2290 top_segment_4_1.bb1.t4 GND 0.3316f
C2291 top_segment_4_1.bb1.t7 GND 0.18395f
C2292 top_segment_4_1.bb1.n7 GND 0.28895f
C2293 top_segment_4_1.bb1.n8 GND 0.05749f
C2294 top_segment_4_1.bb1.n9 GND 0.08242f
C2295 top_segment_4_1.bb1.n10 GND 0.04698f
C2296 top_segment_4_1.bb1.t0 GND 0.09083f
C2297 a_35435_18774.t5 GND 0.03016f
C2298 a_35435_18774.t4 GND 0.14825f
C2299 a_35435_18774.n0 GND 0.16973f
C2300 a_35435_18774.t7 GND 0.15058f
C2301 a_35435_18774.n1 GND 0.279f
C2302 a_35435_18774.t6 GND 0.15058f
C2303 a_35435_18774.t2 GND 0.14825f
C2304 a_35435_18774.t3 GND 0.03016f
C2305 a_35435_18774.n2 GND 0.16973f
C2306 a_35435_18774.n3 GND 0.29912f
C2307 a_35435_18774.t0 GND 0.05237f
C2308 a_35435_18774.n4 GND 0.83928f
C2309 a_35435_18774.t1 GND 0.03278f
C2310 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t2 GND 0.02802f
C2311 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t3 GND 0.02802f
C2312 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n0 GND 0.06682f
C2313 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.Y GND 0.21666f
C2314 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n1 GND 0.13128f
C2315 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t4 GND 0.76823f
C2316 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n2 GND 16.1392f
C2317 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n3 GND 0.04085f
C2318 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t0 GND 0.04311f
C2319 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.t1 GND 0.04311f
C2320 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.IN.n4 GND 0.09469f
C2321 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t1 GND 0.04142f
C2322 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t2 GND 0.04142f
C2323 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n0 GND 0.09096f
C2324 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x1.Y GND 0.20814f
C2325 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n1 GND 0.03924f
C2326 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t5 GND 0.06443f
C2327 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t7 GND 0.03797f
C2328 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t6 GND 0.06443f
C2329 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t8 GND 0.03797f
C2330 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n2 GND 0.1081f
C2331 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n3 GND 0.16037f
C2332 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_10.x2.A GND 0.01074f
C2333 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n4 GND 0.04836f
C2334 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t4 GND 0.55071f
C2335 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n5 GND 15.822f
C2336 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n6 GND 0.02963f
C2337 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t3 GND 0.02692f
C2338 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.t0 GND 0.02692f
C2339 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n7 GND 0.06419f
C2340 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_1/lvsf_0.INB.n8 GND 0.12611f
C2341 top_segment_3_0.rseg_3_v3_0.v9.t1 GND 0.20441f
C2342 top_segment_3_0.rseg_3_v3_0.v9.t2 GND 0.03593f
C2343 top_segment_3_0.rseg_3_v3_0.v9.n0 GND 5.13537f
C2344 top_segment_3_0.rseg_3_v3_0.v9.t0 GND 0.22429f
C2345 top_segment_3_0.rseg_3_v3_0.v10.t1 GND 0.09859f
C2346 top_segment_3_0.rseg_3_v3_0.v10.t2 GND 0.01938f
C2347 top_segment_3_0.rseg_3_v3_0.v10.n0 GND 2.39212f
C2348 top_segment_3_0.rseg_3_v3_0.v10.t0 GND 0.08991f
C2349 a_33403_7938.t1 GND 0.10872f
C2350 a_33403_7938.t2 GND 0.13049f
C2351 a_33403_7938.n0 GND 6.09434f
C2352 a_33403_7938.t0 GND 0.06644f
C2353 a_22406_19162.t2 GND 0.06748f
C2354 a_22406_19162.t1 GND 0.053f
C2355 a_22406_19162.n0 GND 2.83277f
C2356 a_22406_19162.t3 GND 0.08959f
C2357 a_22406_19162.n1 GND 2.82036f
C2358 a_22406_19162.t0 GND 0.03679f
C2359 a_17271_7938.t2 GND 0.03667f
C2360 a_17271_7938.t1 GND 0.03722f
C2361 a_17271_7938.n0 GND 2.59201f
C2362 a_17271_7938.t0 GND 0.0341f
C2363 a_22176_17121.t1 GND 0.07067f
C2364 a_22176_17121.t2 GND 0.05945f
C2365 a_22176_17121.n0 GND 2.30243f
C2366 a_22176_17121.t5 GND 0.05945f
C2367 a_22176_17121.n1 GND 1.38823f
C2368 a_22176_17121.t4 GND 0.05945f
C2369 a_22176_17121.n2 GND 1.3619f
C2370 a_22176_17121.t3 GND 0.05907f
C2371 a_22176_17121.n3 GND 1.47888f
C2372 a_22176_17121.t0 GND 0.06045f
C2373 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t1 GND 0.01506f
C2374 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t2 GND 0.08868f
C2375 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.t0 GND 0.09157f
C2376 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v28.n0 GND 1.45797f
C2377 a_15162_6674.t3 GND 0.09282f
C2378 a_15162_6674.t2 GND 0.07318f
C2379 a_15162_6674.n0 GND 5.4585f
C2380 a_15162_6674.t1 GND 0.07318f
C2381 a_15162_6674.n1 GND 2.6889f
C2382 a_15162_6674.t4 GND 0.07479f
C2383 a_15162_6674.n2 GND 3.75672f
C2384 a_15162_6674.t0 GND 0.0819f
C2385 top_segment_3_0.b[6].t1 GND 0.09761f
C2386 top_segment_3_0.b[6].n0 GND 0.04002f
C2387 top_segment_3_0.b[6].n1 GND 0.08615f
C2388 top_segment_3_0.b[6].n2 GND 0.0572f
C2389 top_segment_3_0.b[6].t2 GND 0.19391f
C2390 top_segment_3_0.b[6].t7 GND 0.19298f
C2391 top_segment_3_0.b[6].n3 GND 0.605f
C2392 top_segment_3_0.b[6].t8 GND 0.19298f
C2393 top_segment_3_0.b[6].n4 GND 0.30296f
C2394 top_segment_3_0.b[6].t3 GND 0.19298f
C2395 top_segment_3_0.b[6].n5 GND 0.30296f
C2396 top_segment_3_0.b[6].t9 GND 0.19298f
C2397 top_segment_3_0.b[6].n6 GND 0.30296f
C2398 top_segment_3_0.b[6].t4 GND 0.19298f
C2399 top_segment_3_0.b[6].n7 GND 0.30296f
C2400 top_segment_3_0.b[6].t6 GND 0.19298f
C2401 top_segment_3_0.b[6].n8 GND 0.30296f
C2402 top_segment_3_0.b[6].t10 GND 0.19298f
C2403 top_segment_3_0.b[6].n9 GND 0.30296f
C2404 top_segment_3_0.b[6].t5 GND 0.19298f
C2405 top_segment_3_0.b[6].n10 GND 0.24595f
C2406 top_segment_3_0.b[6].n11 GND 15.8955f
C2407 top_segment_3_0.b[6].n12 GND 0.06157f
C2408 top_segment_3_0.b[6].t0 GND 0.09351f
C2409 top_segment_3_0.b[6].n13 GND 0.04837f
C2410 a_19646_19162.t1 GND 0.19205f
C2411 a_19646_19162.t3 GND 0.1673f
C2412 a_19646_19162.t2 GND 0.0575f
C2413 a_19646_19162.n0 GND 4.4887f
C2414 a_19646_19162.n1 GND 5.71483f
C2415 a_19646_19162.t0 GND 0.07964f
C2416 top_segment_2_0.DEC0[1].t17 GND 0.14561f
C2417 top_segment_2_0.DEC0[1].n0 GND 0.18624f
C2418 top_segment_2_0.DEC0[1].t7 GND 0.14561f
C2419 top_segment_2_0.DEC0[1].n1 GND 0.23751f
C2420 top_segment_2_0.DEC0[1].t21 GND 0.14561f
C2421 top_segment_2_0.DEC0[1].n2 GND 0.23751f
C2422 top_segment_2_0.DEC0[1].t9 GND 0.14561f
C2423 top_segment_2_0.DEC0[1].n3 GND 0.23751f
C2424 top_segment_2_0.DEC0[1].t5 GND 0.14561f
C2425 top_segment_2_0.DEC0[1].n4 GND 0.23751f
C2426 top_segment_2_0.DEC0[1].t15 GND 0.14561f
C2427 top_segment_2_0.DEC0[1].n5 GND 0.23751f
C2428 top_segment_2_0.DEC0[1].t8 GND 0.14561f
C2429 top_segment_2_0.DEC0[1].n6 GND 0.23751f
C2430 top_segment_2_0.DEC0[1].t19 GND 0.14561f
C2431 top_segment_2_0.DEC0[1].n7 GND 0.22308f
C2432 top_segment_2_0.DEC0[1].t4 GND 0.14635f
C2433 top_segment_2_0.DEC0[1].t11 GND 0.14561f
C2434 top_segment_2_0.DEC0[1].n8 GND 0.47428f
C2435 top_segment_2_0.DEC0[1].t2 GND 0.14561f
C2436 top_segment_2_0.DEC0[1].n9 GND 0.23751f
C2437 top_segment_2_0.DEC0[1].t14 GND 0.14561f
C2438 top_segment_2_0.DEC0[1].n10 GND 0.23751f
C2439 top_segment_2_0.DEC0[1].t18 GND 0.14561f
C2440 top_segment_2_0.DEC0[1].n11 GND 0.23751f
C2441 top_segment_2_0.DEC0[1].t3 GND 0.14561f
C2442 top_segment_2_0.DEC0[1].n12 GND 0.23751f
C2443 top_segment_2_0.DEC0[1].t16 GND 0.14561f
C2444 top_segment_2_0.DEC0[1].n13 GND 0.23751f
C2445 top_segment_2_0.DEC0[1].t6 GND 0.14561f
C2446 top_segment_2_0.DEC0[1].n14 GND 0.23751f
C2447 top_segment_2_0.DEC0[1].t13 GND 0.14561f
C2448 top_segment_2_0.DEC0[1].n15 GND 0.17196f
C2449 top_segment_2_0.DEC0[1].n16 GND 16.048f
C2450 top_segment_2_0.DEC0[1].t1 GND 0.1204f
C2451 top_segment_2_0.DEC0[1].t0 GND 0.10238f
C2452 top_segment_2_0.DEC0[1].n17 GND 0.82365f
C2453 top_segment_2_0.DEC0[1].t12 GND 0.47802f
C2454 top_segment_2_0.DEC0[1].t20 GND 0.47604f
C2455 top_segment_2_0.DEC0[1].n18 GND 0.75563f
C2456 top_segment_2_0.DEC0[1].n19 GND 0.48747f
C2457 top_segment_2_0.DEC0[1].t10 GND 0.50273f
C2458 top_segment_2_0.DEC0[1].n20 GND 1.05121f
C2459 a_29589_6674.t4 GND 0.10032f
C2460 a_29589_6674.t1 GND 0.08434f
C2461 a_29589_6674.n0 GND 3.60497f
C2462 a_29589_6674.t2 GND 0.07983f
C2463 a_29589_6674.n1 GND 2.75522f
C2464 a_29589_6674.t3 GND 0.14569f
C2465 a_29589_6674.n2 GND 5.84981f
C2466 a_29589_6674.t0 GND 0.07983f
C2467 top_segment_1_0.rseg_1_v3_1.v20.t2 GND -0.04304f
C2468 top_segment_1_0.rseg_1_v3_1.v20.t1 GND -0.04297f
C2469 top_segment_1_0.rseg_1_v3_1.v20.n0 GND -0.74314f
C2470 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t3 GND 0.0272f
C2471 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t2 GND 0.0272f
C2472 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n0 GND 0.06485f
C2473 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x1.Y GND 0.21025f
C2474 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n1 GND 0.1274f
C2475 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t13 GND 0.06508f
C2476 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t18 GND 0.03835f
C2477 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t11 GND 0.06508f
C2478 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t17 GND 0.03835f
C2479 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n2 GND 0.1092f
C2480 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n3 GND 0.162f
C2481 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.A GND 0.01085f
C2482 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n4 GND 0.04886f
C2483 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t9 GND 0.06917f
C2484 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t15 GND 0.04317f
C2485 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n5 GND 0.13623f
C2486 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.B GND 0.01674f
C2487 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n6 GND 0.06232f
C2488 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t20 GND 0.06917f
C2489 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t6 GND 0.04317f
C2490 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n7 GND 0.13618f
C2491 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.B GND 0.01715f
C2492 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n8 GND 0.046f
C2493 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n9 GND 0.71314f
C2494 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[0] GND 1.82836f
C2495 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t14 GND 0.25867f
C2496 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n10 GND 5.84879f
C2497 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x1/x1.B GND 0.01799f
C2498 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t16 GND 0.04317f
C2499 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t5 GND 0.06917f
C2500 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n11 GND 0.13609f
C2501 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n12 GND 0.12915f
C2502 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[6] GND 0.18f
C2503 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n13 GND 0.89598f
C2504 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t10 GND 0.07051f
C2505 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t7 GND 0.04428f
C2506 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n14 GND 0.09547f
C2507 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x2.C GND -0.02483f
C2508 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n15 GND 0.41728f
C2509 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n16 GND 1.14727f
C2510 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x5.A GND 0.01994f
C2511 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t12 GND 0.04344f
C2512 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t19 GND 0.06949f
C2513 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n17 GND 0.12217f
C2514 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n18 GND 0.19259f
C2515 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n19 GND 1.11131f
C2516 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t4 GND 0.04344f
C2517 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t8 GND 0.06949f
C2518 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n20 GND 0.12266f
C2519 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x8.A GND 0.01585f
C2520 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n21 GND 0.13712f
C2521 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n22 GND 5.41443f
C2522 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n23 GND 8.07493f
C2523 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n24 GND 1.01356f
C2524 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n25 GND 0.02993f
C2525 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n26 GND 0.03964f
C2526 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t1 GND 0.04184f
C2527 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.t0 GND 0.04184f
C2528 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.INB.n27 GND 0.09189f
C2529 top_segment_1_0.rseg_1_v3_1.v8.t1 GND 0.0341f
C2530 top_segment_1_0.rseg_1_v3_1.v8.t2 GND 0.12376f
C2531 top_segment_1_0.rseg_1_v3_1.v8.t0 GND 0.363f
C2532 top_segment_1_0.rseg_1_v3_1.v8.n0 GND 2.62718f
C2533 top_segment_2_0.rseg_2_v3_0.v36.t1 GND 0.09876f
C2534 top_segment_2_0.rseg_2_v3_0.v36.t2 GND 0.01345f
C2535 top_segment_2_0.rseg_2_v3_0.v36.n0 GND 1.88582f
C2536 top_segment_2_0.rseg_2_v3_0.v36.t0 GND 0.10196f
C2537 top_segment_2_0.rseg_2_v3_0.v40.t1 GND 0.16127f
C2538 top_segment_2_0.rseg_2_v3_0.v40.t2 GND 0.02546f
C2539 top_segment_2_0.rseg_2_v3_0.v40.n0 GND 4.57733f
C2540 top_segment_2_0.rseg_2_v3_0.v40.t0 GND 0.63594f
C2541 top_segment_2_0.rseg_2_v3_0.v23.t1 GND 0.09015f
C2542 top_segment_2_0.rseg_2_v3_0.v23.t2 GND 0.01519f
C2543 top_segment_2_0.rseg_2_v3_0.v23.n0 GND 1.90489f
C2544 top_segment_2_0.rseg_2_v3_0.v23.t0 GND 0.08977f
C2545 top_segment_2_0.rseg_2_v3_0.v22.t1 GND 0.0165f
C2546 top_segment_2_0.rseg_2_v3_0.v22.t2 GND 0.0952f
C2547 top_segment_2_0.rseg_2_v3_0.v22.n0 GND 2.09304f
C2548 top_segment_2_0.rseg_2_v3_0.v22.t0 GND 0.09527f
C2549 a_18493_7938.t2 GND 0.07897f
C2550 a_18493_7938.t1 GND 0.06395f
C2551 a_18493_7938.n0 GND 5.77629f
C2552 a_18493_7938.t0 GND 0.08079f
C2553 a_15438_6674.t3 GND 0.09293f
C2554 a_15438_6674.t2 GND 0.07283f
C2555 a_15438_6674.n0 GND 5.53481f
C2556 a_15438_6674.t1 GND 0.07283f
C2557 a_15438_6674.n1 GND 2.64424f
C2558 a_15438_6674.t4 GND 0.07429f
C2559 a_15438_6674.n2 GND 3.92477f
C2560 a_15438_6674.t0 GND 0.08331f
C2561 a_28879_6674.t4 GND 0.0892f
C2562 a_28879_6674.t1 GND 0.09588f
C2563 a_28879_6674.n0 GND 3.63616f
C2564 a_28879_6674.t2 GND 0.07875f
C2565 a_28879_6674.n1 GND 2.9429f
C2566 a_28879_6674.t3 GND 0.14222f
C2567 a_28879_6674.n2 GND 5.73614f
C2568 a_28879_6674.t0 GND 0.07875f
C2569 a_18099_7938.t2 GND 0.08071f
C2570 a_18099_7938.t1 GND 0.08167f
C2571 a_18099_7938.n0 GND 5.66782f
C2572 a_18099_7938.t0 GND 0.0698f
C2573 a_13154_5238.t1 GND 0.08343f
C2574 a_13154_5238.t2 GND 0.06448f
C2575 a_13154_5238.n0 GND 4.80455f
C2576 a_13154_5238.t4 GND 0.08172f
C2577 a_13154_5238.t3 GND 0.06448f
C2578 a_13154_5238.n1 GND 3.71167f
C2579 a_13154_5238.n2 GND 4.09447f
C2580 a_13154_5238.t0 GND 0.0952f
C2581 top_segment_2_0.rseg_2_v3_0.v1.t1 GND 0.01856f
C2582 top_segment_2_0.rseg_2_v3_0.v1.t2 GND 0.10649f
C2583 top_segment_2_0.rseg_2_v3_0.v1.n0 GND 1.95994f
C2584 top_segment_2_0.rseg_2_v3_0.v1.t0 GND 0.11501f
C2585 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t1 GND 0.01293f
C2586 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t2 GND 0.09801f
C2587 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.t0 GND 0.10101f
C2588 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v37.n0 GND 1.62769f
C2589 a_14452_6674.t3 GND 0.09398f
C2590 a_14452_6674.t2 GND 0.07505f
C2591 a_14452_6674.n0 GND 5.374f
C2592 a_14452_6674.t1 GND 0.07505f
C2593 a_14452_6674.n1 GND 2.89621f
C2594 a_14452_6674.t4 GND 0.08121f
C2595 a_14452_6674.n2 GND 3.82467f
C2596 a_14452_6674.t0 GND 0.07983f
C2597 a_17823_7938.t2 GND 0.07488f
C2598 a_17823_7938.t1 GND 0.07606f
C2599 a_17823_7938.n0 GND 5.28272f
C2600 a_17823_7938.t0 GND 0.06634f
C2601 top_segment_3_0.rseg_3_v3_0.v12.t1 GND 0.10511f
C2602 top_segment_3_0.rseg_3_v3_0.v12.t2 GND 0.10221f
C2603 top_segment_3_0.rseg_3_v3_0.v12.n0 GND 2.37213f
C2604 top_segment_3_0.rseg_3_v3_0.v12.t0 GND 0.02055f
C2605 top_segment_2_0.rseg_2_v3_0.v7.t1 GND 0.02493f
C2606 top_segment_2_0.rseg_2_v3_0.v7.t2 GND 0.09805f
C2607 top_segment_2_0.rseg_2_v3_0.v7.n0 GND 2.57844f
C2608 top_segment_2_0.rseg_2_v3_0.v7.t0 GND 0.09858f
C2609 top_segment_2_0.rseg_2_v3_0.v8.t1 GND 0.02096f
C2610 top_segment_2_0.rseg_2_v3_0.v8.t2 GND 0.52014f
C2611 top_segment_2_0.rseg_2_v3_0.v8.n0 GND 4.09913f
C2612 top_segment_2_0.rseg_2_v3_0.v8.t0 GND 0.15978f
C2613 top_segment_2_0.rseg_2_v3_0.v25.t1 GND 0.21167f
C2614 top_segment_2_0.rseg_2_v3_0.v25.t2 GND 0.03472f
C2615 top_segment_2_0.rseg_2_v3_0.v25.n0 GND 4.61554f
C2616 top_segment_2_0.rseg_2_v3_0.v25.t0 GND 0.23808f
C2617 top_segment_2_0.rseg_2_v3_0.v26.t2 GND 0.08819f
C2618 top_segment_2_0.rseg_2_v3_0.v26.t1 GND 0.09894f
C2619 top_segment_2_0.rseg_2_v3_0.v26.n0 GND 1.89904f
C2620 top_segment_2_0.rseg_2_v3_0.v26.t0 GND 0.01383f
C2621 a_27429_5238.t4 GND 0.14276f
C2622 a_27429_5238.t1 GND 0.08249f
C2623 a_27429_5238.n0 GND 4.59159f
C2624 a_27429_5238.t2 GND 0.15799f
C2625 a_27429_5238.n1 GND 4.32313f
C2626 a_27429_5238.t3 GND 0.17484f
C2627 a_27429_5238.n2 GND 6.44471f
C2628 a_27429_5238.t0 GND 0.08249f
C2629 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t3 GND 0.21159f
C2630 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t1 GND 0.22082f
C2631 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t0 GND 0.21829f
C2632 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n0 GND 2.05618f
C2633 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.n1 GND 0.68941f
C2634 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S4.t2 GND 0.43691f
C2635 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t0 GND 0.05358f
C2636 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t8 GND 0.85572f
C2637 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n0 GND 0.12606f
C2638 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t4 GND 0.08482f
C2639 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n1 GND 0.05712f
C2640 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t2 GND 0.08482f
C2641 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t5 GND 0.01718f
C2642 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n2 GND 0.1007f
C2643 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t3 GND 0.01718f
C2644 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n3 GND 0.13843f
C2645 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n4 GND 0.05663f
C2646 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t14 GND 0.12218f
C2647 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n5 GND 0.07605f
C2648 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t18 GND 0.12218f
C2649 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n6 GND 0.0851f
C2650 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t9 GND 0.12218f
C2651 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n7 GND 0.0851f
C2652 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t17 GND 0.12218f
C2653 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n8 GND 0.05779f
C2654 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t6 GND 0.12218f
C2655 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n9 GND 0.06025f
C2656 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t12 GND 0.12218f
C2657 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n10 GND 0.0851f
C2658 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t10 GND 0.12218f
C2659 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n11 GND 0.0851f
C2660 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t16 GND 0.12218f
C2661 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n12 GND 0.08168f
C2662 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t11 GND 0.12218f
C2663 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n13 GND 0.06025f
C2664 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t7 GND 0.12218f
C2665 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n14 GND 0.0851f
C2666 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t15 GND 0.12218f
C2667 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n15 GND 0.0851f
C2668 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t13 GND 0.12218f
C2669 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n16 GND 0.08168f
C2670 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n17 GND 0.27847f
C2671 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n18 GND 0.75769f
C2672 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n19 GND 0.13016f
C2673 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n20 GND 0.39284f
C2674 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n21 GND 0.26288f
C2675 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.t1 GND 0.05626f
C2676 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNDEC.n22 GND 0.23923f
C2677 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t5 GND 0.04207f
C2678 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t3 GND 0.04207f
C2679 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t4 GND 0.15904f
C2680 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t11 GND 0.16048f
C2681 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t12 GND 0.15996f
C2682 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n0 GND 0.19996f
C2683 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t9 GND 0.16046f
C2684 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t13 GND 0.15996f
C2685 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n1 GND 0.19556f
C2686 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n2 GND 0.04891f
C2687 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n3 GND 0.08386f
C2688 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t2 GND 0.15904f
C2689 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t1 GND 0.0423f
C2690 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t0 GND 0.04183f
C2691 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n4 GND 0.16659f
C2692 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t7 GND 0.15996f
C2693 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n5 GND 0.18631f
C2694 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t8 GND 0.15996f
C2695 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n6 GND 0.10596f
C2696 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t6 GND 0.16046f
C2697 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.t10 GND 0.15996f
C2698 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n7 GND 0.19556f
C2699 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n8 GND 0.04891f
C2700 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n9 GND 0.08386f
C2701 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n10 GND 0.06653f
C2702 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.D0.n11 GND 0.14113f
C2703 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t1 GND 0.01292f
C2704 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t2 GND 0.10105f
C2705 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.t0 GND 0.09788f
C2706 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v21.n0 GND 1.62825f
C2707 top_segment_2_0.rseg_2_v3_0.v43.t2 GND 0.01471f
C2708 top_segment_2_0.rseg_2_v3_0.v43.t1 GND 0.10178f
C2709 top_segment_2_0.rseg_2_v3_0.v43.n0 GND 2.07892f
C2710 top_segment_2_0.rseg_2_v3_0.v43.t0 GND 0.10459f
C2711 top_segment_2_0.rseg_2_v3_0.v44.t1 GND 0.10286f
C2712 top_segment_2_0.rseg_2_v3_0.v44.t2 GND 0.01467f
C2713 top_segment_2_0.rseg_2_v3_0.v44.n0 GND 2.07652f
C2714 top_segment_2_0.rseg_2_v3_0.v44.t0 GND 0.10595f
C2715 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t1 GND 0.03028f
C2716 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t3 GND 0.03028f
C2717 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n0 GND 0.06649f
C2718 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n1 GND 0.02868f
C2719 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t12 GND 0.0471f
C2720 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t9 GND 0.02775f
C2721 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t11 GND 0.0471f
C2722 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t8 GND 0.02775f
C2723 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n2 GND 0.07902f
C2724 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n3 GND 0.11723f
C2725 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n4 GND 0.03535f
C2726 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t13 GND 0.03129f
C2727 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t6 GND 0.05012f
C2728 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n5 GND 0.09554f
C2729 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n6 GND 0.15506f
C2730 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n7 GND 0.75373f
C2731 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t4 GND 0.03124f
C2732 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t7 GND 0.05005f
C2733 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n8 GND 0.09952f
C2734 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t10 GND 0.03129f
C2735 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t5 GND 0.05012f
C2736 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n9 GND 0.0954f
C2737 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n10 GND 0.01346f
C2738 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n11 GND 0.34761f
C2739 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n12 GND 8.72639f
C2740 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n13 GND 6.93802f
C2741 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n14 GND 0.02166f
C2742 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t0 GND 0.01968f
C2743 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].t2 GND 0.01968f
C2744 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n15 GND 0.04693f
C2745 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[9].n16 GND 0.09219f
C2746 a_26443_5238.t4 GND 0.13945f
C2747 a_26443_5238.t1 GND 0.0817f
C2748 a_26443_5238.n0 GND 5.49877f
C2749 a_26443_5238.t2 GND 0.17983f
C2750 a_26443_5238.n1 GND 4.84462f
C2751 a_26443_5238.t3 GND 0.17181f
C2752 a_26443_5238.n2 GND 5.30212f
C2753 a_26443_5238.t0 GND 0.0817f
C2754 top_segment_3_0.rseg_3_v3_0.v5.t2 GND 0.09431f
C2755 top_segment_3_0.rseg_3_v3_0.v5.t1 GND 0.01555f
C2756 top_segment_3_0.rseg_3_v3_0.v5.n0 GND 1.89943f
C2757 top_segment_3_0.rseg_3_v3_0.v5.t0 GND 0.09071f
C2758 top_segment_2_0.DEC1[0].t6 GND 0.16908f
C2759 top_segment_2_0.DEC1[0].t3 GND 0.16823f
C2760 top_segment_2_0.DEC1[0].n0 GND 0.50612f
C2761 top_segment_2_0.DEC1[0].t8 GND 0.16908f
C2762 top_segment_2_0.DEC1[0].t5 GND 0.16823f
C2763 top_segment_2_0.DEC1[0].n1 GND 0.54795f
C2764 top_segment_2_0.DEC1[0].n2 GND 0.13418f
C2765 top_segment_2_0.DEC1[0].t9 GND 0.16629f
C2766 top_segment_2_0.DEC1[0].n3 GND 15.1749f
C2767 top_segment_2_0.DEC1[0].t0 GND 0.13933f
C2768 top_segment_2_0.DEC1[0].t1 GND 0.11828f
C2769 top_segment_2_0.DEC1[0].n4 GND 1.15353f
C2770 top_segment_2_0.DEC1[0].t2 GND 0.55227f
C2771 top_segment_2_0.DEC1[0].t7 GND 0.54999f
C2772 top_segment_2_0.DEC1[0].n5 GND 0.91171f
C2773 top_segment_2_0.DEC1[0].t4 GND 0.54999f
C2774 top_segment_2_0.DEC1[0].n6 GND 0.47041f
C2775 top_segment_2_0.DEC1[0].n7 GND 0.86048f
C2776 top_segment_2_0.DEC1[3].t5 GND 0.16429f
C2777 top_segment_2_0.DEC1[3].t3 GND 0.16346f
C2778 top_segment_2_0.DEC1[3].n0 GND 0.47064f
C2779 top_segment_2_0.DEC1[3].t8 GND 0.16429f
C2780 top_segment_2_0.DEC1[3].t4 GND 0.16346f
C2781 top_segment_2_0.DEC1[3].n1 GND 0.53242f
C2782 top_segment_2_0.DEC1[3].n2 GND 0.15152f
C2783 top_segment_2_0.DEC1[3].t7 GND 0.16158f
C2784 top_segment_2_0.DEC1[3].n3 GND 15.2195f
C2785 top_segment_2_0.DEC1[3].t1 GND 0.13506f
C2786 top_segment_2_0.DEC1[3].t0 GND 0.11495f
C2787 top_segment_2_0.DEC1[3].n4 GND 0.69706f
C2788 top_segment_2_0.DEC1[3].t2 GND 0.53685f
C2789 top_segment_2_0.DEC1[3].t6 GND 0.53459f
C2790 top_segment_2_0.DEC1[3].n5 GND 0.89852f
C2791 top_segment_2_0.DEC1[3].t9 GND 0.53459f
C2792 top_segment_2_0.DEC1[3].n6 GND 0.78982f
C2793 top_segment_2_0.DEC1[3].n7 GND 1.21743f
C2794 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t2 GND 0.0223f
C2795 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t1 GND 0.12905f
C2796 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.t0 GND 0.42097f
C2797 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v56.n0 GND 2.85985f
C2798 top_segment_4_1.DEC3.t1 GND 0.08409f
C2799 top_segment_4_1.DEC3.n0 GND 0.03448f
C2800 top_segment_4_1.DEC3.n1 GND 0.07422f
C2801 top_segment_4_1.DEC3.n2 GND 0.04927f
C2802 top_segment_4_1.DEC3.t9 GND 0.16704f
C2803 top_segment_4_1.DEC3.t14 GND 0.16625f
C2804 top_segment_4_1.DEC3.n3 GND 0.52118f
C2805 top_segment_4_1.DEC3.t10 GND 0.16625f
C2806 top_segment_4_1.DEC3.n4 GND 0.26099f
C2807 top_segment_4_1.DEC3.t12 GND 0.16625f
C2808 top_segment_4_1.DEC3.n5 GND 0.26099f
C2809 top_segment_4_1.DEC3.t13 GND 0.16625f
C2810 top_segment_4_1.DEC3.n6 GND 0.26099f
C2811 top_segment_4_1.DEC3.t16 GND 0.16625f
C2812 top_segment_4_1.DEC3.n7 GND 0.26099f
C2813 top_segment_4_1.DEC3.t17 GND 0.16625f
C2814 top_segment_4_1.DEC3.n8 GND 0.26099f
C2815 top_segment_4_1.DEC3.t2 GND 0.16625f
C2816 top_segment_4_1.DEC3.n9 GND 0.2138f
C2817 top_segment_4_1.DEC3.t15 GND 0.16704f
C2818 top_segment_4_1.DEC3.t4 GND 0.16625f
C2819 top_segment_4_1.DEC3.n10 GND 0.52118f
C2820 top_segment_4_1.DEC3.t6 GND 0.16625f
C2821 top_segment_4_1.DEC3.n11 GND 0.26099f
C2822 top_segment_4_1.DEC3.t7 GND 0.16625f
C2823 top_segment_4_1.DEC3.n12 GND 0.21681f
C2824 top_segment_4_1.DEC3.t8 GND 0.16704f
C2825 top_segment_4_1.DEC3.t11 GND 0.16625f
C2826 top_segment_4_1.DEC3.n13 GND 0.52118f
C2827 top_segment_4_1.DEC3.t5 GND 0.16625f
C2828 top_segment_4_1.DEC3.n14 GND 0.26099f
C2829 top_segment_4_1.DEC3.t3 GND 0.16625f
C2830 top_segment_4_1.DEC3.n15 GND 0.21681f
C2831 top_segment_4_1.DEC3.n16 GND 0.2093f
C2832 top_segment_4_1.DEC3.n17 GND 16.7136f
C2833 top_segment_4_1.DEC3.n18 GND 0.07943f
C2834 top_segment_4_1.DEC3.t0 GND 0.08056f
C2835 top_segment_4_1.DEC3.n19 GND 0.04167f
C2836 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t1 GND 0.05407f
C2837 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t2 GND 0.03615f
C2838 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t3 GND 0.02256f
C2839 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n0 GND 0.07188f
C2840 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t4 GND 0.0362f
C2841 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t5 GND 0.0226f
C2842 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n1 GND 0.06891f
C2843 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n2 GND 0.02012f
C2844 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n3 GND 4.68779f
C2845 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].t0 GND 0.07769f
C2846 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n4 GND 0.107f
C2847 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[1].n5 GND 0.02567f
C2848 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t1 GND 0.05236f
C2849 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t8 GND 0.04377f
C2850 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t9 GND 0.02732f
C2851 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n0 GND 0.08703f
C2852 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t6 GND 0.04383f
C2853 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t7 GND 0.02737f
C2854 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n1 GND 0.08343f
C2855 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n2 GND 0.01642f
C2856 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n3 GND 0.0358f
C2857 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n4 GND 5.85791f
C2858 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t4 GND 0.04386f
C2859 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t5 GND 0.02739f
C2860 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n5 GND 0.0822f
C2861 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n6 GND 0.02224f
C2862 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n7 GND 0.2998f
C2863 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n8 GND 0.13919f
C2864 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t2 GND 0.02648f
C2865 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t3 GND 0.02648f
C2866 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n9 GND 0.05886f
C2867 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].t0 GND 0.12167f
C2868 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[1].n10 GND 0.29364f
C2869 top_segment_2_0.rseg_2_v3_0.v39.t1 GND 0.10272f
C2870 top_segment_2_0.rseg_2_v3_0.v39.t2 GND 0.01601f
C2871 top_segment_2_0.rseg_2_v3_0.v39.n0 GND 2.08049f
C2872 top_segment_2_0.rseg_2_v3_0.v39.t0 GND 0.10078f
C2873 a_23510_19162.t1 GND 0.15594f
C2874 a_23510_19162.t3 GND 0.06377f
C2875 a_23510_19162.n0 GND 5.11593f
C2876 a_23510_19162.t2 GND 0.10224f
C2877 a_23510_19162.n1 GND 3.89706f
C2878 a_23510_19162.t0 GND 0.06506f
C2879 top_segment_2_0.DEC0[2].t2 GND 0.14295f
C2880 top_segment_2_0.DEC0[2].t14 GND 0.14218f
C2881 top_segment_2_0.DEC0[2].n0 GND 0.50006f
C2882 top_segment_2_0.DEC0[2].t11 GND 0.14218f
C2883 top_segment_2_0.DEC0[2].n1 GND 0.25042f
C2884 top_segment_2_0.DEC0[2].t19 GND 0.14218f
C2885 top_segment_2_0.DEC0[2].n2 GND 0.22448f
C2886 top_segment_2_0.DEC0[2].t13 GND 0.14218f
C2887 top_segment_2_0.DEC0[2].n3 GND 0.19854f
C2888 top_segment_2_0.DEC0[2].t21 GND 0.14218f
C2889 top_segment_2_0.DEC0[2].n4 GND 0.25042f
C2890 top_segment_2_0.DEC0[2].t17 GND 0.14218f
C2891 top_segment_2_0.DEC0[2].n5 GND 0.25042f
C2892 top_segment_2_0.DEC0[2].t12 GND 0.14218f
C2893 top_segment_2_0.DEC0[2].n6 GND 0.23356f
C2894 top_segment_2_0.DEC0[2].t4 GND 0.14295f
C2895 top_segment_2_0.DEC0[2].t20 GND 0.14218f
C2896 top_segment_2_0.DEC0[2].n7 GND 0.50006f
C2897 top_segment_2_0.DEC0[2].t5 GND 0.14218f
C2898 top_segment_2_0.DEC0[2].n8 GND 0.25042f
C2899 top_segment_2_0.DEC0[2].t8 GND 0.14218f
C2900 top_segment_2_0.DEC0[2].n9 GND 0.25042f
C2901 top_segment_2_0.DEC0[2].t6 GND 0.14218f
C2902 top_segment_2_0.DEC0[2].n10 GND 0.25042f
C2903 top_segment_2_0.DEC0[2].t15 GND 0.14218f
C2904 top_segment_2_0.DEC0[2].n11 GND 0.25042f
C2905 top_segment_2_0.DEC0[2].t10 GND 0.14218f
C2906 top_segment_2_0.DEC0[2].n12 GND 0.25042f
C2907 top_segment_2_0.DEC0[2].t9 GND 0.14218f
C2908 top_segment_2_0.DEC0[2].n13 GND 0.25042f
C2909 top_segment_2_0.DEC0[2].t16 GND 0.14218f
C2910 top_segment_2_0.DEC0[2].n14 GND 0.1892f
C2911 top_segment_2_0.DEC0[2].n15 GND 14.7419f
C2912 top_segment_2_0.DEC0[2].t18 GND 0.4559f
C2913 top_segment_2_0.DEC0[2].t1 GND 0.09968f
C2914 top_segment_2_0.DEC0[2].t0 GND 0.11713f
C2915 top_segment_2_0.DEC0[2].n16 GND 0.6449f
C2916 top_segment_2_0.DEC0[2].n17 GND 0.51336f
C2917 top_segment_2_0.DEC0[2].t7 GND 0.46557f
C2918 top_segment_2_0.DEC0[2].t3 GND 0.46361f
C2919 top_segment_2_0.DEC0[2].n18 GND 1.03065f
C2920 top_segment_2_0.DEC0[2].n19 GND 0.7664f
C2921 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t3 GND 0.02821f
C2922 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t2 GND 0.02821f
C2923 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n0 GND 0.06728f
C2924 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n1 GND 0.13217f
C2925 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t13 GND 0.07176f
C2926 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t16 GND 0.04479f
C2927 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n2 GND 0.14268f
C2928 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t4 GND 0.07186f
C2929 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t8 GND 0.04486f
C2930 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n3 GND 0.13678f
C2931 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n4 GND 0.02691f
C2932 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n5 GND 0.06791f
C2933 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t9 GND 0.04479f
C2934 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t14 GND 0.07176f
C2935 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n6 GND 0.14129f
C2936 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n7 GND 0.19926f
C2937 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n8 GND 0.69128f
C2938 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t10 GND 0.07196f
C2939 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t7 GND 0.04495f
C2940 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n9 GND 0.13234f
C2941 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n10 GND 0.10406f
C2942 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n11 GND 0.77672f
C2943 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t15 GND 0.04479f
C2944 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t6 GND 0.07176f
C2945 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n12 GND 0.14129f
C2946 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n13 GND 0.19036f
C2947 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n14 GND 0.75233f
C2948 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t11 GND 0.07186f
C2949 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t12 GND 0.04486f
C2950 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n15 GND 0.13678f
C2951 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n16 GND 0.30498f
C2952 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n17 GND 1.04101f
C2953 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t17 GND 0.04479f
C2954 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t5 GND 0.07176f
C2955 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n18 GND 0.14124f
C2956 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n19 GND 0.13864f
C2957 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n20 GND 4.55762f
C2958 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n21 GND 12.0001f
C2959 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n22 GND 0.56248f
C2960 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n23 GND 0.04112f
C2961 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t0 GND 0.04341f
C2962 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].t1 GND 0.04341f
C2963 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[1].n24 GND 0.09533f
C2964 top_segment_1_0.rseg_1_v3_1.v25.t0 GND 0.04645f
C2965 top_segment_1_0.rseg_1_v3_1.v25.t2 GND 0.13937f
C2966 top_segment_1_0.rseg_1_v3_1.v25.t1 GND 0.14921f
C2967 top_segment_1_0.rseg_1_v3_1.v25.n0 GND 2.57872f
C2968 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t3 GND 0.02481f
C2969 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t2 GND 0.02481f
C2970 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n0 GND 0.05916f
C2971 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x2.Y GND 0.1918f
C2972 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n1 GND 0.11622f
C2973 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.A GND 0.01088f
C2974 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t8 GND 0.06318f
C2975 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t4 GND 0.03945f
C2976 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n2 GND 0.12027f
C2977 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n3 GND 0.07308f
C2978 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.A GND 0.01088f
C2979 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t5 GND 0.06318f
C2980 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t7 GND 0.03945f
C2981 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n4 GND 0.12027f
C2982 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n5 GND 0.03223f
C2983 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n6 GND 0.66246f
C2984 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.b[0] GND 2.72474f
C2985 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t6 GND 0.23963f
C2986 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n7 GND 11.603f
C2987 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n8 GND 1.68418f
C2988 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n9 GND 0.03616f
C2989 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t1 GND 0.03817f
C2990 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.t0 GND 0.03817f
C2991 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.IN.n10 GND 0.08382f
C2992 top_segment_3_0.b[4].t1 GND 0.10561f
C2993 top_segment_3_0.b[4].n0 GND 0.0433f
C2994 top_segment_3_0.b[4].n1 GND 0.09321f
C2995 top_segment_3_0.b[4].n2 GND 0.06188f
C2996 top_segment_3_0.b[4].t2 GND 0.20879f
C2997 top_segment_3_0.b[4].n3 GND 0.27086f
C2998 top_segment_3_0.b[4].t3 GND 0.20979f
C2999 top_segment_3_0.b[4].n4 GND 0.545f
C3000 top_segment_3_0.b[4].t4 GND 0.20647f
C3001 top_segment_3_0.b[4].n5 GND 15.6438f
C3002 top_segment_3_0.b[4].n6 GND 0.06662f
C3003 top_segment_3_0.b[4].t0 GND 0.10117f
C3004 top_segment_3_0.b[4].n7 GND 0.05233f
C3005 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t1 GND 0.02948f
C3006 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t2 GND 0.02948f
C3007 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n0 GND 0.07028f
C3008 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n1 GND 0.13808f
C3009 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t10 GND 0.07054f
C3010 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t7 GND 0.04157f
C3011 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t4 GND 0.07054f
C3012 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t13 GND 0.04157f
C3013 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n2 GND 0.11836f
C3014 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n3 GND 0.17559f
C3015 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n4 GND 0.05295f
C3016 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t8 GND 0.04679f
C3017 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t12 GND 0.07497f
C3018 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n5 GND 0.14751f
C3019 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n6 GND 0.23906f
C3020 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n7 GND 1.13361f
C3021 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t6 GND 0.04687f
C3022 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t11 GND 0.07507f
C3023 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n8 GND 0.14345f
C3024 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n9 GND 0.63171f
C3025 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n10 GND 1.9824f
C3026 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t5 GND 0.04689f
C3027 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t9 GND 0.07509f
C3028 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n11 GND 0.14293f
C3029 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n12 GND 0.27598f
C3030 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n13 GND 12.0537f
C3031 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n14 GND 9.98745f
C3032 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n15 GND 0.03244f
C3033 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n16 GND 0.04296f
C3034 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t3 GND 0.04535f
C3035 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].t0 GND 0.04535f
C3036 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.bb[8].n17 GND 0.09959f
C3037 top_segment_2_0.rseg_2_v3_0.v6.t2 GND 0.08522f
C3038 top_segment_2_0.rseg_2_v3_0.v6.t1 GND 0.01499f
C3039 top_segment_2_0.rseg_2_v3_0.v6.n0 GND 2.01508f
C3040 top_segment_2_0.rseg_2_v3_0.v6.t0 GND 0.08471f
C3041 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t0 GND 0.02742f
C3042 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t1 GND 0.15083f
C3043 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.t2 GND 0.16899f
C3044 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v25.n0 GND 2.83612f
C3045 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t0 GND 0.02265f
C3046 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t2 GND 0.13251f
C3047 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.t1 GND 0.39729f
C3048 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v24.n0 GND 2.76756f
C3049 a_13900_6674.t3 GND 0.03957f
C3050 a_13900_6674.t4 GND 0.04498f
C3051 a_13900_6674.n0 GND 2.05844f
C3052 a_13900_6674.t2 GND 0.04733f
C3053 a_13900_6674.t1 GND 0.03831f
C3054 a_13900_6674.n1 GND 2.62168f
C3055 a_13900_6674.n2 GND 1.51138f
C3056 a_13900_6674.t0 GND 0.03831f
C3057 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t1 GND 0.07426f
C3058 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t4 GND 0.04735f
C3059 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t5 GND 0.02955f
C3060 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n0 GND 0.09326f
C3061 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n1 GND 0.04267f
C3062 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t2 GND 0.04735f
C3063 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t3 GND 0.02955f
C3064 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n2 GND 0.09323f
C3065 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n3 GND 0.03149f
C3066 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n4 GND 0.48165f
C3067 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n5 GND 5.99489f
C3068 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n6 GND 0.25011f
C3069 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].n7 GND 0.02569f
C3070 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.bb[0].t0 GND 0.10587f
C3071 top_segment_3_0.bb[5].t1 GND 0.08958f
C3072 top_segment_3_0.bb[5].n0 GND 0.03673f
C3073 top_segment_3_0.bb[5].n1 GND 0.07907f
C3074 top_segment_3_0.bb[5].n2 GND 0.05249f
C3075 top_segment_3_0.bb[5].t3 GND 0.17711f
C3076 top_segment_3_0.bb[5].n3 GND 0.21367f
C3077 top_segment_3_0.bb[5].t5 GND 0.17796f
C3078 top_segment_3_0.bb[5].t6 GND 0.17711f
C3079 top_segment_3_0.bb[5].n4 GND 0.55525f
C3080 top_segment_3_0.bb[5].t4 GND 0.17711f
C3081 top_segment_3_0.bb[5].n5 GND 0.27805f
C3082 top_segment_3_0.bb[5].n6 GND 0.1851f
C3083 top_segment_3_0.bb[5].t8 GND 0.17514f
C3084 top_segment_3_0.bb[5].n7 GND 13.1384f
C3085 top_segment_3_0.bb[5].t7 GND 0.31329f
C3086 top_segment_3_0.bb[5].t2 GND 0.1738f
C3087 top_segment_3_0.bb[5].n8 GND 0.273f
C3088 top_segment_3_0.bb[5].n9 GND 0.05431f
C3089 top_segment_3_0.bb[5].n10 GND 0.07787f
C3090 top_segment_3_0.bb[5].n11 GND 0.04439f
C3091 top_segment_3_0.bb[5].t0 GND 0.08582f
C3092 a_14416_5238.t1 GND 0.04927f
C3093 a_14416_5238.t2 GND 0.03722f
C3094 a_14416_5238.n0 GND 2.56635f
C3095 a_14416_5238.t4 GND 0.04824f
C3096 a_14416_5238.t3 GND 0.03722f
C3097 a_14416_5238.n1 GND 2.76876f
C3098 a_14416_5238.n2 GND 1.74851f
C3099 a_14416_5238.t0 GND 0.04443f
C3100 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t1 GND 0.01247f
C3101 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t2 GND 0.09059f
C3102 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.t0 GND 0.08855f
C3103 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v23.n0 GND 1.58122f
C3104 top_segment_4_1.DEC1.t1 GND 0.08516f
C3105 top_segment_4_1.DEC1.n0 GND 0.03492f
C3106 top_segment_4_1.DEC1.n1 GND 0.07516f
C3107 top_segment_4_1.DEC1.n2 GND 0.0499f
C3108 top_segment_4_1.DEC1.t11 GND 0.16917f
C3109 top_segment_4_1.DEC1.t5 GND 0.16836f
C3110 top_segment_4_1.DEC1.n3 GND 0.52781f
C3111 top_segment_4_1.DEC1.t14 GND 0.16836f
C3112 top_segment_4_1.DEC1.n4 GND 0.26431f
C3113 top_segment_4_1.DEC1.t16 GND 0.16836f
C3114 top_segment_4_1.DEC1.n5 GND 0.26431f
C3115 top_segment_4_1.DEC1.t12 GND 0.16836f
C3116 top_segment_4_1.DEC1.n6 GND 0.26431f
C3117 top_segment_4_1.DEC1.t13 GND 0.16836f
C3118 top_segment_4_1.DEC1.n7 GND 0.26431f
C3119 top_segment_4_1.DEC1.t15 GND 0.16836f
C3120 top_segment_4_1.DEC1.n8 GND 0.26431f
C3121 top_segment_4_1.DEC1.t3 GND 0.16649f
C3122 top_segment_4_1.DEC1.t2 GND 0.16917f
C3123 top_segment_4_1.DEC1.t9 GND 0.16969f
C3124 top_segment_4_1.DEC1.t7 GND 0.16882f
C3125 top_segment_4_1.DEC1.n9 GND 0.57115f
C3126 top_segment_4_1.DEC1.t6 GND 0.16882f
C3127 top_segment_4_1.DEC1.n10 GND 0.28601f
C3128 top_segment_4_1.DEC1.t10 GND 0.16882f
C3129 top_segment_4_1.DEC1.n11 GND 0.28601f
C3130 top_segment_4_1.DEC1.t8 GND 0.16882f
C3131 top_segment_4_1.DEC1.n12 GND 0.28601f
C3132 top_segment_4_1.DEC1.t17 GND 0.16882f
C3133 top_segment_4_1.DEC1.n13 GND 0.28601f
C3134 top_segment_4_1.DEC1.n14 GND 0.43945f
C3135 top_segment_4_1.DEC1.t4 GND 0.16649f
C3136 top_segment_4_1.DEC1.n15 GND 0.42862f
C3137 top_segment_4_1.DEC1.n16 GND 0.20782f
C3138 top_segment_4_1.DEC1.n17 GND 13.6678f
C3139 top_segment_4_1.DEC1.n18 GND 13.4839f
C3140 top_segment_4_1.DEC1.n19 GND 0.06924f
C3141 top_segment_4_1.DEC1.t0 GND 0.08158f
C3142 top_segment_4_1.DEC1.n20 GND 0.0422f
C3143 top_segment_1_0.rseg_1_v3_1.v10.t1 GND 0.01319f
C3144 top_segment_1_0.rseg_1_v3_1.v10.t0 GND 0.03696f
C3145 top_segment_1_0.rseg_1_v3_1.v10.t2 GND 0.0369f
C3146 top_segment_1_0.rseg_1_v3_1.v10.n0 GND 0.66059f
C3147 top_segment_4_1.b1.t0 GND 0.09468f
C3148 top_segment_4_1.b1.n0 GND 0.03882f
C3149 top_segment_4_1.b1.n1 GND 0.08356f
C3150 top_segment_4_1.b1.n2 GND 0.05548f
C3151 top_segment_4_1.b1.t1 GND 0.0907f
C3152 top_segment_4_1.b1.n3 GND 0.01146f
C3153 top_segment_4_1.b1.t4 GND 0.18808f
C3154 top_segment_4_1.b1.n4 GND 0.42232f
C3155 top_segment_4_1.b1.t5 GND 0.1851f
C3156 top_segment_4_1.b1.n5 GND 8.8209f
C3157 top_segment_4_1.b1.t2 GND 0.17858f
C3158 top_segment_4_1.b1.t3 GND 0.17611f
C3159 top_segment_4_1.b1.n6 GND 1.94256f
C3160 top_segment_4_1.b1.n7 GND 13.6325f
C3161 top_segment_4_1.b1.n8 GND 0.05972f
C3162 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/sky130_fd_sc_hvl__inv_1_3.Y GND 0.48818f
C3163 top_segment_4_1.DEC0.t1 GND 0.08559f
C3164 top_segment_4_1.DEC0.n0 GND 0.03509f
C3165 top_segment_4_1.DEC0.n1 GND 0.07555f
C3166 top_segment_4_1.DEC0.n2 GND 0.05016f
C3167 top_segment_4_1.DEC0.t5 GND 0.17003f
C3168 top_segment_4_1.DEC0.t15 GND 0.16922f
C3169 top_segment_4_1.DEC0.n3 GND 0.53051f
C3170 top_segment_4_1.DEC0.t9 GND 0.16922f
C3171 top_segment_4_1.DEC0.n4 GND 0.26566f
C3172 top_segment_4_1.DEC0.t11 GND 0.16922f
C3173 top_segment_4_1.DEC0.n5 GND 0.22069f
C3174 top_segment_4_1.DEC0.t17 GND 0.17003f
C3175 top_segment_4_1.DEC0.t16 GND 0.16922f
C3176 top_segment_4_1.DEC0.n6 GND 0.53051f
C3177 top_segment_4_1.DEC0.t8 GND 0.16922f
C3178 top_segment_4_1.DEC0.n7 GND 0.26566f
C3179 top_segment_4_1.DEC0.t14 GND 0.16922f
C3180 top_segment_4_1.DEC0.n8 GND 0.22069f
C3181 top_segment_4_1.DEC0.n9 GND 0.64939f
C3182 top_segment_4_1.DEC0.t6 GND 0.16922f
C3183 top_segment_4_1.DEC0.n10 GND 1.05429f
C3184 top_segment_4_1.DEC0.t12 GND 0.16922f
C3185 top_segment_4_1.DEC0.n11 GND 0.26566f
C3186 top_segment_4_1.DEC0.t10 GND 0.16922f
C3187 top_segment_4_1.DEC0.n12 GND 0.26566f
C3188 top_segment_4_1.DEC0.t7 GND 0.16922f
C3189 top_segment_4_1.DEC0.n13 GND 0.26566f
C3190 top_segment_4_1.DEC0.t13 GND 0.16922f
C3191 top_segment_4_1.DEC0.n14 GND 0.26566f
C3192 top_segment_4_1.DEC0.t3 GND 0.16922f
C3193 top_segment_4_1.DEC0.n15 GND 0.26566f
C3194 top_segment_4_1.DEC0.t2 GND 0.16922f
C3195 top_segment_4_1.DEC0.n16 GND 0.26566f
C3196 top_segment_4_1.DEC0.t4 GND 0.16922f
C3197 top_segment_4_1.DEC0.n17 GND 14.7335f
C3198 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dec2b[0] GND 0.13752f
C3199 top_segment_4_1.DEC0.n18 GND 12.4597f
C3200 top_segment_4_1.DEC0.n19 GND 0.06984f
C3201 top_segment_4_1.DEC0.t0 GND 0.082f
C3202 top_segment_4_1.DEC0.n20 GND 0.04241f
C3203 a_19045_7938.t2 GND 0.04106f
C3204 a_19045_7938.t1 GND 0.03172f
C3205 a_19045_7938.n0 GND 2.9852f
C3206 a_19045_7938.t0 GND 0.04203f
C3207 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t2 GND 0.01441f
C3208 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t1 GND 0.08695f
C3209 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.t0 GND 0.07745f
C3210 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v26.n0 GND 1.43576f
C3211 a_29155_6674.t4 GND 0.0933f
C3212 a_29155_6674.t1 GND 0.08812f
C3213 a_29155_6674.n0 GND 3.52034f
C3214 a_29155_6674.t2 GND 0.07942f
C3215 a_29155_6674.n1 GND 2.88984f
C3216 a_29155_6674.t3 GND 0.14424f
C3217 a_29155_6674.n2 GND 5.80531f
C3218 a_29155_6674.t0 GND 0.07942f
C3219 a_33679_7938.t1 GND 0.05535f
C3220 a_33679_7938.t2 GND 0.06636f
C3221 a_33679_7938.n0 GND 3.04622f
C3222 a_33679_7938.t0 GND 0.03208f
C3223 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t4 GND 0.15112f
C3224 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n0 GND 0.31314f
C3225 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t5 GND 0.03061f
C3226 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n1 GND 0.09861f
C3227 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t17 GND 0.19802f
C3228 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n3 GND 0.13878f
C3229 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t10 GND 0.19802f
C3230 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n4 GND 0.14564f
C3231 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t13 GND 0.19802f
C3232 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n5 GND 0.14564f
C3233 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t15 GND 0.19802f
C3234 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n6 GND 0.10675f
C3235 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t11 GND 0.19802f
C3236 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n7 GND 0.10675f
C3237 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t9 GND 0.19802f
C3238 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n8 GND 0.14564f
C3239 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t12 GND 0.19802f
C3240 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n9 GND 0.14564f
C3241 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t7 GND 0.19802f
C3242 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n10 GND 0.14408f
C3243 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t8 GND 0.19802f
C3244 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n11 GND 0.10675f
C3245 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t16 GND 0.19802f
C3246 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n12 GND 0.14564f
C3247 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t6 GND 0.19802f
C3248 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n13 GND 0.14564f
C3249 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t14 GND 0.19802f
C3250 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n14 GND 0.10859f
C3251 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n15 GND 0.39639f
C3252 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n16 GND 0.8517f
C3253 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t3 GND 0.03061f
C3254 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n17 GND 0.08691f
C3255 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t2 GND 0.15112f
C3256 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n18 GND 0.11384f
C3257 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n19 GND 0.67032f
C3258 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t0 GND 0.09915f
C3259 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n20 GND 0.53323f
C3260 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.t1 GND 0.09577f
C3261 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPDEC.n21 GND 0.14399f
C3262 a_19922_19162.t2 GND 0.11548f
C3263 a_19922_19162.t3 GND 0.04818f
C3264 a_19922_19162.n0 GND 3.58176f
C3265 a_19922_19162.t1 GND 0.03156f
C3266 a_19922_19162.n1 GND 2.4369f
C3267 a_19922_19162.t0 GND 0.08612f
C3268 top_segment_4_1.b3.t1 GND 0.07211f
C3269 top_segment_4_1.b3.n0 GND 0.02957f
C3270 top_segment_4_1.b3.n1 GND 0.06365f
C3271 top_segment_4_1.b3.n2 GND 0.04226f
C3272 top_segment_4_1.b3.t3 GND 0.14257f
C3273 top_segment_4_1.b3.n3 GND 0.1747f
C3274 top_segment_4_1.b3.t18 GND 0.14257f
C3275 top_segment_4_1.b3.n4 GND 0.22382f
C3276 top_segment_4_1.b3.t7 GND 0.14257f
C3277 top_segment_4_1.b3.n5 GND 0.22382f
C3278 top_segment_4_1.b3.t11 GND 0.14257f
C3279 top_segment_4_1.b3.n6 GND 0.22382f
C3280 top_segment_4_1.b3.t4 GND 0.14257f
C3281 top_segment_4_1.b3.n7 GND 0.22382f
C3282 top_segment_4_1.b3.t6 GND 0.14257f
C3283 top_segment_4_1.b3.n8 GND 0.22382f
C3284 top_segment_4_1.b3.t16 GND 0.14325f
C3285 top_segment_4_1.b3.n9 GND 0.37214f
C3286 top_segment_4_1.b3.t10 GND 0.14098f
C3287 top_segment_4_1.b3.n10 GND 2.18424f
C3288 top_segment_4_1.b3.t15 GND 0.14325f
C3289 top_segment_4_1.b3.n11 GND 0.33381f
C3290 top_segment_4_1.b3.t2 GND 0.14098f
C3291 top_segment_4_1.b3.n12 GND 2.06846f
C3292 top_segment_4_1.b3.n13 GND 9.29285f
C3293 top_segment_4_1.b3.t19 GND 0.13639f
C3294 top_segment_4_1.b3.t9 GND 0.1357f
C3295 top_segment_4_1.b3.n14 GND 0.44201f
C3296 top_segment_4_1.b3.t13 GND 0.1357f
C3297 top_segment_4_1.b3.n15 GND 0.22135f
C3298 top_segment_4_1.b3.t5 GND 0.1357f
C3299 top_segment_4_1.b3.n16 GND 0.22135f
C3300 top_segment_4_1.b3.t8 GND 0.1357f
C3301 top_segment_4_1.b3.n17 GND 0.22135f
C3302 top_segment_4_1.b3.t14 GND 0.13588f
C3303 top_segment_4_1.b3.t17 GND 0.1357f
C3304 top_segment_4_1.b3.n18 GND 0.19705f
C3305 top_segment_4_1.b3.n19 GND 0.149f
C3306 top_segment_4_1.b3.t12 GND 0.13414f
C3307 top_segment_4_1.b3.n20 GND 1.98463f
C3308 top_segment_4_1.b3.n21 GND 8.77348f
C3309 top_segment_4_1.b3.n22 GND 0.04549f
C3310 top_segment_4_1.b3.t0 GND 0.06908f
C3311 top_segment_4_1.b3.n23 GND 0.03573f
C3312 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t0 GND 0.39374f
C3313 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t3 GND 0.19462f
C3314 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t2 GND 0.21619f
C3315 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n0 GND 1.60492f
C3316 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.t1 GND 0.20263f
C3317 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S1.n1 GND 3.37677f
C3318 a_18217_7938.t2 GND 0.0805f
C3319 a_18217_7938.t1 GND 0.06677f
C3320 a_18217_7938.n0 GND 5.8709f
C3321 a_18217_7938.t0 GND 0.08183f
C3322 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t1 GND 0.02431f
C3323 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t2 GND 0.02431f
C3324 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n0 GND 0.05796f
C3325 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_2.x2.Y GND 0.18793f
C3326 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n1 GND 0.11387f
C3327 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_3.A GND 0.01066f
C3328 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t13 GND 0.0619f
C3329 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t18 GND 0.03865f
C3330 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n2 GND 0.11784f
C3331 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n3 GND 0.07161f
C3332 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.dec_logic_0/sky130_fd_sc_hd__nand2_1_1.A GND 0.01066f
C3333 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t4 GND 0.0619f
C3334 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t7 GND 0.03865f
C3335 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n4 GND 0.11784f
C3336 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n5 GND 0.03158f
C3337 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n6 GND 0.64907f
C3338 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.b[0] GND 1.66982f
C3339 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t17 GND 0.23188f
C3340 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n7 GND 5.28977f
C3341 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[6] GND 0.11568f
C3342 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t8 GND 0.03865f
C3343 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t14 GND 0.0619f
C3344 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n8 GND 0.118f
C3345 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x2.A GND 0.0167f
C3346 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n9 GND 0.21334f
C3347 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n10 GND 0.62504f
C3348 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t15 GND 0.06302f
C3349 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t10 GND 0.03957f
C3350 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n11 GND 0.09737f
C3351 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x1.B GND 0.03102f
C3352 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n12 GND 0.34887f
C3353 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n13 GND 0.85432f
C3354 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t16 GND 0.03865f
C3355 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t6 GND 0.0619f
C3356 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n14 GND 0.11826f
C3357 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x2/x3.A GND 0.01299f
C3358 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n15 GND 0.25368f
C3359 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n16 GND 0.89808f
C3360 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x2.A GND 0.01066f
C3361 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t11 GND 0.0619f
C3362 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t12 GND 0.03865f
C3363 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n17 GND 0.11784f
C3364 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n18 GND 0.1843f
C3365 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n19 GND 0.83617f
C3366 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t5 GND 0.03865f
C3367 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t9 GND 0.0619f
C3368 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n20 GND 0.11809f
C3369 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.logic_shift_seg2_0.x7.A GND 0.0153f
C3370 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n21 GND 0.21398f
C3371 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n22 GND 4.36182f
C3372 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n23 GND 8.09385f
C3373 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n24 GND 0.43725f
C3374 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n25 GND 0.03543f
C3375 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t0 GND 0.0374f
C3376 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.t3 GND 0.0374f
C3377 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_7/lvsf_0.IN.n26 GND 0.08213f
C3378 a_35435_18538.t3 GND 0.05539f
C3379 a_35435_18538.t2 GND 0.05331f
C3380 a_35435_18538.n0 GND 0.5884f
C3381 a_35435_18538.t0 GND 0.09815f
C3382 a_35435_18538.n1 GND 1.64869f
C3383 a_35435_18538.t1 GND 0.05605f
C3384 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t24 GND 2.65181f
C3385 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t1 GND 0.10532f
C3386 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t0 GND 0.39669f
C3387 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n0 GND 0.35115f
C3388 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t2 GND 0.39669f
C3389 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n1 GND 0.16403f
C3390 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t3 GND 0.10454f
C3391 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n2 GND 0.19634f
C3392 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n3 GND 0.89301f
C3393 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t5 GND 0.03518f
C3394 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t4 GND 0.04509f
C3395 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n4 GND 0.51038f
C3396 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t15 GND 0.2035f
C3397 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t17 GND 0.20271f
C3398 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n5 GND 0.41896f
C3399 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t28 GND 0.20271f
C3400 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n6 GND 0.17856f
C3401 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t25 GND 0.20271f
C3402 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n7 GND 0.17856f
C3403 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t11 GND 0.20271f
C3404 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n8 GND 0.17856f
C3405 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t8 GND 0.20271f
C3406 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n9 GND 0.17856f
C3407 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t16 GND 0.20271f
C3408 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n10 GND 0.17856f
C3409 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t19 GND 0.20271f
C3410 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n11 GND 0.17856f
C3411 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t22 GND 0.20271f
C3412 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n12 GND 0.17856f
C3413 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t20 GND 0.20271f
C3414 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n13 GND 0.17856f
C3415 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t23 GND 0.20271f
C3416 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n14 GND 0.17856f
C3417 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t27 GND 0.20271f
C3418 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n15 GND 0.17856f
C3419 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t7 GND 0.20271f
C3420 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n16 GND 0.17856f
C3421 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t10 GND 0.20271f
C3422 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n17 GND 0.17856f
C3423 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t13 GND 0.20271f
C3424 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n18 GND 0.17856f
C3425 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t14 GND 0.20271f
C3426 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n19 GND 0.17856f
C3427 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t18 GND 0.20271f
C3428 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n20 GND 0.17856f
C3429 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t21 GND 0.20271f
C3430 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n21 GND 0.17856f
C3431 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t26 GND 0.20271f
C3432 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n22 GND 0.17856f
C3433 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t6 GND 0.20271f
C3434 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n23 GND 0.17856f
C3435 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t9 GND 0.20271f
C3436 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n24 GND 0.17856f
C3437 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.t12 GND 0.20271f
C3438 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n25 GND 0.16737f
C3439 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n26 GND 1.68902f
C3440 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBPLV.n27 GND 2.3067f
C3441 a_21596_17121.t3 GND 0.07113f
C3442 a_21596_17121.t4 GND 0.05948f
C3443 a_21596_17121.n0 GND 2.3636f
C3444 a_21596_17121.t1 GND 0.05948f
C3445 a_21596_17121.n1 GND 1.41357f
C3446 a_21596_17121.t2 GND 0.05948f
C3447 a_21596_17121.n2 GND 1.49069f
C3448 a_21596_17121.t5 GND 0.06059f
C3449 a_21596_17121.n3 GND 1.66289f
C3450 a_21596_17121.t0 GND 0.05908f
C3451 a_32851_7938.t2 GND 0.12718f
C3452 a_32851_7938.t1 GND 0.07284f
C3453 a_32851_7938.n0 GND 6.19294f
C3454 a_32851_7938.t0 GND 0.10705f
C3455 top_segment_4_1.b2.t1 GND 0.088f
C3456 top_segment_4_1.b2.n0 GND 0.03608f
C3457 top_segment_4_1.b2.n1 GND 0.07767f
C3458 top_segment_4_1.b2.n2 GND 0.05156f
C3459 top_segment_4_1.b2.t8 GND 0.17397f
C3460 top_segment_4_1.b2.n3 GND 0.20692f
C3461 top_segment_4_1.b2.t9 GND 0.17397f
C3462 top_segment_4_1.b2.n4 GND 0.27312f
C3463 top_segment_4_1.b2.t4 GND 0.17481f
C3464 top_segment_4_1.b2.n5 GND 0.45411f
C3465 top_segment_4_1.b2.t7 GND 0.17204f
C3466 top_segment_4_1.b2.n6 GND 9.43278f
C3467 top_segment_4_1.b2.t3 GND 0.16643f
C3468 top_segment_4_1.b2.t5 GND 0.16559f
C3469 top_segment_4_1.b2.n7 GND 0.48732f
C3470 top_segment_4_1.b2.t2 GND 0.16643f
C3471 top_segment_4_1.b2.n8 GND 0.41221f
C3472 top_segment_4_1.b2.t6 GND 0.16368f
C3473 top_segment_4_1.b2.n9 GND 1.87395f
C3474 top_segment_4_1.b2.n10 GND 12.201f
C3475 top_segment_4_1.b2.n11 GND 0.05551f
C3476 top_segment_4_1.b2.t0 GND 0.0843f
C3477 top_segment_4_1.b2.n12 GND 0.0436f
C3478 a_13588_5238.t3 GND 0.08408f
C3479 a_13588_5238.t2 GND 0.0646f
C3480 a_13588_5238.n0 GND 3.95828f
C3481 a_13588_5238.t1 GND 0.08235f
C3482 a_13588_5238.t4 GND 0.0646f
C3483 a_13588_5238.n1 GND 4.76416f
C3484 a_13588_5238.n2 GND 3.79219f
C3485 a_13588_5238.t0 GND 0.08975f
C3486 top_segment_4_1.DEC2.t1 GND 0.08474f
C3487 top_segment_4_1.DEC2.n0 GND 0.03475f
C3488 top_segment_4_1.DEC2.n1 GND 0.0748f
C3489 top_segment_4_1.DEC2.n2 GND 0.04966f
C3490 top_segment_4_1.DEC2.t10 GND 0.16835f
C3491 top_segment_4_1.DEC2.t4 GND 0.16754f
C3492 top_segment_4_1.DEC2.n3 GND 0.52525f
C3493 top_segment_4_1.DEC2.t6 GND 0.16754f
C3494 top_segment_4_1.DEC2.n4 GND 0.26303f
C3495 top_segment_4_1.DEC2.t14 GND 0.16754f
C3496 top_segment_4_1.DEC2.n5 GND 0.26303f
C3497 top_segment_4_1.DEC2.t16 GND 0.16754f
C3498 top_segment_4_1.DEC2.n6 GND 0.26303f
C3499 top_segment_4_1.DEC2.t5 GND 0.16754f
C3500 top_segment_4_1.DEC2.n7 GND 0.26303f
C3501 top_segment_4_1.DEC2.t13 GND 0.16754f
C3502 top_segment_4_1.DEC2.n8 GND 0.26303f
C3503 top_segment_4_1.DEC2.t15 GND 0.16568f
C3504 top_segment_4_1.DEC2.t17 GND 0.16835f
C3505 top_segment_4_1.DEC2.t8 GND 0.16835f
C3506 top_segment_4_1.DEC2.t12 GND 0.16754f
C3507 top_segment_4_1.DEC2.n9 GND 0.52525f
C3508 top_segment_4_1.DEC2.t11 GND 0.16754f
C3509 top_segment_4_1.DEC2.n10 GND 0.26303f
C3510 top_segment_4_1.DEC2.t9 GND 0.16754f
C3511 top_segment_4_1.DEC2.n11 GND 0.26303f
C3512 top_segment_4_1.DEC2.t2 GND 0.16754f
C3513 top_segment_4_1.DEC2.n12 GND 0.26303f
C3514 top_segment_4_1.DEC2.t3 GND 0.16754f
C3515 top_segment_4_1.DEC2.n13 GND 0.26303f
C3516 top_segment_4_1.DEC2.n14 GND 0.43732f
C3517 top_segment_4_1.DEC2.t7 GND 0.16568f
C3518 top_segment_4_1.DEC2.n15 GND 0.42527f
C3519 top_segment_4_1.DEC2.n16 GND 0.19515f
C3520 top_segment_4_1.DEC2.n17 GND 15.7048f
C3521 top_segment_4_1.DEC2.n18 GND 0.08218f
C3522 top_segment_4_1.DEC2.t0 GND 0.08119f
C3523 top_segment_4_1.DEC2.n19 GND 0.04199f
C3524 a_31905_7938.t2 GND 0.05347f
C3525 a_31905_7938.t1 GND 0.03963f
C3526 a_31905_7938.n0 GND 2.76188f
C3527 a_31905_7938.t0 GND 0.04502f
C3528 top_segment_4_1.bb2.t1 GND 0.0857f
C3529 top_segment_4_1.bb2.n0 GND 0.03514f
C3530 top_segment_4_1.bb2.n1 GND 0.07564f
C3531 top_segment_4_1.bb2.n2 GND 0.05022f
C3532 top_segment_4_1.bb2.t4 GND 0.17025f
C3533 top_segment_4_1.bb2.t5 GND 0.16944f
C3534 top_segment_4_1.bb2.n3 GND 0.53119f
C3535 top_segment_4_1.bb2.t3 GND 0.16944f
C3536 top_segment_4_1.bb2.n4 GND 0.215f
C3537 top_segment_4_1.bb2.n5 GND 0.17708f
C3538 top_segment_4_1.bb2.t8 GND 0.16755f
C3539 top_segment_4_1.bb2.n6 GND 8.8549f
C3540 top_segment_4_1.bb2.t9 GND 0.16209f
C3541 top_segment_4_1.bb2.t11 GND 0.16128f
C3542 top_segment_4_1.bb2.n7 GND 0.49611f
C3543 top_segment_4_1.bb2.t2 GND 0.16209f
C3544 top_segment_4_1.bb2.n8 GND 0.37997f
C3545 top_segment_4_1.bb2.t7 GND 0.15942f
C3546 top_segment_4_1.bb2.n9 GND 1.79953f
C3547 top_segment_4_1.bb2.n10 GND 11.7595f
C3548 top_segment_4_1.bb2.t10 GND 0.29972f
C3549 top_segment_4_1.bb2.t6 GND 0.16627f
C3550 top_segment_4_1.bb2.n11 GND 0.26118f
C3551 top_segment_4_1.bb2.n12 GND 0.05196f
C3552 top_segment_4_1.bb2.n13 GND 0.0745f
C3553 top_segment_4_1.bb2.n14 GND 0.04247f
C3554 top_segment_4_1.bb2.t0 GND 0.0821f
C3555 top_segment_3_0.bb[4].t1 GND 0.09672f
C3556 top_segment_3_0.bb[4].n0 GND 0.03966f
C3557 top_segment_3_0.bb[4].n1 GND 0.08537f
C3558 top_segment_3_0.bb[4].n2 GND 0.05668f
C3559 top_segment_3_0.bb[4].t2 GND 0.19122f
C3560 top_segment_3_0.bb[4].n3 GND 0.24119f
C3561 top_segment_3_0.bb[4].t4 GND 0.19213f
C3562 top_segment_3_0.bb[4].n4 GND 0.49912f
C3563 top_segment_3_0.bb[4].t6 GND 0.18909f
C3564 top_segment_3_0.bb[4].n5 GND 14.5942f
C3565 top_segment_3_0.bb[4].t3 GND 0.33825f
C3566 top_segment_3_0.bb[4].t5 GND 0.18764f
C3567 top_segment_3_0.bb[4].n6 GND 0.29475f
C3568 top_segment_3_0.bb[4].n7 GND 0.05864f
C3569 top_segment_3_0.bb[4].n8 GND 0.08407f
C3570 top_segment_3_0.bb[4].n9 GND 0.04793f
C3571 top_segment_3_0.bb[4].t0 GND 0.09266f
C3572 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t1 GND 0.04329f
C3573 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t2 GND 0.04329f
C3574 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n0 GND 0.09506f
C3575 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n1 GND 0.04101f
C3576 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t13 GND 0.04474f
C3577 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t6 GND 0.07165f
C3578 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n2 GND 0.13662f
C3579 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n3 GND 0.1482f
C3580 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n4 GND 0.5264f
C3581 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t4 GND 0.07295f
C3582 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t15 GND 0.04581f
C3583 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n5 GND 0.09982f
C3584 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n6 GND 0.12298f
C3585 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t9 GND 0.07295f
C3586 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t5 GND 0.04581f
C3587 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n7 GND 0.11271f
C3588 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n8 GND 0.15523f
C3589 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n9 GND 0.50079f
C3590 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n10 GND 0.64061f
C3591 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t12 GND 0.04476f
C3592 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t16 GND 0.07168f
C3593 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n11 GND 0.13717f
C3594 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n12 GND 0.47666f
C3595 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n13 GND 1.2109f
C3596 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t8 GND 0.07156f
C3597 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t11 GND 0.04466f
C3598 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n14 GND 0.1408f
C3599 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n15 GND 0.1064f
C3600 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n16 GND 0.7135f
C3601 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t7 GND 0.04466f
C3602 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t10 GND 0.07156f
C3603 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n17 GND 0.14228f
C3604 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t14 GND 0.04474f
C3605 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t17 GND 0.07165f
C3606 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n18 GND 0.1364f
C3607 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n19 GND 0.01603f
C3608 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n20 GND 0.16255f
C3609 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n21 GND 12.0678f
C3610 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n22 GND 8.45355f
C3611 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t3 GND 0.02814f
C3612 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].t0 GND 0.02814f
C3613 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n23 GND 0.06709f
C3614 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[8].n24 GND 0.1318f
C3615 top_segment_3_0.bb[6].t0 GND 0.0937f
C3616 top_segment_3_0.bb[6].n0 GND 0.03842f
C3617 top_segment_3_0.bb[6].n1 GND 0.0827f
C3618 top_segment_3_0.bb[6].n2 GND 0.05491f
C3619 top_segment_3_0.bb[6].t1 GND 0.08977f
C3620 top_segment_3_0.bb[6].n3 GND 0.01134f
C3621 top_segment_3_0.bb[6].t6 GND 0.18615f
C3622 top_segment_3_0.bb[6].t11 GND 0.18526f
C3623 top_segment_3_0.bb[6].n4 GND 0.58079f
C3624 top_segment_3_0.bb[6].t5 GND 0.18526f
C3625 top_segment_3_0.bb[6].n5 GND 0.29084f
C3626 top_segment_3_0.bb[6].t10 GND 0.18526f
C3627 top_segment_3_0.bb[6].n6 GND 0.29084f
C3628 top_segment_3_0.bb[6].t12 GND 0.18526f
C3629 top_segment_3_0.bb[6].n7 GND 0.29084f
C3630 top_segment_3_0.bb[6].t8 GND 0.18526f
C3631 top_segment_3_0.bb[6].n8 GND 0.29084f
C3632 top_segment_3_0.bb[6].t2 GND 0.18526f
C3633 top_segment_3_0.bb[6].n9 GND 0.29084f
C3634 top_segment_3_0.bb[6].t4 GND 0.18526f
C3635 top_segment_3_0.bb[6].n10 GND 0.29022f
C3636 top_segment_3_0.bb[6].t9 GND 0.18526f
C3637 top_segment_3_0.bb[6].n11 GND 0.19865f
C3638 top_segment_3_0.bb[6].n12 GND 16.0287f
C3639 top_segment_3_0.bb[6].t3 GND 0.3277f
C3640 top_segment_3_0.bb[6].t7 GND 0.18179f
C3641 top_segment_3_0.bb[6].n13 GND 0.28556f
C3642 top_segment_3_0.bb[6].n14 GND 0.05681f
C3643 top_segment_3_0.bb[6].n15 GND 0.08145f
C3644 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t1 GND 0.04173f
C3645 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.sky130_fd_sc_hd__inv_1_0.Y GND 0.08421f
C3646 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t0 GND 0.06405f
C3647 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.t2 GND 0.14686f
C3648 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.SB[3] GND 2.03364f
C3649 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.SB[3] GND 0.20139f
C3650 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.INB.n0 GND 0.12812f
C3651 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t1 GND 0.06182f
C3652 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t5 GND 0.21263f
C3653 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[3] GND 3.59225f
C3654 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[3] GND 0.2209f
C3655 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t4 GND 0.04704f
C3656 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t3 GND 0.02938f
C3657 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n0 GND 0.08811f
C3658 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n1 GND 0.02491f
C3659 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n2 GND 0.32297f
C3660 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n3 GND 0.16531f
C3661 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x3/x3.Y GND 0.14996f
C3662 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n4 GND 0.02367f
C3663 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t0 GND 0.02839f
C3664 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.t2 GND 0.02839f
C3665 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n5 GND 0.08229f
C3666 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_2/lvsf_0.IN.n6 GND 0.01239f
C3667 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t1 GND 0.0305f
C3668 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t2 GND 0.0305f
C3669 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n0 GND 0.07274f
C3670 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n1 GND 0.1429f
C3671 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t8 GND 0.073f
C3672 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t13 GND 0.04302f
C3673 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t18 GND 0.073f
C3674 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t10 GND 0.04302f
C3675 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n2 GND 0.12249f
C3676 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n3 GND 0.18172f
C3677 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n4 GND 0.0548f
C3678 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t5 GND 0.07759f
C3679 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t9 GND 0.04842f
C3680 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n5 GND 0.15426f
C3681 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t14 GND 0.07769f
C3682 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t17 GND 0.04851f
C3683 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n6 GND 0.14788f
C3684 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n7 GND 0.04318f
C3685 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t15 GND 0.04851f
C3686 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t6 GND 0.07769f
C3687 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n8 GND 0.14809f
C3688 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n9 GND 0.25203f
C3689 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n10 GND 0.72876f
C3690 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t4 GND 0.07749f
C3691 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t16 GND 0.04834f
C3692 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n11 GND 0.1591f
C3693 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n12 GND 1.10696f
C3694 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t12 GND 0.04966f
C3695 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t19 GND 0.07909f
C3696 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n13 GND 0.10732f
C3697 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n14 GND 1.43878f
C3698 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t7 GND 0.04966f
C3699 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t11 GND 0.07909f
C3700 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n15 GND 0.10732f
C3701 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n16 GND 5.7562f
C3702 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n17 GND 11.8589f
C3703 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n18 GND 1.22867f
C3704 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n19 GND 0.03358f
C3705 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n20 GND 0.04446f
C3706 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t3 GND 0.04693f
C3707 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].t0 GND 0.04693f
C3708 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_1.bb[1].n21 GND 0.10307f
C3709 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t2 GND 0.03736f
C3710 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t3 GND 0.03736f
C3711 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n0 GND 0.08204f
C3712 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_7.x1.Y GND 0.18772f
C3713 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n1 GND 0.03539f
C3714 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t6 GND 0.05811f
C3715 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t10 GND 0.03424f
C3716 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t5 GND 0.05811f
C3717 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t9 GND 0.03424f
C3718 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n2 GND 0.0975f
C3719 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n3 GND 0.14465f
C3720 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n4 GND 0.04362f
C3721 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t11 GND 0.06176f
C3722 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t4 GND 0.03854f
C3723 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n5 GND 0.12163f
C3724 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_2.B GND 0.01494f
C3725 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n6 GND 0.05564f
C3726 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t7 GND 0.06176f
C3727 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t8 GND 0.03854f
C3728 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n7 GND 0.12159f
C3729 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.dec_logic_0/sky130_fd_sc_hd__nand2_1_0.B GND 0.01532f
C3730 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n8 GND 0.04107f
C3731 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n9 GND 0.63673f
C3732 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/dec_2_0/decoder_2to4_0.bb[0] GND 2.63598f
C3733 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t12 GND 0.23379f
C3734 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n10 GND 10.3706f
C3735 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n11 GND 2.64516f
C3736 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n12 GND 0.02673f
C3737 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t0 GND 0.02428f
C3738 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.t1 GND 0.02428f
C3739 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n13 GND 0.0579f
C3740 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_5/lvsf_0.INB.n14 GND 0.11375f
C3741 a_32181_7938.t1 GND 0.09175f
C3742 a_32181_7938.t2 GND 0.10894f
C3743 a_32181_7938.n0 GND 5.52296f
C3744 a_32181_7938.t0 GND 0.07635f
C3745 a_26167_5238.t4 GND 0.13813f
C3746 a_26167_5238.t1 GND 0.0814f
C3747 a_26167_5238.n0 GND 5.35733f
C3748 a_26167_5238.t2 GND 0.17912f
C3749 a_26167_5238.n1 GND 4.85263f
C3750 a_26167_5238.t3 GND 0.17054f
C3751 a_26167_5238.n2 GND 5.33946f
C3752 a_26167_5238.t0 GND 0.0814f
C3753 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t0 GND 0.37557f
C3754 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t3 GND 0.19527f
C3755 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t2 GND 0.19937f
C3756 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n0 GND 1.75815f
C3757 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n1 GND 2.71685f
C3758 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.t1 GND 0.19137f
C3759 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S3.n2 GND 0.35177f
C3760 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t4 GND 0.07548f
C3761 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t3 GND 0.07543f
C3762 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n0 GND 0.1418f
C3763 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t1 GND 0.07543f
C3764 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t0 GND 0.28512f
C3765 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t6 GND 0.2877f
C3766 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t7 GND 0.28677f
C3767 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n1 GND 0.35847f
C3768 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t12 GND 0.28766f
C3769 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t8 GND 0.28677f
C3770 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n2 GND 0.35058f
C3771 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n3 GND 0.08769f
C3772 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n4 GND 0.15103f
C3773 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t2 GND 0.28512f
C3774 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t10 GND 0.28766f
C3775 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t11 GND 0.28677f
C3776 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n5 GND 0.35058f
C3777 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t9 GND 0.2877f
C3778 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t13 GND 0.28677f
C3779 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n6 GND 0.35847f
C3780 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n7 GND 0.08769f
C3781 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n8 GND 0.15103f
C3782 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n9 GND 0.1243f
C3783 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n10 GND 0.13769f
C3784 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n11 GND 0.35047f
C3785 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.n12 GND 0.26235f
C3786 top_dcell_routing_0.top_dcell_bias_0/top_bias_lvsf_dec_0.cm2_pcell_0.cm2_pcell2_0.S0.t5 GND 0.07543f
C3787 top_segment_1_0.rseg_1_v3_1.v56.t1 GND 0.03703f
C3788 top_segment_1_0.rseg_1_v3_1.v56.t0 GND 0.12367f
C3789 top_segment_1_0.rseg_1_v3_1.v56.t2 GND 0.36626f
C3790 top_segment_1_0.rseg_1_v3_1.v56.n0 GND 2.56501f
C3791 a_28327_6674.t4 GND 0.04115f
C3792 a_28327_6674.t1 GND 0.05703f
C3793 a_28327_6674.n0 GND 1.94212f
C3794 a_28327_6674.t2 GND 0.03868f
C3795 a_28327_6674.n1 GND 1.52384f
C3796 a_28327_6674.t3 GND 0.06894f
C3797 a_28327_6674.n2 GND 2.78956f
C3798 a_28327_6674.t0 GND 0.03868f
C3799 top_segment_2_0.DEC2[3].t1 GND 0.08361f
C3800 top_segment_2_0.DEC2[3].t0 GND 0.09824f
C3801 top_segment_2_0.DEC2[3].n0 GND 0.50703f
C3802 top_segment_2_0.DEC2[3].t8 GND 0.3905f
C3803 top_segment_2_0.DEC2[3].t6 GND 0.38885f
C3804 top_segment_2_0.DEC2[3].n1 GND 0.65358f
C3805 top_segment_2_0.DEC2[3].t9 GND 0.38885f
C3806 top_segment_2_0.DEC2[3].n2 GND 0.57451f
C3807 top_segment_2_0.DEC2[3].n3 GND 0.88555f
C3808 top_segment_2_0.DEC2[3].t11 GND 0.11913f
C3809 top_segment_2_0.DEC2[3].t22 GND 0.11753f
C3810 top_segment_2_0.DEC2[3].n4 GND 7.35149f
C3811 top_segment_2_0.DEC2[3].t13 GND 0.1195f
C3812 top_segment_2_0.DEC2[3].t10 GND 0.1189f
C3813 top_segment_2_0.DEC2[3].n5 GND 0.38728f
C3814 top_segment_2_0.DEC2[3].t12 GND 0.1189f
C3815 top_segment_2_0.DEC2[3].n6 GND 0.19394f
C3816 top_segment_2_0.DEC2[3].t15 GND 0.1189f
C3817 top_segment_2_0.DEC2[3].n7 GND 0.19394f
C3818 top_segment_2_0.DEC2[3].t18 GND 0.1189f
C3819 top_segment_2_0.DEC2[3].n8 GND 0.19394f
C3820 top_segment_2_0.DEC2[3].t19 GND 0.1189f
C3821 top_segment_2_0.DEC2[3].n9 GND 0.19394f
C3822 top_segment_2_0.DEC2[3].t23 GND 0.1189f
C3823 top_segment_2_0.DEC2[3].n10 GND 0.19394f
C3824 top_segment_2_0.DEC2[3].t2 GND 0.11753f
C3825 top_segment_2_0.DEC2[3].t14 GND 0.1195f
C3826 top_segment_2_0.DEC2[3].t7 GND 0.1199f
C3827 top_segment_2_0.DEC2[3].t20 GND 0.11925f
C3828 top_segment_2_0.DEC2[3].n11 GND 0.41942f
C3829 top_segment_2_0.DEC2[3].t3 GND 0.11925f
C3830 top_segment_2_0.DEC2[3].n12 GND 0.21004f
C3831 top_segment_2_0.DEC2[3].t24 GND 0.11925f
C3832 top_segment_2_0.DEC2[3].n13 GND 0.21004f
C3833 top_segment_2_0.DEC2[3].t21 GND 0.11925f
C3834 top_segment_2_0.DEC2[3].n14 GND 0.21004f
C3835 top_segment_2_0.DEC2[3].t4 GND 0.11925f
C3836 top_segment_2_0.DEC2[3].n15 GND 0.21004f
C3837 top_segment_2_0.DEC2[3].n16 GND 0.32389f
C3838 top_segment_2_0.DEC2[3].t17 GND 0.11753f
C3839 top_segment_2_0.DEC2[3].n17 GND 0.40813f
C3840 top_segment_2_0.DEC2[3].n18 GND 0.3895f
C3841 top_segment_2_0.DEC2[3].n19 GND 0.0959f
C3842 top_segment_2_0.DEC2[3].n20 GND 10.4542f
C3843 top_segment_2_0.DEC2[3].t16 GND 0.22097f
C3844 top_segment_2_0.DEC2[3].t5 GND 0.12258f
C3845 top_segment_2_0.DEC2[3].n21 GND 0.19255f
C3846 top_segment_2_0.DEC2[3].n22 GND 0.03361f
C3847 top_segment_2_0.DEC2[3].n23 GND 0.26303f
C3848 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t0 GND 0.07568f
C3849 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t2 GND 0.01404f
C3850 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t1 GND 0.01404f
C3851 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n0 GND 0.06081f
C3852 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t4 GND 0.02235f
C3853 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t5 GND 0.03579f
C3854 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n1 GND 0.06697f
C3855 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n2 GND 0.01729f
C3856 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.t3 GND 0.1888f
C3857 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.S[4] GND 3.43312f
C3858 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.S[4] GND 0.36483f
C3859 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n3 GND 0.30007f
C3860 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n4 GND 0.10839f
C3861 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.seg_selector_lvsf_0/lvsf_inv_3/lvsf_0.IN.n5 GND 0.04586f
C3862 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.seg_selector_logic_0.x4/x3.Y GND 0.04408f
C3863 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t2 GND 0.04411f
C3864 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t3 GND 0.04411f
C3865 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n0 GND 0.09687f
C3866 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.buffer_bus_0/buffer_cell_5.x2.Y GND 0.22166f
C3867 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n1 GND 0.04179f
C3868 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t4 GND 0.73789f
C3869 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n2 GND 16.6536f
C3870 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t0 GND 0.02867f
C3871 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.t1 GND 0.02867f
C3872 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n3 GND 0.06836f
C3873 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.lvsf_7bit_0/lvsf_buff_2/lvsf_0.IN.n4 GND 0.1343f
C3874 top_segment_2_0.rseg_2_v3_0.v10.t1 GND -0.04356f
C3875 top_segment_2_0.rseg_2_v3_0.v10.n0 GND -0.90533f
C3876 top_segment_2_0.rseg_2_v3_0.v10.t0 GND -0.0437f
C3877 a_19094_19162.t2 GND 0.12781f
C3878 a_19094_19162.t1 GND 0.05892f
C3879 a_19094_19162.n0 GND 4.03512f
C3880 a_19094_19162.t3 GND 0.06702f
C3881 a_19094_19162.n1 GND 5.04796f
C3882 a_19094_19162.t0 GND 0.16318f
C3883 top_segment_2_0.DEC0[0].t16 GND 0.13816f
C3884 top_segment_2_0.DEC0[0].n0 GND 0.17342f
C3885 top_segment_2_0.DEC0[0].t8 GND 0.13816f
C3886 top_segment_2_0.DEC0[0].n1 GND 0.22536f
C3887 top_segment_2_0.DEC0[0].t20 GND 0.13816f
C3888 top_segment_2_0.DEC0[0].n2 GND 0.22536f
C3889 top_segment_2_0.DEC0[0].t15 GND 0.13816f
C3890 top_segment_2_0.DEC0[0].n3 GND 0.22536f
C3891 top_segment_2_0.DEC0[0].t4 GND 0.13816f
C3892 top_segment_2_0.DEC0[0].n4 GND 0.22536f
C3893 top_segment_2_0.DEC0[0].t2 GND 0.13887f
C3894 top_segment_2_0.DEC0[0].t9 GND 0.13816f
C3895 top_segment_2_0.DEC0[0].n5 GND 0.45002f
C3896 top_segment_2_0.DEC0[0].t18 GND 0.13816f
C3897 top_segment_2_0.DEC0[0].n6 GND 0.22536f
C3898 top_segment_2_0.DEC0[0].t3 GND 0.13816f
C3899 top_segment_2_0.DEC0[0].n7 GND 0.22536f
C3900 top_segment_2_0.DEC0[0].t11 GND 0.13816f
C3901 top_segment_2_0.DEC0[0].n8 GND 0.22536f
C3902 top_segment_2_0.DEC0[0].t10 GND 0.13816f
C3903 top_segment_2_0.DEC0[0].n9 GND 0.22536f
C3904 top_segment_2_0.DEC0[0].t13 GND 0.13816f
C3905 top_segment_2_0.DEC0[0].n10 GND 0.22536f
C3906 top_segment_2_0.DEC0[0].t5 GND 0.13816f
C3907 top_segment_2_0.DEC0[0].n11 GND 0.22536f
C3908 top_segment_2_0.DEC0[0].t12 GND 0.13816f
C3909 top_segment_2_0.DEC0[0].n12 GND 0.22536f
C3910 top_segment_2_0.DEC0[0].t19 GND 0.13816f
C3911 top_segment_2_0.DEC0[0].n13 GND 0.22536f
C3912 top_segment_2_0.DEC0[0].t7 GND 0.13816f
C3913 top_segment_2_0.DEC0[0].n14 GND 0.22536f
C3914 top_segment_2_0.DEC0[0].n15 GND 0.1517f
C3915 top_segment_2_0.DEC0[0].t17 GND 0.13657f
C3916 top_segment_2_0.DEC0[0].n16 GND 15.1085f
C3917 top_segment_2_0.DEC0[0].t0 GND 0.11443f
C3918 top_segment_2_0.DEC0[0].t1 GND 0.09714f
C3919 top_segment_2_0.DEC0[0].n17 GND 0.94738f
C3920 top_segment_2_0.DEC0[0].t14 GND 0.45357f
C3921 top_segment_2_0.DEC0[0].t21 GND 0.4517f
C3922 top_segment_2_0.DEC0[0].n18 GND 0.74878f
C3923 top_segment_2_0.DEC0[0].t6 GND 0.4517f
C3924 top_segment_2_0.DEC0[0].n19 GND 0.38634f
C3925 top_segment_2_0.DEC0[0].n20 GND 0.7067f
C3926 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t1 GND 0.01248f
C3927 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t2 GND 0.09426f
C3928 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.t0 GND 0.09768f
C3929 top_segment_4_1.rseg_4_routing_0/rseg_4_v3_0.v53.n0 GND 1.54809f
C3930 top_segment_1_0.rseg_1_v3_1.v9.t1 GND 0.04754f
C3931 top_segment_1_0.rseg_1_v3_1.v9.t2 GND 0.14298f
C3932 top_segment_1_0.rseg_1_v3_1.v9.t0 GND 0.14263f
C3933 top_segment_1_0.rseg_1_v3_1.v9.n0 GND 2.55569f
C3934 a_28603_6674.t1 GND 0.0855f
C3935 a_28603_6674.t2 GND 0.10458f
C3936 a_28603_6674.n0 GND 3.75935f
C3937 a_28603_6674.t3 GND 0.07805f
C3938 a_28603_6674.n1 GND 2.99489f
C3939 a_28603_6674.t4 GND 0.14007f
C3940 a_28603_6674.n2 GND 5.65951f
C3941 a_28603_6674.t0 GND 0.07805f
C3942 top_segment_2_0.DEC2[0].t1 GND 0.09748f
C3943 top_segment_2_0.DEC2[0].t0 GND 0.08275f
C3944 top_segment_2_0.DEC2[0].n0 GND 0.80704f
C3945 top_segment_2_0.DEC2[0].t15 GND 0.38639f
C3946 top_segment_2_0.DEC2[0].t7 GND 0.38479f
C3947 top_segment_2_0.DEC2[0].n1 GND 0.63787f
C3948 top_segment_2_0.DEC2[0].t20 GND 0.38479f
C3949 top_segment_2_0.DEC2[0].n2 GND 0.32912f
C3950 top_segment_2_0.DEC2[0].n3 GND 0.60202f
C3951 top_segment_2_0.DEC2[0].t18 GND 0.11796f
C3952 top_segment_2_0.DEC2[0].t6 GND 0.11634f
C3953 top_segment_2_0.DEC2[0].n4 GND 3.73702f
C3954 top_segment_2_0.DEC2[0].t21 GND 0.1183f
C3955 top_segment_2_0.DEC2[0].t14 GND 0.1177f
C3956 top_segment_2_0.DEC2[0].n5 GND 0.38336f
C3957 top_segment_2_0.DEC2[0].t19 GND 0.1177f
C3958 top_segment_2_0.DEC2[0].n6 GND 0.19198f
C3959 top_segment_2_0.DEC2[0].t9 GND 0.1177f
C3960 top_segment_2_0.DEC2[0].n7 GND 0.1585f
C3961 top_segment_2_0.DEC2[0].t23 GND 0.1183f
C3962 top_segment_2_0.DEC2[0].t8 GND 0.1177f
C3963 top_segment_2_0.DEC2[0].n8 GND 0.38336f
C3964 top_segment_2_0.DEC2[0].t4 GND 0.1177f
C3965 top_segment_2_0.DEC2[0].n9 GND 0.19198f
C3966 top_segment_2_0.DEC2[0].t24 GND 0.1177f
C3967 top_segment_2_0.DEC2[0].n10 GND 0.1585f
C3968 top_segment_2_0.DEC2[0].n11 GND 0.20637f
C3969 top_segment_2_0.DEC2[0].t10 GND 0.1183f
C3970 top_segment_2_0.DEC2[0].t17 GND 0.1177f
C3971 top_segment_2_0.DEC2[0].n12 GND 0.38336f
C3972 top_segment_2_0.DEC2[0].t13 GND 0.1177f
C3973 top_segment_2_0.DEC2[0].n13 GND 0.19198f
C3974 top_segment_2_0.DEC2[0].t16 GND 0.1177f
C3975 top_segment_2_0.DEC2[0].n14 GND 0.19198f
C3976 top_segment_2_0.DEC2[0].t22 GND 0.1177f
C3977 top_segment_2_0.DEC2[0].n15 GND 0.19198f
C3978 top_segment_2_0.DEC2[0].t12 GND 0.1177f
C3979 top_segment_2_0.DEC2[0].n16 GND 0.19198f
C3980 top_segment_2_0.DEC2[0].t2 GND 0.1177f
C3981 top_segment_2_0.DEC2[0].n17 GND 0.19198f
C3982 top_segment_2_0.DEC2[0].t5 GND 0.1177f
C3983 top_segment_2_0.DEC2[0].n18 GND 0.15678f
C3984 top_segment_2_0.DEC2[0].n19 GND 3.06972f
C3985 top_segment_2_0.DEC2[0].n20 GND 10.845f
C3986 top_segment_2_0.DEC2[0].t11 GND 0.21873f
C3987 top_segment_2_0.DEC2[0].t3 GND 0.12134f
C3988 top_segment_2_0.DEC2[0].n21 GND 0.1906f
C3989 top_segment_2_0.DEC2[0].n22 GND 0.03327f
C3990 top_segment_2_0.DEC2[0].n23 GND 0.26302f
C3991 top_segment_2_0.rseg_2_v3_0.v5.t2 GND 0.0447f
C3992 top_segment_2_0.rseg_2_v3_0.v5.t1 GND 0.19887f
C3993 top_segment_2_0.rseg_2_v3_0.v5.n0 GND 4.85619f
C3994 top_segment_2_0.rseg_2_v3_0.v5.t0 GND 0.20023f
C3995 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t2 GND 0.02605f
C3996 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t3 GND 0.02605f
C3997 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n0 GND 0.06212f
C3998 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n1 GND 0.12205f
C3999 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t5 GND 0.06645f
C4000 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t16 GND 0.04151f
C4001 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n2 GND 0.12322f
C4002 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t13 GND 0.06618f
C4003 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t8 GND 0.04129f
C4004 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n3 GND 0.13445f
C4005 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n4 GND 0.15582f
C4006 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t4 GND 0.04136f
C4007 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t9 GND 0.06626f
C4008 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n5 GND 0.13065f
C4009 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n6 GND 0.08905f
C4010 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n7 GND 0.49955f
C4011 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n8 GND 0.84298f
C4012 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t10 GND 0.04136f
C4013 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t17 GND 0.06626f
C4014 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n9 GND 0.13038f
C4015 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n10 GND 0.08233f
C4016 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n11 GND 0.58676f
C4017 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t12 GND 0.06626f
C4018 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t15 GND 0.04136f
C4019 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n12 GND 0.13038f
C4020 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n13 GND 0.05851f
C4021 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t11 GND 0.06626f
C4022 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t14 GND 0.04136f
C4023 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n14 GND 0.13175f
C4024 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t6 GND 0.06635f
C4025 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t7 GND 0.04143f
C4026 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n15 GND 0.1263f
C4027 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n16 GND 0.0229f
C4028 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n17 GND 0.03311f
C4029 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n18 GND 0.46233f
C4030 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n19 GND 11.365f
C4031 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n20 GND 7.93634f
C4032 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n21 GND 0.03797f
C4033 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t0 GND 0.04008f
C4034 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].t1 GND 0.04008f
C4035 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.dcell_lv_0.b[9].n22 GND 0.08803f
C4036 top_segment_2_0.DEC2[2].t24 GND 0.39716f
C4037 top_segment_2_0.DEC2[2].t1 GND 0.10204f
C4038 top_segment_2_0.DEC2[2].t0 GND 0.08684f
C4039 top_segment_2_0.DEC2[2].n0 GND 0.56182f
C4040 top_segment_2_0.DEC2[2].n1 GND 0.44723f
C4041 top_segment_2_0.DEC2[2].t2 GND 0.40559f
C4042 top_segment_2_0.DEC2[2].t15 GND 0.40388f
C4043 top_segment_2_0.DEC2[2].n2 GND 0.89787f
C4044 top_segment_2_0.DEC2[2].n3 GND 0.66766f
C4045 top_segment_2_0.DEC2[2].t3 GND 0.12415f
C4046 top_segment_2_0.DEC2[2].t9 GND 0.12207f
C4047 top_segment_2_0.DEC2[2].n4 GND 6.72012f
C4048 top_segment_2_0.DEC2[2].t22 GND 0.12412f
C4049 top_segment_2_0.DEC2[2].t13 GND 0.1235f
C4050 top_segment_2_0.DEC2[2].n5 GND 0.40225f
C4051 top_segment_2_0.DEC2[2].t18 GND 0.1235f
C4052 top_segment_2_0.DEC2[2].n6 GND 0.20144f
C4053 top_segment_2_0.DEC2[2].t21 GND 0.1235f
C4054 top_segment_2_0.DEC2[2].n7 GND 0.20144f
C4055 top_segment_2_0.DEC2[2].t11 GND 0.1235f
C4056 top_segment_2_0.DEC2[2].n8 GND 0.20144f
C4057 top_segment_2_0.DEC2[2].t5 GND 0.1235f
C4058 top_segment_2_0.DEC2[2].n9 GND 0.20144f
C4059 top_segment_2_0.DEC2[2].t20 GND 0.1235f
C4060 top_segment_2_0.DEC2[2].n10 GND 0.20144f
C4061 top_segment_2_0.DEC2[2].t7 GND 0.12207f
C4062 top_segment_2_0.DEC2[2].t8 GND 0.12412f
C4063 top_segment_2_0.DEC2[2].t6 GND 0.12454f
C4064 top_segment_2_0.DEC2[2].t17 GND 0.12386f
C4065 top_segment_2_0.DEC2[2].n11 GND 0.43564f
C4066 top_segment_2_0.DEC2[2].t4 GND 0.12386f
C4067 top_segment_2_0.DEC2[2].n12 GND 0.21816f
C4068 top_segment_2_0.DEC2[2].t23 GND 0.12386f
C4069 top_segment_2_0.DEC2[2].n13 GND 0.21816f
C4070 top_segment_2_0.DEC2[2].t19 GND 0.12386f
C4071 top_segment_2_0.DEC2[2].n14 GND 0.21816f
C4072 top_segment_2_0.DEC2[2].t14 GND 0.12386f
C4073 top_segment_2_0.DEC2[2].n15 GND 0.21816f
C4074 top_segment_2_0.DEC2[2].n16 GND 0.33641f
C4075 top_segment_2_0.DEC2[2].t10 GND 0.12207f
C4076 top_segment_2_0.DEC2[2].n17 GND 0.42016f
C4077 top_segment_2_0.DEC2[2].n18 GND 0.4247f
C4078 top_segment_2_0.DEC2[2].n19 GND 0.09752f
C4079 top_segment_2_0.DEC2[2].n20 GND 11.1617f
C4080 top_segment_2_0.DEC2[2].t12 GND 0.22951f
C4081 top_segment_2_0.DEC2[2].t16 GND 0.12732f
C4082 top_segment_2_0.DEC2[2].n21 GND 0.19999f
C4083 top_segment_2_0.DEC2[2].n22 GND 0.03491f
C4084 top_segment_2_0.DEC2[2].n23 GND 0.27706f
C4085 top_segment_2_0.rseg_2_v3_0.v41.t2 GND 0.20596f
C4086 top_segment_2_0.rseg_2_v3_0.v41.t1 GND 0.22743f
C4087 top_segment_2_0.rseg_2_v3_0.v41.n0 GND 4.83206f
C4088 top_segment_2_0.rseg_2_v3_0.v41.t0 GND 0.03454f
C4089 top_segment_2_0.rseg_2_v3_0.v42.t1 GND 0.09067f
C4090 top_segment_2_0.rseg_2_v3_0.v42.t2 GND 0.10022f
C4091 top_segment_2_0.rseg_2_v3_0.v42.n0 GND 2.09413f
C4092 top_segment_2_0.rseg_2_v3_0.v42.t0 GND 0.01498f
C4093 a_18769_7938.t2 GND 0.08054f
C4094 a_18769_7938.t1 GND 0.08241f
C4095 a_18769_7938.n0 GND 5.87337f
C4096 a_18769_7938.t0 GND 0.06369f
C4097 a_15714_6674.t3 GND 0.08487f
C4098 a_15714_6674.t4 GND 0.07389f
C4099 a_15714_6674.n0 GND 4.0948f
C4100 a_15714_6674.t2 GND 0.07249f
C4101 a_15714_6674.n1 GND 2.60041f
C4102 a_15714_6674.t1 GND 0.07249f
C4103 a_15714_6674.n2 GND 5.60801f
C4104 a_15714_6674.t0 GND 0.09304f
C4105 top_segment_4_1.bb3.t1 GND 0.07082f
C4106 top_segment_4_1.bb3.n0 GND 0.02904f
C4107 top_segment_4_1.bb3.n1 GND 0.06251f
C4108 top_segment_4_1.bb3.n2 GND 0.0415f
C4109 top_segment_4_1.bb3.t11 GND 0.1407f
C4110 top_segment_4_1.bb3.n3 GND 0.32652f
C4111 top_segment_4_1.bb3.t20 GND 0.13847f
C4112 top_segment_4_1.bb3.n4 GND 3.60149f
C4113 top_segment_4_1.bb3.t17 GND 0.1407f
C4114 top_segment_4_1.bb3.t2 GND 0.14002f
C4115 top_segment_4_1.bb3.n5 GND 0.43898f
C4116 top_segment_4_1.bb3.t6 GND 0.14002f
C4117 top_segment_4_1.bb3.n6 GND 0.21982f
C4118 top_segment_4_1.bb3.t10 GND 0.14002f
C4119 top_segment_4_1.bb3.n7 GND 0.179f
C4120 top_segment_4_1.bb3.t12 GND 0.14002f
C4121 top_segment_4_1.bb3.n8 GND 0.21982f
C4122 top_segment_4_1.bb3.t5 GND 0.14002f
C4123 top_segment_4_1.bb3.n9 GND 0.21982f
C4124 top_segment_4_1.bb3.t21 GND 0.14002f
C4125 top_segment_4_1.bb3.n10 GND 0.21982f
C4126 top_segment_4_1.bb3.n11 GND 0.14634f
C4127 top_segment_4_1.bb3.t7 GND 0.13847f
C4128 top_segment_4_1.bb3.n12 GND 1.91133f
C4129 top_segment_4_1.bb3.n13 GND 7.65499f
C4130 top_segment_4_1.bb3.t9 GND 0.13396f
C4131 top_segment_4_1.bb3.t16 GND 0.13328f
C4132 top_segment_4_1.bb3.n14 GND 0.43411f
C4133 top_segment_4_1.bb3.t19 GND 0.13328f
C4134 top_segment_4_1.bb3.n15 GND 0.15775f
C4135 top_segment_4_1.bb3.t8 GND 0.13328f
C4136 top_segment_4_1.bb3.n16 GND 0.20387f
C4137 top_segment_4_1.bb3.t15 GND 0.13328f
C4138 top_segment_4_1.bb3.n17 GND 0.21739f
C4139 top_segment_4_1.bb3.t18 GND 0.13328f
C4140 top_segment_4_1.bb3.n18 GND 0.21739f
C4141 top_segment_4_1.bb3.t14 GND 0.13396f
C4142 top_segment_4_1.bb3.n19 GND 0.36306f
C4143 top_segment_4_1.bb3.t3 GND 0.13174f
C4144 top_segment_4_1.bb3.n20 GND 1.9148f
C4145 top_segment_4_1.bb3.n21 GND 7.47526f
C4146 top_segment_4_1.bb3.t4 GND 0.24769f
C4147 top_segment_4_1.bb3.t13 GND 0.1374f
C4148 top_segment_4_1.bb3.n22 GND 0.21584f
C4149 top_segment_4_1.bb3.n23 GND 0.04294f
C4150 top_segment_4_1.bb3.n24 GND 0.06157f
C4151 top_segment_4_1.bb3.n25 GND 0.0351f
C4152 top_segment_4_1.bb3.t0 GND 0.06785f
C4153 VDDH.n0 GND 0.01561f
C4154 VDDH.n1 GND 0.03219f
C4155 VDDH.t258 GND 0.03662f
C4156 VDDH.n2 GND 0.04259f
C4157 VDDH.n3 GND 0.0882f
C4158 VDDH.n4 GND 0.02471f
C4159 VDDH.n5 GND 0.21919f
C4160 VDDH.n6 GND 0.02123f
C4161 VDDH.n7 GND 0.05927f
C4162 VDDH.n8 GND 0.03219f
C4163 VDDH.t245 GND 0.03662f
C4164 VDDH.n9 GND 0.04259f
C4165 VDDH.n10 GND 0.01562f
C4166 VDDH.n11 GND 0.03006f
C4167 VDDH.n12 GND 0.01153f
C4168 VDDH.n13 GND 0.01999f
C4169 VDDH.n14 GND 0.03738f
C4170 VDDH.n15 GND 0.23532f
C4171 VDDH.n17 GND 0.31189f
C4172 VDDH.n18 GND 0.09419f
C4173 VDDH.n19 GND 0.01627f
C4174 VDDH.n20 GND 0.05347f
C4175 VDDH.n22 GND 0.0562f
C4176 VDDH.n23 GND 0.03219f
C4177 VDDH.t241 GND 0.03662f
C4178 VDDH.n24 GND 0.01846f
C4179 VDDH.n25 GND 0.03219f
C4180 VDDH.t252 GND 0.03662f
C4181 VDDH.n26 GND 0.04563f
C4182 VDDH.n27 GND 0.04857f
C4183 VDDH.n28 GND 0.03754f
C4184 VDDH.n29 GND 0.08984f
C4185 VDDH.n30 GND 0.05371f
C4186 VDDH.n31 GND 0.09494f
C4187 VDDH.t184 GND 0.55363f
C4188 VDDH.t7 GND 0.14037f
C4189 VDDH.t40 GND 0.4098f
C4190 VDDH.t74 GND 0.69582f
C4191 VDDH.t28 GND 0.23466f
C4192 VDDH.n32 GND 0.17373f
C4193 VDDH.n33 GND 0.04266f
C4194 VDDH.n34 GND 0.02417f
C4195 VDDH.n35 GND 0.03362f
C4196 VDDH.n36 GND 0.02892f
C4197 VDDH.n38 GND 0.01083f
C4198 VDDH.t8 GND 0.14037f
C4199 VDDH.t76 GND 0.18136f
C4200 VDDH.n42 GND 0.12441f
C4201 VDDH.t5 GND 0.23686f
C4202 VDDH.n50 GND 0.01083f
C4203 VDDH.n53 GND 0.01066f
C4204 VDDH.n55 GND 0.02091f
C4205 VDDH.n61 GND 0.01129f
C4206 VDDH.n62 GND 0.04266f
C4207 VDDH.n63 GND 0.02417f
C4208 VDDH.n66 GND 0.02091f
C4209 VDDH.n69 GND 0.01083f
C4210 VDDH.n71 GND 0.01083f
C4211 VDDH.n73 GND 0.17589f
C4212 VDDH.n81 GND 0.03048f
C4213 VDDH.n82 GND 0.03048f
C4214 VDDH.n83 GND 0.02444f
C4215 VDDH.t211 GND 0.0237f
C4216 VDDH.t45 GND 0.09137f
C4217 VDDH.n88 GND 0.04469f
C4218 VDDH.n92 GND 0.03063f
C4219 VDDH.n94 GND 0.02091f
C4220 VDDH.n95 GND 0.05247f
C4221 VDDH.t83 GND 0.0237f
C4222 VDDH.n100 GND 0.02691f
C4223 VDDH.n101 GND 0.0237f
C4224 VDDH.t171 GND 0.02296f
C4225 VDDH.n102 GND 0.02691f
C4226 VDDH.n108 GND 0.02091f
C4227 VDDH.n113 GND 0.04493f
C4228 VDDH.t164 GND 0.07343f
C4229 VDDH.t29 GND 0.07321f
C4230 VDDH.n114 GND 0.04469f
C4231 VDDH.t62 GND 0.0237f
C4232 VDDH.t270 GND 0.0237f
C4233 VDDH.n116 GND 0.02691f
C4234 VDDH.t152 GND 0.02296f
C4235 VDDH.t278 GND 0.0237f
C4236 VDDH.n126 GND 0.02091f
C4237 VDDH.t233 GND 0.0237f
C4238 VDDH.n137 GND 0.02691f
C4239 VDDH.n138 GND 0.0237f
C4240 VDDH.n139 GND 0.02691f
C4241 VDDH.t162 GND 0.02296f
C4242 VDDH.n140 GND 0.02444f
C4243 VDDH.t100 GND 0.0237f
C4244 VDDH.n144 GND 0.02091f
C4245 VDDH.n148 GND 0.03048f
C4246 VDDH.t87 GND 0.0237f
C4247 VDDH.n150 GND 0.02691f
C4248 VDDH.t85 GND 0.02296f
C4249 VDDH.n156 GND 0.0225f
C4250 VDDH.n157 GND 0.17589f
C4251 VDDH.n158 GND 0.17589f
C4252 VDDH.n166 GND 0.03048f
C4253 VDDH.n167 GND 0.02444f
C4254 VDDH.t268 GND 0.0237f
C4255 VDDH.n172 GND 0.02444f
C4256 VDDH.n175 GND 0.04493f
C4257 VDDH.t27 GND 0.07343f
C4258 VDDH.t2 GND 0.07321f
C4259 VDDH.n176 GND 0.04469f
C4260 VDDH.n181 GND 0.03063f
C4261 VDDH.n183 GND 0.02091f
C4262 VDDH.t173 GND 0.0237f
C4263 VDDH.n189 GND 0.02691f
C4264 VDDH.n190 GND 0.0237f
C4265 VDDH.t167 GND 0.02296f
C4266 VDDH.n191 GND 0.02691f
C4267 VDDH.n197 GND 0.02091f
C4268 VDDH.n202 GND 0.04493f
C4269 VDDH.t305 GND 0.07343f
C4270 VDDH.t207 GND 0.07321f
C4271 VDDH.n203 GND 0.04469f
C4272 VDDH.t38 GND 0.0237f
C4273 VDDH.t286 GND 0.0237f
C4274 VDDH.n205 GND 0.02691f
C4275 VDDH.t146 GND 0.02296f
C4276 VDDH.t49 GND 0.0237f
C4277 VDDH.n215 GND 0.02091f
C4278 VDDH.t231 GND 0.0237f
C4279 VDDH.n226 GND 0.02691f
C4280 VDDH.n227 GND 0.0237f
C4281 VDDH.n228 GND 0.02691f
C4282 VDDH.t235 GND 0.02296f
C4283 VDDH.n229 GND 0.02444f
C4284 VDDH.t0 GND 0.06847f
C4285 VDDH.n230 GND 0.0237f
C4286 VDDH.t158 GND 0.04465f
C4287 VDDH.n231 GND 0.03048f
C4288 VDDH.n233 GND 0.03163f
C4289 VDDH.n241 GND 0.03163f
C4290 VDDH.n243 GND 0.02091f
C4291 VDDH.n245 GND 0.17589f
C4292 VDDH.n247 GND 0.03612f
C4293 VDDH.t272 GND 0.06847f
C4294 VDDH.n257 GND 0.02091f
C4295 VDDH.n259 GND 0.03612f
C4296 VDDH.n263 GND 0.0237f
C4297 VDDH.t240 GND 0.07565f
C4298 VDDH.t122 GND 0.07565f
C4299 VDDH.t169 GND 0.04465f
C4300 VDDH.n264 GND 0.03029f
C4301 VDDH.t81 GND 0.04465f
C4302 VDDH.t197 GND 0.07565f
C4303 VDDH.t187 GND 0.07565f
C4304 VDDH.t150 GND 0.04465f
C4305 VDDH.t288 GND 0.04465f
C4306 VDDH.n266 GND 0.03612f
C4307 VDDH.t186 GND 0.07565f
C4308 VDDH.t92 GND 0.07565f
C4309 VDDH.t160 GND 0.04465f
C4310 VDDH.t303 GND 0.09367f
C4311 VDDH.t156 GND 0.04465f
C4312 VDDH.t65 GND 0.06847f
C4313 VDDH.n270 GND 0.02091f
C4314 VDDH.n272 GND 1.08268f
C4315 VDDH.n273 GND 0.03908f
C4316 VDDH.n274 GND 0.03908f
C4317 VDDH.n275 GND 0.03347f
C4318 VDDH.n276 GND 0.01657f
C4319 VDDH.n277 GND 0.05788f
C4320 VDDH.n278 GND 0.04399f
C4321 VDDH.t242 GND 0.48674f
C4322 VDDH.t21 GND 0.57101f
C4323 VDDH.n279 GND 0.29614f
C4324 VDDH.t12 GND 0.3174f
C4325 VDDH.t24 GND 0.33169f
C4326 VDDH.n280 GND 0.0313f
C4327 VDDH.n281 GND 0.0371f
C4328 VDDH.n283 GND 0.01785f
C4329 VDDH.n284 GND 0.0389f
C4330 VDDH.n285 GND 0.03474f
C4331 VDDH.n286 GND 0.03441f
C4332 VDDH.n287 GND 0.03219f
C4333 VDDH.t264 GND 0.03662f
C4334 VDDH.n288 GND 0.04259f
C4335 VDDH.n289 GND 0.02343f
C4336 VDDH.t255 GND 0.03662f
C4337 VDDH.n290 GND 0.05303f
C4338 VDDH.n291 GND 0.03332f
C4339 VDDH.n292 GND 0.03908f
C4340 VDDH.n293 GND 0.03032f
C4341 VDDH.n294 GND 0.01174f
C4342 VDDH.n295 GND 0.01123f
C4343 VDDH.n296 GND 0.01228f
C4344 VDDH.n297 GND 0.04104f
C4345 VDDH.n298 GND 0.29614f
C4346 VDDH.t16 GND 0.55526f
C4347 VDDH.t14 GND 0.59228f
C4348 VDDH.t249 GND 0.48674f
C4349 VDDH.n299 GND 0.33745f
C4350 VDDH.n300 GND 0.0371f
C4351 VDDH.n302 GND 0.02828f
C4352 VDDH.t248 GND 0.03662f
C4353 VDDH.n303 GND 0.01657f
C4354 VDDH.n304 GND 0.02402f
C4355 VDDH.n305 GND 0.09853f
C4356 VDDH.n306 GND 0.01431f
C4357 VDDH.n307 GND 0.03008f
C4358 VDDH.n308 GND 0.04074f
C4359 VDDH.t33 GND 0.08378f
C4360 VDDH.t306 GND 0.08168f
C4361 VDDH.t36 GND 0.08378f
C4362 VDDH.t177 GND 0.08378f
C4363 VDDH.t307 GND 0.08378f
C4364 VDDH.n310 GND 0.09853f
C4365 VDDH.n312 GND 0.02399f
C4366 VDDH.n313 GND 0.02223f
C4367 VDDH.t217 GND 0.08168f
C4368 VDDH.t213 GND 0.08378f
C4369 VDDH.t210 GND 0.08378f
C4370 VDDH.t216 GND 0.08378f
C4371 VDDH.t35 GND 0.08378f
C4372 VDDH.t179 GND 0.08378f
C4373 VDDH.t34 GND 0.07422f
C4374 VDDH.n314 GND 0.06466f
C4375 VDDH.t215 GND 0.07422f
C4376 VDDH.t219 GND 0.08378f
C4377 VDDH.t214 GND 0.08378f
C4378 VDDH.t218 GND 0.08378f
C4379 VDDH.n315 GND 0.01947f
C4380 VDDH.n316 GND 0.02692f
C4381 VDDH.n317 GND 0.10378f
C4382 VDDH.n318 GND 0.03536f
C4383 VDDH.t90 GND 0.08168f
C4384 VDDH.t284 GND 0.08803f
C4385 VDDH.t176 GND 0.08803f
C4386 VDDH.t237 GND 0.08803f
C4387 VDDH.t277 GND 0.06496f
C4388 VDDH.t281 GND 0.06481f
C4389 VDDH.n319 GND 0.03534f
C4390 VDDH.n321 GND 0.01462f
C4391 VDDH.n322 GND 0.02476f
C4392 VDDH.t280 GND 0.08803f
C4393 VDDH.t56 GND 0.08803f
C4394 VDDH.t58 GND 0.08378f
C4395 VDDH.t57 GND 0.07422f
C4396 VDDH.n324 GND 0.06466f
C4397 VDDH.t55 GND 0.07422f
C4398 VDDH.t52 GND 0.08378f
C4399 VDDH.t51 GND 0.08378f
C4400 VDDH.n325 GND 0.02476f
C4401 VDDH.n327 GND 0.08243f
C4402 VDDH.t53 GND 0.07422f
C4403 VDDH.n329 GND 0.06466f
C4404 VDDH.t141 GND 0.07422f
C4405 VDDH.t64 GND 0.08378f
C4406 VDDH.t60 GND 0.08168f
C4407 VDDH.t61 GND 0.08378f
C4408 VDDH.n330 GND 0.0138f
C4409 VDDH.n331 GND 0.01467f
C4410 VDDH.n332 GND 0.02492f
C4411 VDDH.t59 GND 0.08378f
C4412 VDDH.n333 GND 0.02492f
C4413 VDDH.n335 GND 0.01462f
C4414 VDDH.n336 GND 0.01299f
C4415 VDDH.n337 GND 0.02215f
C4416 VDDH.t54 GND 0.08378f
C4417 VDDH.n338 GND 0.02215f
C4418 VDDH.n339 GND 0.01299f
C4419 VDDH.n340 GND 0.02082f
C4420 VDDH.n341 GND 0.02707f
C4421 VDDH.n342 GND 0.04605f
C4422 VDDH.n343 GND 0.02307f
C4423 VDDH.n344 GND 0.01897f
C4424 VDDH.n345 GND 0.04605f
C4425 VDDH.n346 GND 0.02236f
C4426 VDDH.n347 GND 0.02053f
C4427 VDDH.n349 GND 0.01919f
C4428 VDDH.n350 GND 0.02236f
C4429 VDDH.n351 GND 0.04084f
C4430 VDDH.t220 GND 0.08378f
C4431 VDDH.n352 GND 0.04084f
C4432 VDDH.n353 GND 0.04074f
C4433 VDDH.n354 GND 0.04084f
C4434 VDDH.t178 GND 0.08378f
C4435 VDDH.n355 GND 0.04084f
C4436 VDDH.n356 GND 0.02236f
C4437 VDDH.n357 GND 0.01919f
C4438 VDDH.n358 GND 1.85667f
C4439 VDDH.n359 GND 9.8115f
C4440 VDDH.n360 GND 0.06363f
C4441 VDDH.n361 GND 0.03089f
C4442 VDDH.n362 GND 0.02085f
C4443 VDDH.n363 GND 0.01657f
C4444 VDDH.n364 GND 0.03267f
C4445 VDDH.n365 GND 0.01174f
C4446 VDDH.n366 GND 0.03134f
C4447 VDDH.n367 GND 0.03756f
C4448 VDDH.n368 GND 0.03383f
C4449 VDDH.t261 GND 0.03662f
C4450 VDDH.n369 GND 0.01884f
C4451 VDDH.n370 GND 0.02403f
C4452 VDDH.n371 GND 0.0641f
C4453 VDDH.n372 GND 0.1005f
C4454 VDDH.n373 GND 0.08296f
C4455 VDDH.n374 GND 0.07253f
C4456 VDDH.n375 GND 0.1213f
C4457 VDDH.n376 GND 5.9128f
C4458 VDDH.n377 GND 0.01503f
C4459 VDDH.n378 GND 0.09451f
C4460 VDDH.n379 GND 0.01778f
C4461 VDDH.n380 GND 0.01499f
C4462 VDDH.n381 GND 0.01351f
C4463 VDDH.n382 GND 0.02579f
C4464 VDDH.n383 GND 0.09451f
C4465 VDDH.n384 GND 0.09451f
C4466 VDDH.t107 GND 0.08168f
C4467 VDDH.t105 GND 0.08378f
C4468 VDDH.t106 GND 0.08378f
C4469 VDDH.t121 GND 0.06284f
C4470 VDDH.t109 GND 0.08168f
C4471 VDDH.t120 GND 0.08378f
C4472 VDDH.t118 GND 0.08378f
C4473 VDDH.t110 GND 0.06284f
C4474 VDDH.n386 GND 0.01943f
C4475 VDDH.n387 GND 0.01248f
C4476 VDDH.n388 GND 0.09451f
C4477 VDDH.n389 GND 0.09451f
C4478 VDDH.t203 GND 0.08168f
C4479 VDDH.t126 GND 0.08378f
C4480 VDDH.t297 GND 0.08378f
C4481 VDDH.t299 GND 0.06284f
C4482 VDDH.n391 GND 0.02639f
C4483 VDDH.n392 GND 0.01473f
C4484 VDDH.n393 GND 0.01775f
C4485 VDDH.n394 GND 0.09451f
C4486 VDDH.n395 GND 0.09451f
C4487 VDDH.t123 GND 0.08168f
C4488 VDDH.t125 GND 0.08378f
C4489 VDDH.t300 GND 0.08378f
C4490 VDDH.t200 GND 0.06284f
C4491 VDDH.n398 GND 0.0193f
C4492 VDDH.n399 GND 0.09451f
C4493 VDDH.n400 GND 0.09451f
C4494 VDDH.t309 GND 0.08168f
C4495 VDDH.t139 GND 0.08378f
C4496 VDDH.t135 GND 0.08378f
C4497 VDDH.t134 GND 0.06284f
C4498 VDDH.t140 GND 0.08168f
C4499 VDDH.t130 GND 0.08378f
C4500 VDDH.t129 GND 0.08378f
C4501 VDDH.t127 GND 0.06284f
C4502 VDDH.n401 GND 0.02639f
C4503 VDDH.n404 GND 0.0277f
C4504 VDDH.n406 GND 0.02377f
C4505 VDDH.n407 GND 0.09451f
C4506 VDDH.n408 GND 0.09451f
C4507 VDDH.t223 GND 0.08168f
C4508 VDDH.t142 GND 0.08378f
C4509 VDDH.t225 GND 0.08378f
C4510 VDDH.t227 GND 0.06284f
C4511 VDDH.t191 GND 0.08168f
C4512 VDDH.t145 GND 0.08378f
C4513 VDDH.t144 GND 0.08378f
C4514 VDDH.t228 GND 0.06284f
C4515 VDDH.n409 GND 0.01943f
C4516 VDDH.n411 GND 0.03906f
C4517 VDDH.n413 GND 0.09451f
C4518 VDDH.n414 GND 0.09451f
C4519 VDDH.t70 GND 0.08168f
C4520 VDDH.t239 GND 0.08378f
C4521 VDDH.t73 GND 0.08378f
C4522 VDDH.t98 GND 0.06284f
C4523 VDDH.t238 GND 0.08168f
C4524 VDDH.t97 GND 0.08378f
C4525 VDDH.t72 GND 0.08378f
C4526 VDDH.t71 GND 0.06284f
C4527 VDDH.n415 GND 0.03156f
C4528 VDDH.n416 GND 0.02115f
C4529 VDDH.n417 GND 0.02005f
C4530 VDDH.n418 GND 0.03958f
C4531 VDDH.n419 GND 0.02001f
C4532 VDDH.n420 GND 0.03958f
C4533 VDDH.n421 GND 0.01351f
C4534 VDDH.n422 GND 0.09451f
C4535 VDDH.t282 GND 0.08168f
C4536 VDDH.t99 GND 0.08378f
C4537 VDDH.t103 GND 0.08378f
C4538 VDDH.t104 GND 0.06284f
C4539 VDDH.n423 GND 0.04189f
C4540 VDDH.t91 GND 0.06284f
C4541 VDDH.t102 GND 0.08378f
C4542 VDDH.t285 GND 0.08378f
C4543 VDDH.t283 GND 0.08168f
C4544 VDDH.n424 GND 0.09451f
C4545 VDDH.n426 GND 0.02319f
C4546 VDDH.n427 GND 0.01535f
C4547 VDDH.n428 GND 0.02489f
C4548 VDDH.n429 GND 0.12061f
C4549 VDDH.n430 GND 0.12061f
C4550 VDDH.t112 GND 0.08168f
C4551 VDDH.t113 GND 0.08378f
C4552 VDDH.t267 GND 0.08378f
C4553 VDDH.t111 GND 0.08803f
C4554 VDDH.t275 GND 0.08803f
C4555 VDDH.t276 GND 0.08378f
C4556 VDDH.t166 GND 0.06921f
C4557 VDDH.t48 GND 0.08593f
C4558 VDDH.t43 GND 0.09228f
C4559 VDDH.t37 GND 0.08803f
C4560 VDDH.t188 GND 0.08803f
C4561 VDDH.t190 GND 0.08803f
C4562 VDDH.t189 GND 0.08803f
C4563 VDDH.t165 GND 0.06071f
C4564 VDDH.n431 GND 0.02115f
C4565 VDDH.n432 GND 0.03857f
C4566 VDDH.n433 GND 0.06549f
C4567 VDDH.n434 GND 0.04189f
C4568 VDDH.n435 GND 0.06549f
C4569 VDDH.n436 GND 0.03526f
C4570 VDDH.n437 GND 0.02489f
C4571 VDDH.n439 GND 0.01703f
C4572 VDDH.n440 GND 0.0137f
C4573 VDDH.n441 GND 0.03958f
C4574 VDDH.n442 GND 0.04189f
C4575 VDDH.n443 GND 0.03958f
C4576 VDDH.n444 GND 0.02001f
C4577 VDDH.n445 GND 0.03906f
C4578 VDDH.n446 GND 0.01451f
C4579 VDDH.n447 GND 0.01781f
C4580 VDDH.n448 GND 0.09451f
C4581 VDDH.n450 GND 0.09451f
C4582 VDDH.t128 GND 0.08168f
C4583 VDDH.t136 GND 0.08378f
C4584 VDDH.t138 GND 0.08378f
C4585 VDDH.t132 GND 0.06284f
C4586 VDDH.n451 GND 0.02001f
C4587 VDDH.n452 GND 0.03958f
C4588 VDDH.t133 GND 0.08168f
C4589 VDDH.t131 GND 0.08378f
C4590 VDDH.t137 GND 0.08378f
C4591 VDDH.t308 GND 0.06284f
C4592 VDDH.n453 GND 0.04189f
C4593 VDDH.n454 GND 0.03958f
C4594 VDDH.n455 GND 0.01375f
C4595 VDDH.n456 GND 0.01751f
C4596 VDDH.n457 GND 0.01621f
C4597 VDDH.n458 GND 0.01538f
C4598 VDDH.n459 GND 0.01751f
C4599 VDDH.n460 GND 0.01625f
C4600 VDDH.n461 GND 0.03958f
C4601 VDDH.n462 GND 0.04189f
C4602 VDDH.n463 GND 0.03958f
C4603 VDDH.n464 GND 0.02168f
C4604 VDDH.n465 GND 0.0277f
C4605 VDDH.n466 GND 0.01944f
C4606 VDDH.n467 GND 0.09451f
C4607 VDDH.n468 GND 0.09451f
C4608 VDDH.t143 GND 0.08168f
C4609 VDDH.t193 GND 0.08378f
C4610 VDDH.t195 GND 0.08378f
C4611 VDDH.t196 GND 0.06284f
C4612 VDDH.n469 GND 0.01917f
C4613 VDDH.n470 GND 0.0193f
C4614 VDDH.n471 GND 0.02168f
C4615 VDDH.n472 GND 0.03958f
C4616 VDDH.t222 GND 0.08168f
C4617 VDDH.t226 GND 0.08378f
C4618 VDDH.t194 GND 0.08378f
C4619 VDDH.t192 GND 0.06284f
C4620 VDDH.n473 GND 0.04189f
C4621 VDDH.n474 GND 0.03958f
C4622 VDDH.n476 GND 0.01775f
C4623 VDDH.n477 GND 0.01556f
C4624 VDDH.n478 GND 0.01538f
C4625 VDDH.n479 GND 0.01775f
C4626 VDDH.n480 GND 0.01526f
C4627 VDDH.n481 GND 0.01775f
C4628 VDDH.n483 GND 0.03958f
C4629 VDDH.n484 GND 0.04189f
C4630 VDDH.n485 GND 0.03958f
C4631 VDDH.n486 GND 0.02001f
C4632 VDDH.n487 GND 0.01835f
C4633 VDDH.n488 GND 0.01835f
C4634 VDDH.n490 GND 0.01778f
C4635 VDDH.n491 GND 0.02001f
C4636 VDDH.n492 GND 0.03958f
C4637 VDDH.t201 GND 0.08168f
C4638 VDDH.t199 GND 0.08378f
C4639 VDDH.t198 GND 0.08378f
C4640 VDDH.t202 GND 0.06284f
C4641 VDDH.n493 GND 0.04189f
C4642 VDDH.n494 GND 0.03958f
C4643 VDDH.n496 GND 0.01775f
C4644 VDDH.n497 GND 0.02579f
C4645 VDDH.n498 GND 0.02001f
C4646 VDDH.n499 GND 0.03958f
C4647 VDDH.t124 GND 0.08168f
C4648 VDDH.t298 GND 0.08378f
C4649 VDDH.t296 GND 0.08378f
C4650 VDDH.t295 GND 0.06284f
C4651 VDDH.n500 GND 0.04189f
C4652 VDDH.n501 GND 0.03958f
C4653 VDDH.n502 GND 0.01917f
C4654 VDDH.n503 GND 0.01751f
C4655 VDDH.n506 GND 0.01805f
C4656 VDDH.n507 GND 0.02168f
C4657 VDDH.n508 GND 0.03958f
C4658 VDDH.n509 GND 0.04189f
C4659 VDDH.n510 GND 0.03958f
C4660 VDDH.n511 GND 0.02001f
C4661 VDDH.n512 GND 0.01457f
C4662 VDDH.n513 GND 0.0151f
C4663 VDDH.n514 GND 0.01443f
C4664 VDDH.n516 GND 0.09451f
C4665 VDDH.t108 GND 0.08168f
C4666 VDDH.t94 GND 0.08378f
C4667 VDDH.t117 GND 0.08378f
C4668 VDDH.t119 GND 0.06284f
C4669 VDDH.t96 GND 0.08168f
C4670 VDDH.t95 GND 0.08378f
C4671 VDDH.t116 GND 0.08378f
C4672 VDDH.t93 GND 0.06284f
C4673 VDDH.n517 GND 0.03958f
C4674 VDDH.n518 GND 0.04189f
C4675 VDDH.n519 GND 0.03958f
C4676 VDDH.n520 GND 0.02168f
C4677 VDDH.n521 GND 0.07771f
C4678 VDDH.n522 GND 3.8727f
C4679 VDDH.t208 GND 0.02075f
C4680 VDDH.n523 GND 0.43289f
C4681 VDDH.n524 GND 5.52519f
C4682 VDDH.n525 GND 7.97003f
C4683 VDDH.n526 GND 0.39499f
C4684 VDDH.n527 GND 0.03163f
C4685 VDDH.n531 GND 0.02091f
C4686 VDDH.n536 GND 0.0237f
C4687 VDDH.n537 GND 0.03029f
C4688 VDDH.n538 GND 0.03048f
C4689 VDDH.n539 GND 0.03048f
C4690 VDDH.n540 GND 0.03029f
C4691 VDDH.t301 GND 0.06847f
C4692 VDDH.n541 GND 0.0237f
C4693 VDDH.n546 GND 0.03163f
C4694 VDDH.n547 GND 0.17149f
C4695 VDDH.n548 GND 0.17589f
C4696 VDDH.n550 GND 0.02091f
C4697 VDDH.n552 GND 0.03612f
C4698 VDDH.n553 GND 0.03048f
C4699 VDDH.n554 GND 0.03029f
C4700 VDDH.t229 GND 0.04465f
C4701 VDDH.t69 GND 0.07348f
C4702 VDDH.t209 GND 0.07546f
C4703 VDDH.n555 GND 0.04493f
C4704 VDDH.n561 GND 0.03063f
C4705 VDDH.n563 GND 0.02091f
C4706 VDDH.n566 GND 0.0225f
C4707 VDDH.n569 GND 0.04469f
C4708 VDDH.t175 GND 0.07321f
C4709 VDDH.t310 GND 0.07343f
C4710 VDDH.n570 GND 0.04493f
C4711 VDDH.n571 GND 0.02444f
C4712 VDDH.n574 GND 0.02691f
C4713 VDDH.n575 GND 0.0237f
C4714 VDDH.n576 GND 0.03048f
C4715 VDDH.n577 GND 0.03063f
C4716 VDDH.n578 GND 0.02091f
C4717 VDDH.n584 GND 0.0225f
C4718 VDDH.n585 GND 0.17589f
C4719 VDDH.n586 GND 0.17589f
C4720 VDDH.n588 GND 0.02091f
C4721 VDDH.n594 GND 0.02691f
C4722 VDDH.n595 GND 0.0237f
C4723 VDDH.n596 GND 0.03048f
C4724 VDDH.n597 GND 0.03063f
C4725 VDDH.n599 GND 0.02091f
C4726 VDDH.n602 GND 0.0225f
C4727 VDDH.n605 GND 0.04469f
C4728 VDDH.t9 GND 0.07321f
C4729 VDDH.t75 GND 0.07343f
C4730 VDDH.n606 GND 0.04493f
C4731 VDDH.n612 GND 0.03063f
C4732 VDDH.n614 GND 0.02091f
C4733 VDDH.n617 GND 0.0225f
C4734 VDDH.n620 GND 0.04469f
C4735 VDDH.t221 GND 0.07321f
C4736 VDDH.t274 GND 0.07343f
C4737 VDDH.n621 GND 0.04493f
C4738 VDDH.n622 GND 0.02444f
C4739 VDDH.n625 GND 0.02691f
C4740 VDDH.n626 GND 0.0237f
C4741 VDDH.n627 GND 0.03048f
C4742 VDDH.n628 GND 0.03063f
C4743 VDDH.n629 GND 0.02091f
C4744 VDDH.n635 GND 0.0225f
C4745 VDDH.n636 GND 0.19516f
C4746 VDDH.n637 GND 0.06935f
C4747 VDDH.n638 GND 0.01129f
C4748 VDDH.n644 GND 0.02091f
C4749 VDDH.n646 GND 0.01129f
C4750 VDDH.n651 GND 0.1168f
C4751 VDDH.n657 GND 0.02091f
C4752 VDDH.n659 GND 0.03019f
C4753 VDDH.n660 GND 0.02589f
C4754 VDDH.n661 GND 0.01673f
C4755 VDDH.n662 GND 0.02892f
C4756 VDDH.n663 GND 0.02735f
C4757 VDDH.n664 GND 0.03019f
C4758 VDDH.n665 GND 0.02589f
C4759 VDDH.n666 GND 0.01673f
C4760 VDDH.n667 GND 0.04543f
C4761 VDDH.n668 GND 0.26477f
C4762 VDDH.t41 GND 0.33952f
C4763 VDDH.t180 GND 0.23053f
C4764 VDDH.t294 GND 0.1888f
C4765 VDDH.n670 GND 0.17042f
C4766 VDDH.t204 GND 0.30488f
C4767 VDDH.t32 GND 0.38014f
C4768 VDDH.n671 GND 0.27524f
C4769 VDDH.t148 GND 1.70981f
C4770 VDDH.t44 GND 0.09002f
C4771 VDDH.n672 GND 0.40183f
C4772 VDDH.n673 GND 0.04719f
C4773 VDDH.n674 GND 0.02289f
C4774 VDDH.n675 GND 0.05045f
C4775 VDDH.n676 GND 0.05605f
C4776 VDDH.n677 GND 0.08459f
C4777 VDDH.n679 GND 0.03275f
C4778 VDDH.n680 GND 0.01306f
C4779 VDDH.n682 GND 0.01317f
C4780 VDDH.n683 GND 0.02881f
C4781 VDDH.n684 GND 0.03156f
C4782 VDDH.n685 GND 0.02679f
C4783 VDDH.n686 GND 0.01415f
C4784 VDDH.n687 GND 0.05506f
C4785 VDDH.n688 GND 0.07563f
C4786 VDDH.n689 GND 0.02916f
C4787 VDDH.n690 GND 0.03283f
C4788 VDDH.n691 GND 0.02807f
C4789 VDDH.n692 GND 0.04941f
C4790 VDDH.n693 GND 0.33709f
C4791 VDDH.t154 GND 0.41901f
C4792 VDDH.t155 GND 0.41901f
C4793 VDDH.n694 GND 0.45072f
C4794 VDDH.n695 GND 0.02081f
C4795 VDDH.n698 GND 0.03292f
C4796 VDDH.n699 GND 0.03478f
C4797 VDDH.n700 GND 0.05343f
C4798 VDDH.n701 GND 0.04505f
C4799 VDDH.n702 GND 0.02587f
C4800 VDDH.n703 GND 0.02416f
C4801 VDDH.n704 GND 0.01668f
C4802 VDDH.n705 GND 0.04355f
C4803 VDDH.n706 GND 0.02099f
C4804 top_segment_3_0.b[5].t0 GND 0.09866f
C4805 top_segment_3_0.b[5].n0 GND 0.04045f
C4806 top_segment_3_0.b[5].n1 GND 0.08708f
C4807 top_segment_3_0.b[5].n2 GND 0.05782f
C4808 top_segment_3_0.b[5].t1 GND 0.09452f
C4809 top_segment_3_0.b[5].n3 GND 0.01194f
C4810 top_segment_3_0.b[5].t2 GND 0.19507f
C4811 top_segment_3_0.b[5].n4 GND 0.25416f
C4812 top_segment_3_0.b[5].t5 GND 0.19507f
C4813 top_segment_3_0.b[5].n5 GND 0.30624f
C4814 top_segment_3_0.b[5].t4 GND 0.196f
C4815 top_segment_3_0.b[5].t6 GND 0.19507f
C4816 top_segment_3_0.b[5].n6 GND 0.61154f
C4817 top_segment_3_0.b[5].n7 GND 0.20386f
C4818 top_segment_3_0.b[5].t3 GND 0.1929f
C4819 top_segment_3_0.b[5].n8 GND 13.9648f
C4820 top_segment_3_0.b[5].n9 GND 0.06224f
C4821 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t1 GND 0.04119f
C4822 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t7 GND 0.03353f
C4823 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t8 GND 0.02094f
C4824 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n0 GND 0.06383f
C4825 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n1 GND 0.03879f
C4826 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t4 GND 0.03353f
C4827 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t6 GND 0.02094f
C4828 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n2 GND 0.06383f
C4829 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n3 GND 0.01711f
C4830 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n4 GND 0.35016f
C4831 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n5 GND 4.38855f
C4832 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n6 GND 0.18482f
C4833 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t2 GND 0.02026f
C4834 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t3 GND 0.02026f
C4835 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n7 GND 0.04503f
C4836 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t0 GND 0.07496f
C4837 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t9 GND 0.02096f
C4838 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].t5 GND 0.03356f
C4839 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n8 GND 0.06289f
C4840 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n9 GND 0.05268f
C4841 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n10 GND 0.14872f
C4842 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.decoder_3_0/decoder_2to4_2.b[0].n11 GND 0.12975f
C4843 VDD.n0 GND 0.01865f
C4844 VDD.n15 GND 0.01039f
C4845 VDD.n19 GND 0.01039f
C4846 VDD.n23 GND 0.01039f
C4847 VDD.n27 GND 0.01039f
C4848 VDD.n31 GND 0.01039f
C4849 VDD.n35 GND 0.01039f
C4850 VDD.n39 GND 0.01039f
C4851 VDD.n43 GND 0.01039f
C4852 VDD.n46 GND 0.14175f
C4853 VDD.n47 GND 3.73304f
C4854 VDD.n81 GND 0.01746f
C4855 VDD.t182 GND 0.01144f
C4856 VDD.n83 GND 0.01545f
C4857 VDD.n84 GND 0.01268f
C4858 VDD.n89 GND 0.02837f
C4859 VDD.n115 GND 0.01268f
C4860 VDD.n141 GND 0.01337f
C4861 VDD.n142 GND 0.01545f
C4862 VDD.n147 GND 0.02837f
C4863 VDD.n148 GND 0.10888f
C4864 VDD.n149 GND 0.19392f
C4865 VDD.n150 GND 6.89573f
C4866 VDD.n153 GND 0.06728f
C4867 VDD.t14 GND 0.02779f
C4868 VDD.n161 GND 0.04824f
C4869 VDD.t43 GND 0.02779f
C4870 VDD.n163 GND 0.06697f
C4871 VDD.n198 GND 0.01889f
C4872 VDD.t174 GND 0.01066f
C4873 VDD.t71 GND 0.01533f
C4874 VDD.t67 GND 0.01428f
C4875 VDD.n238 GND 0.01452f
C4876 VDD.n276 GND 0.01224f
C4877 VDD.t169 GND 0.0123f
C4878 VDD.n277 GND 0.01013f
C4879 VDD.n279 GND 0.02586f
C4880 VDD.n280 GND 0.03539f
C4881 VDD.n282 GND 0.01917f
C4882 VDD.n295 GND 0.01031f
C4883 VDD.t161 GND 0.01037f
C4884 VDD.n312 GND 0.01091f
C4885 VDD.t69 GND 0.02901f
C4886 VDD.n313 GND 0.02981f
C4887 VDD.n314 GND 0.01287f
C4888 VDD.n315 GND 0.0662f
C4889 VDD.n316 GND 0.02986f
C4890 VDD.n317 GND 0.01332f
C4891 VDD.n331 GND 0.03982f
C4892 VDD.n335 GND 0.09635f
C4893 VDD.n336 GND 0.0844f
C4894 VDD.n337 GND 4.61645f
C4895 VDD.n338 GND 1.73773f
C4896 VDD.n339 GND 0.20085f
C4897 VDD.n439 GND 0.01039f
C4898 VDD.t98 GND 0.0143f
C4899 VDD.n440 GND 0.01387f
C4900 a_26719_5238.t1 GND 0.12364f
C4901 a_26719_5238.t3 GND 0.07206f
C4902 a_26719_5238.n0 GND 4.94854f
C4903 a_26719_5238.t4 GND 0.15859f
C4904 a_26719_5238.n1 GND 4.24803f
C4905 a_26719_5238.t2 GND 0.15202f
C4906 a_26719_5238.n2 GND 4.62506f
C4907 a_26719_5238.t0 GND 0.07206f
C4908 top_segment_2_0.DEC2[1].t0 GND 0.10226f
C4909 top_segment_2_0.DEC2[1].t1 GND 0.08695f
C4910 top_segment_2_0.DEC2[1].n0 GND 0.69951f
C4911 top_segment_2_0.DEC2[1].t17 GND 0.40597f
C4912 top_segment_2_0.DEC2[1].t7 GND 0.4043f
C4913 top_segment_2_0.DEC2[1].n1 GND 0.64174f
C4914 top_segment_2_0.DEC2[1].n2 GND 0.414f
C4915 top_segment_2_0.DEC2[1].t4 GND 0.42696f
C4916 top_segment_2_0.DEC2[1].n3 GND 0.89278f
C4917 top_segment_2_0.DEC2[1].t20 GND 0.12394f
C4918 top_segment_2_0.DEC2[1].t15 GND 0.12224f
C4919 top_segment_2_0.DEC2[1].n4 GND 5.66133f
C4920 top_segment_2_0.DEC2[1].t16 GND 0.12429f
C4921 top_segment_2_0.DEC2[1].t19 GND 0.12366f
C4922 top_segment_2_0.DEC2[1].n5 GND 0.4028f
C4923 top_segment_2_0.DEC2[1].t9 GND 0.12366f
C4924 top_segment_2_0.DEC2[1].n6 GND 0.20171f
C4925 top_segment_2_0.DEC2[1].t22 GND 0.12366f
C4926 top_segment_2_0.DEC2[1].n7 GND 0.20171f
C4927 top_segment_2_0.DEC2[1].t3 GND 0.12366f
C4928 top_segment_2_0.DEC2[1].n8 GND 0.20171f
C4929 top_segment_2_0.DEC2[1].t8 GND 0.12366f
C4930 top_segment_2_0.DEC2[1].n9 GND 0.20171f
C4931 top_segment_2_0.DEC2[1].t11 GND 0.12366f
C4932 top_segment_2_0.DEC2[1].n10 GND 0.20171f
C4933 top_segment_2_0.DEC2[1].n11 GND 0.09544f
C4934 top_segment_2_0.DEC2[1].t12 GND 0.12224f
C4935 top_segment_2_0.DEC2[1].n12 GND 0.10215f
C4936 top_segment_2_0.DEC2[1].t24 GND 0.12429f
C4937 top_segment_2_0.DEC2[1].t13 GND 0.12471f
C4938 top_segment_2_0.DEC2[1].t10 GND 0.12403f
C4939 top_segment_2_0.DEC2[1].n13 GND 0.43623f
C4940 top_segment_2_0.DEC2[1].t5 GND 0.12403f
C4941 top_segment_2_0.DEC2[1].n14 GND 0.21846f
C4942 top_segment_2_0.DEC2[1].t2 GND 0.12403f
C4943 top_segment_2_0.DEC2[1].n15 GND 0.21846f
C4944 top_segment_2_0.DEC2[1].t23 GND 0.12403f
C4945 top_segment_2_0.DEC2[1].n16 GND 0.21846f
C4946 top_segment_2_0.DEC2[1].t6 GND 0.12403f
C4947 top_segment_2_0.DEC2[1].n17 GND 0.21846f
C4948 top_segment_2_0.DEC2[1].n18 GND 0.33687f
C4949 top_segment_2_0.DEC2[1].t18 GND 0.12224f
C4950 top_segment_2_0.DEC2[1].n19 GND 0.42787f
C4951 top_segment_2_0.DEC2[1].n20 GND 2.49587f
C4952 top_segment_2_0.DEC2[1].n21 GND 11.4725f
C4953 top_segment_2_0.DEC2[1].t21 GND 0.22982f
C4954 top_segment_2_0.DEC2[1].t14 GND 0.12749f
C4955 top_segment_2_0.DEC2[1].n22 GND 0.20027f
C4956 top_segment_2_0.DEC2[1].n23 GND 0.03496f
C4957 top_segment_2_0.DEC2[1].n24 GND 0.27468f
C4958 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t8 GND 0.07099f
C4959 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t15 GND 0.0702f
C4960 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n0 GND 0.14656f
C4961 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t16 GND 0.0702f
C4962 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n1 GND 0.06927f
C4963 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t20 GND 0.0702f
C4964 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n2 GND 0.06927f
C4965 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t21 GND 0.0702f
C4966 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n3 GND 0.06927f
C4967 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t25 GND 0.0702f
C4968 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n4 GND 0.06927f
C4969 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t26 GND 0.0702f
C4970 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n5 GND 0.06927f
C4971 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t9 GND 0.0702f
C4972 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n6 GND 0.06927f
C4973 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t10 GND 0.0702f
C4974 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n7 GND 0.06927f
C4975 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t28 GND 0.0702f
C4976 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n8 GND 0.06927f
C4977 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t6 GND 0.0702f
C4978 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n9 GND 0.06927f
C4979 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t11 GND 0.0702f
C4980 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n10 GND 0.06927f
C4981 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t12 GND 0.0702f
C4982 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n11 GND 0.06927f
C4983 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t17 GND 0.0702f
C4984 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n12 GND 0.06927f
C4985 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t18 GND 0.0702f
C4986 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n13 GND 0.06927f
C4987 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t22 GND 0.0702f
C4988 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n14 GND 0.06927f
C4989 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t23 GND 0.0702f
C4990 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n15 GND 0.06927f
C4991 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t7 GND 0.0702f
C4992 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n16 GND 0.06927f
C4993 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t13 GND 0.0702f
C4994 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n17 GND 0.06927f
C4995 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t14 GND 0.0702f
C4996 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n18 GND 0.06927f
C4997 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t19 GND 0.0702f
C4998 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n19 GND 0.06927f
C4999 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t24 GND 0.0702f
C5000 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n20 GND 0.06641f
C5001 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t27 GND 0.27283f
C5002 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n21 GND 0.09448f
C5003 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n22 GND 0.55544f
C5004 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t4 GND 0.04839f
C5005 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n23 GND 0.0364f
C5006 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n24 GND 0.04636f
C5007 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t2 GND 0.04832f
C5008 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n25 GND 0.02822f
C5009 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n26 GND 0.18252f
C5010 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t1 GND 0.0317f
C5011 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n27 GND 0.18304f
C5012 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.t0 GND 0.03062f
C5013 top_dcell_routing_0.top_dcell_bias_0/top_digital_cell_0.VBNLV.n28 GND 0.1181f
.ends

